// This is the unpowered netlist.
module des_Trojan (clk,
    decrypt,
    finish,
    init,
    reset,
    desIn,
    desOut_ff,
    key);
 input clk;
 input decrypt;
 output finish;
 input init;
 input reset;
 input [63:0] desIn;
 output [63:0] desOut_ff;
 input [55:0] key;

 wire \FP[10] ;
 wire \FP[11] ;
 wire \FP[12] ;
 wire \FP[13] ;
 wire \FP[14] ;
 wire \FP[15] ;
 wire \FP[16] ;
 wire \FP[17] ;
 wire \FP[18] ;
 wire \FP[19] ;
 wire \FP[1] ;
 wire \FP[20] ;
 wire \FP[21] ;
 wire \FP[22] ;
 wire \FP[23] ;
 wire \FP[24] ;
 wire \FP[25] ;
 wire \FP[26] ;
 wire \FP[27] ;
 wire \FP[28] ;
 wire \FP[29] ;
 wire \FP[2] ;
 wire \FP[30] ;
 wire \FP[31] ;
 wire \FP[32] ;
 wire \FP[3] ;
 wire \FP[4] ;
 wire \FP[5] ;
 wire \FP[6] ;
 wire \FP[7] ;
 wire \FP[8] ;
 wire \FP[9] ;
 wire \L[10] ;
 wire \L[11] ;
 wire \L[12] ;
 wire \L[13] ;
 wire \L[14] ;
 wire \L[15] ;
 wire \L[16] ;
 wire \L[17] ;
 wire \L[18] ;
 wire \L[19] ;
 wire \L[1] ;
 wire \L[20] ;
 wire \L[21] ;
 wire \L[22] ;
 wire \L[23] ;
 wire \L[24] ;
 wire \L[25] ;
 wire \L[26] ;
 wire \L[27] ;
 wire \L[28] ;
 wire \L[29] ;
 wire \L[2] ;
 wire \L[30] ;
 wire \L[31] ;
 wire \L[32] ;
 wire \L[3] ;
 wire \L[4] ;
 wire \L[5] ;
 wire \L[6] ;
 wire \L[7] ;
 wire \L[8] ;
 wire \L[9] ;
 wire \R[10] ;
 wire \R[11] ;
 wire \R[12] ;
 wire \R[13] ;
 wire \R[14] ;
 wire \R[15] ;
 wire \R[16] ;
 wire \R[17] ;
 wire \R[18] ;
 wire \R[19] ;
 wire \R[1] ;
 wire \R[20] ;
 wire \R[21] ;
 wire \R[22] ;
 wire \R[23] ;
 wire \R[24] ;
 wire \R[25] ;
 wire \R[26] ;
 wire \R[27] ;
 wire \R[28] ;
 wire \R[29] ;
 wire \R[2] ;
 wire \R[30] ;
 wire \R[31] ;
 wire \R[32] ;
 wire \R[3] ;
 wire \R[4] ;
 wire \R[5] ;
 wire \R[6] ;
 wire \R[7] ;
 wire \R[8] ;
 wire \R[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \counter_inst.count[0] ;
 wire \counter_inst.count[1] ;
 wire \counter_inst.count[2] ;
 wire \counter_inst.count[3] ;
 wire \counter_inst.count[4] ;
 wire \fifo.fifo[0][0] ;
 wire \fifo.fifo[0][10] ;
 wire \fifo.fifo[0][11] ;
 wire \fifo.fifo[0][12] ;
 wire \fifo.fifo[0][13] ;
 wire \fifo.fifo[0][14] ;
 wire \fifo.fifo[0][15] ;
 wire \fifo.fifo[0][16] ;
 wire \fifo.fifo[0][17] ;
 wire \fifo.fifo[0][18] ;
 wire \fifo.fifo[0][19] ;
 wire \fifo.fifo[0][1] ;
 wire \fifo.fifo[0][20] ;
 wire \fifo.fifo[0][21] ;
 wire \fifo.fifo[0][22] ;
 wire \fifo.fifo[0][23] ;
 wire \fifo.fifo[0][24] ;
 wire \fifo.fifo[0][25] ;
 wire \fifo.fifo[0][26] ;
 wire \fifo.fifo[0][27] ;
 wire \fifo.fifo[0][28] ;
 wire \fifo.fifo[0][29] ;
 wire \fifo.fifo[0][2] ;
 wire \fifo.fifo[0][30] ;
 wire \fifo.fifo[0][31] ;
 wire \fifo.fifo[0][32] ;
 wire \fifo.fifo[0][33] ;
 wire \fifo.fifo[0][34] ;
 wire \fifo.fifo[0][35] ;
 wire \fifo.fifo[0][36] ;
 wire \fifo.fifo[0][37] ;
 wire \fifo.fifo[0][38] ;
 wire \fifo.fifo[0][39] ;
 wire \fifo.fifo[0][3] ;
 wire \fifo.fifo[0][40] ;
 wire \fifo.fifo[0][41] ;
 wire \fifo.fifo[0][42] ;
 wire \fifo.fifo[0][43] ;
 wire \fifo.fifo[0][44] ;
 wire \fifo.fifo[0][45] ;
 wire \fifo.fifo[0][46] ;
 wire \fifo.fifo[0][47] ;
 wire \fifo.fifo[0][48] ;
 wire \fifo.fifo[0][49] ;
 wire \fifo.fifo[0][4] ;
 wire \fifo.fifo[0][50] ;
 wire \fifo.fifo[0][51] ;
 wire \fifo.fifo[0][52] ;
 wire \fifo.fifo[0][53] ;
 wire \fifo.fifo[0][54] ;
 wire \fifo.fifo[0][55] ;
 wire \fifo.fifo[0][5] ;
 wire \fifo.fifo[0][6] ;
 wire \fifo.fifo[0][7] ;
 wire \fifo.fifo[0][8] ;
 wire \fifo.fifo[0][9] ;
 wire \fifo.fifo[1][0] ;
 wire \fifo.fifo[1][10] ;
 wire \fifo.fifo[1][11] ;
 wire \fifo.fifo[1][12] ;
 wire \fifo.fifo[1][13] ;
 wire \fifo.fifo[1][14] ;
 wire \fifo.fifo[1][15] ;
 wire \fifo.fifo[1][16] ;
 wire \fifo.fifo[1][17] ;
 wire \fifo.fifo[1][18] ;
 wire \fifo.fifo[1][19] ;
 wire \fifo.fifo[1][1] ;
 wire \fifo.fifo[1][20] ;
 wire \fifo.fifo[1][21] ;
 wire \fifo.fifo[1][22] ;
 wire \fifo.fifo[1][23] ;
 wire \fifo.fifo[1][24] ;
 wire \fifo.fifo[1][25] ;
 wire \fifo.fifo[1][26] ;
 wire \fifo.fifo[1][27] ;
 wire \fifo.fifo[1][28] ;
 wire \fifo.fifo[1][29] ;
 wire \fifo.fifo[1][2] ;
 wire \fifo.fifo[1][30] ;
 wire \fifo.fifo[1][31] ;
 wire \fifo.fifo[1][32] ;
 wire \fifo.fifo[1][33] ;
 wire \fifo.fifo[1][34] ;
 wire \fifo.fifo[1][35] ;
 wire \fifo.fifo[1][36] ;
 wire \fifo.fifo[1][37] ;
 wire \fifo.fifo[1][38] ;
 wire \fifo.fifo[1][39] ;
 wire \fifo.fifo[1][3] ;
 wire \fifo.fifo[1][40] ;
 wire \fifo.fifo[1][41] ;
 wire \fifo.fifo[1][42] ;
 wire \fifo.fifo[1][43] ;
 wire \fifo.fifo[1][44] ;
 wire \fifo.fifo[1][45] ;
 wire \fifo.fifo[1][46] ;
 wire \fifo.fifo[1][47] ;
 wire \fifo.fifo[1][48] ;
 wire \fifo.fifo[1][49] ;
 wire \fifo.fifo[1][4] ;
 wire \fifo.fifo[1][50] ;
 wire \fifo.fifo[1][51] ;
 wire \fifo.fifo[1][52] ;
 wire \fifo.fifo[1][53] ;
 wire \fifo.fifo[1][54] ;
 wire \fifo.fifo[1][55] ;
 wire \fifo.fifo[1][5] ;
 wire \fifo.fifo[1][6] ;
 wire \fifo.fifo[1][7] ;
 wire \fifo.fifo[1][8] ;
 wire \fifo.fifo[1][9] ;
 wire \fifo.fifo[2][0] ;
 wire \fifo.fifo[2][10] ;
 wire \fifo.fifo[2][11] ;
 wire \fifo.fifo[2][12] ;
 wire \fifo.fifo[2][13] ;
 wire \fifo.fifo[2][14] ;
 wire \fifo.fifo[2][15] ;
 wire \fifo.fifo[2][16] ;
 wire \fifo.fifo[2][17] ;
 wire \fifo.fifo[2][18] ;
 wire \fifo.fifo[2][19] ;
 wire \fifo.fifo[2][1] ;
 wire \fifo.fifo[2][20] ;
 wire \fifo.fifo[2][21] ;
 wire \fifo.fifo[2][22] ;
 wire \fifo.fifo[2][23] ;
 wire \fifo.fifo[2][24] ;
 wire \fifo.fifo[2][25] ;
 wire \fifo.fifo[2][26] ;
 wire \fifo.fifo[2][27] ;
 wire \fifo.fifo[2][28] ;
 wire \fifo.fifo[2][29] ;
 wire \fifo.fifo[2][2] ;
 wire \fifo.fifo[2][30] ;
 wire \fifo.fifo[2][31] ;
 wire \fifo.fifo[2][32] ;
 wire \fifo.fifo[2][33] ;
 wire \fifo.fifo[2][34] ;
 wire \fifo.fifo[2][35] ;
 wire \fifo.fifo[2][36] ;
 wire \fifo.fifo[2][37] ;
 wire \fifo.fifo[2][38] ;
 wire \fifo.fifo[2][39] ;
 wire \fifo.fifo[2][3] ;
 wire \fifo.fifo[2][40] ;
 wire \fifo.fifo[2][41] ;
 wire \fifo.fifo[2][42] ;
 wire \fifo.fifo[2][43] ;
 wire \fifo.fifo[2][44] ;
 wire \fifo.fifo[2][45] ;
 wire \fifo.fifo[2][46] ;
 wire \fifo.fifo[2][47] ;
 wire \fifo.fifo[2][48] ;
 wire \fifo.fifo[2][49] ;
 wire \fifo.fifo[2][4] ;
 wire \fifo.fifo[2][50] ;
 wire \fifo.fifo[2][51] ;
 wire \fifo.fifo[2][52] ;
 wire \fifo.fifo[2][53] ;
 wire \fifo.fifo[2][54] ;
 wire \fifo.fifo[2][55] ;
 wire \fifo.fifo[2][5] ;
 wire \fifo.fifo[2][6] ;
 wire \fifo.fifo[2][7] ;
 wire \fifo.fifo[2][8] ;
 wire \fifo.fifo[2][9] ;
 wire \fifo.fifo[3][0] ;
 wire \fifo.fifo[3][10] ;
 wire \fifo.fifo[3][11] ;
 wire \fifo.fifo[3][12] ;
 wire \fifo.fifo[3][13] ;
 wire \fifo.fifo[3][14] ;
 wire \fifo.fifo[3][15] ;
 wire \fifo.fifo[3][16] ;
 wire \fifo.fifo[3][17] ;
 wire \fifo.fifo[3][18] ;
 wire \fifo.fifo[3][19] ;
 wire \fifo.fifo[3][1] ;
 wire \fifo.fifo[3][20] ;
 wire \fifo.fifo[3][21] ;
 wire \fifo.fifo[3][22] ;
 wire \fifo.fifo[3][23] ;
 wire \fifo.fifo[3][24] ;
 wire \fifo.fifo[3][25] ;
 wire \fifo.fifo[3][26] ;
 wire \fifo.fifo[3][27] ;
 wire \fifo.fifo[3][28] ;
 wire \fifo.fifo[3][29] ;
 wire \fifo.fifo[3][2] ;
 wire \fifo.fifo[3][30] ;
 wire \fifo.fifo[3][31] ;
 wire \fifo.fifo[3][32] ;
 wire \fifo.fifo[3][33] ;
 wire \fifo.fifo[3][34] ;
 wire \fifo.fifo[3][35] ;
 wire \fifo.fifo[3][36] ;
 wire \fifo.fifo[3][37] ;
 wire \fifo.fifo[3][38] ;
 wire \fifo.fifo[3][39] ;
 wire \fifo.fifo[3][3] ;
 wire \fifo.fifo[3][40] ;
 wire \fifo.fifo[3][41] ;
 wire \fifo.fifo[3][42] ;
 wire \fifo.fifo[3][43] ;
 wire \fifo.fifo[3][44] ;
 wire \fifo.fifo[3][45] ;
 wire \fifo.fifo[3][46] ;
 wire \fifo.fifo[3][47] ;
 wire \fifo.fifo[3][48] ;
 wire \fifo.fifo[3][49] ;
 wire \fifo.fifo[3][4] ;
 wire \fifo.fifo[3][50] ;
 wire \fifo.fifo[3][51] ;
 wire \fifo.fifo[3][52] ;
 wire \fifo.fifo[3][53] ;
 wire \fifo.fifo[3][54] ;
 wire \fifo.fifo[3][55] ;
 wire \fifo.fifo[3][5] ;
 wire \fifo.fifo[3][6] ;
 wire \fifo.fifo[3][7] ;
 wire \fifo.fifo[3][8] ;
 wire \fifo.fifo[3][9] ;
 wire \fifo.fifo[4][0] ;
 wire \fifo.fifo[4][10] ;
 wire \fifo.fifo[4][11] ;
 wire \fifo.fifo[4][12] ;
 wire \fifo.fifo[4][13] ;
 wire \fifo.fifo[4][14] ;
 wire \fifo.fifo[4][15] ;
 wire \fifo.fifo[4][16] ;
 wire \fifo.fifo[4][17] ;
 wire \fifo.fifo[4][18] ;
 wire \fifo.fifo[4][19] ;
 wire \fifo.fifo[4][1] ;
 wire \fifo.fifo[4][20] ;
 wire \fifo.fifo[4][21] ;
 wire \fifo.fifo[4][22] ;
 wire \fifo.fifo[4][23] ;
 wire \fifo.fifo[4][24] ;
 wire \fifo.fifo[4][25] ;
 wire \fifo.fifo[4][26] ;
 wire \fifo.fifo[4][27] ;
 wire \fifo.fifo[4][28] ;
 wire \fifo.fifo[4][29] ;
 wire \fifo.fifo[4][2] ;
 wire \fifo.fifo[4][30] ;
 wire \fifo.fifo[4][31] ;
 wire \fifo.fifo[4][32] ;
 wire \fifo.fifo[4][33] ;
 wire \fifo.fifo[4][34] ;
 wire \fifo.fifo[4][35] ;
 wire \fifo.fifo[4][36] ;
 wire \fifo.fifo[4][37] ;
 wire \fifo.fifo[4][38] ;
 wire \fifo.fifo[4][39] ;
 wire \fifo.fifo[4][3] ;
 wire \fifo.fifo[4][40] ;
 wire \fifo.fifo[4][41] ;
 wire \fifo.fifo[4][42] ;
 wire \fifo.fifo[4][43] ;
 wire \fifo.fifo[4][44] ;
 wire \fifo.fifo[4][45] ;
 wire \fifo.fifo[4][46] ;
 wire \fifo.fifo[4][47] ;
 wire \fifo.fifo[4][48] ;
 wire \fifo.fifo[4][49] ;
 wire \fifo.fifo[4][4] ;
 wire \fifo.fifo[4][50] ;
 wire \fifo.fifo[4][51] ;
 wire \fifo.fifo[4][52] ;
 wire \fifo.fifo[4][53] ;
 wire \fifo.fifo[4][54] ;
 wire \fifo.fifo[4][55] ;
 wire \fifo.fifo[4][5] ;
 wire \fifo.fifo[4][6] ;
 wire \fifo.fifo[4][7] ;
 wire \fifo.fifo[4][8] ;
 wire \fifo.fifo[4][9] ;
 wire \fifo.fifo[5][0] ;
 wire \fifo.fifo[5][10] ;
 wire \fifo.fifo[5][11] ;
 wire \fifo.fifo[5][12] ;
 wire \fifo.fifo[5][13] ;
 wire \fifo.fifo[5][14] ;
 wire \fifo.fifo[5][15] ;
 wire \fifo.fifo[5][16] ;
 wire \fifo.fifo[5][17] ;
 wire \fifo.fifo[5][18] ;
 wire \fifo.fifo[5][19] ;
 wire \fifo.fifo[5][1] ;
 wire \fifo.fifo[5][20] ;
 wire \fifo.fifo[5][21] ;
 wire \fifo.fifo[5][22] ;
 wire \fifo.fifo[5][23] ;
 wire \fifo.fifo[5][24] ;
 wire \fifo.fifo[5][25] ;
 wire \fifo.fifo[5][26] ;
 wire \fifo.fifo[5][27] ;
 wire \fifo.fifo[5][28] ;
 wire \fifo.fifo[5][29] ;
 wire \fifo.fifo[5][2] ;
 wire \fifo.fifo[5][30] ;
 wire \fifo.fifo[5][31] ;
 wire \fifo.fifo[5][32] ;
 wire \fifo.fifo[5][33] ;
 wire \fifo.fifo[5][34] ;
 wire \fifo.fifo[5][35] ;
 wire \fifo.fifo[5][36] ;
 wire \fifo.fifo[5][37] ;
 wire \fifo.fifo[5][38] ;
 wire \fifo.fifo[5][39] ;
 wire \fifo.fifo[5][3] ;
 wire \fifo.fifo[5][40] ;
 wire \fifo.fifo[5][41] ;
 wire \fifo.fifo[5][42] ;
 wire \fifo.fifo[5][43] ;
 wire \fifo.fifo[5][44] ;
 wire \fifo.fifo[5][45] ;
 wire \fifo.fifo[5][46] ;
 wire \fifo.fifo[5][47] ;
 wire \fifo.fifo[5][48] ;
 wire \fifo.fifo[5][49] ;
 wire \fifo.fifo[5][4] ;
 wire \fifo.fifo[5][50] ;
 wire \fifo.fifo[5][51] ;
 wire \fifo.fifo[5][52] ;
 wire \fifo.fifo[5][53] ;
 wire \fifo.fifo[5][54] ;
 wire \fifo.fifo[5][55] ;
 wire \fifo.fifo[5][5] ;
 wire \fifo.fifo[5][6] ;
 wire \fifo.fifo[5][7] ;
 wire \fifo.fifo[5][8] ;
 wire \fifo.fifo[5][9] ;
 wire \fifo.fifo[6][0] ;
 wire \fifo.fifo[6][10] ;
 wire \fifo.fifo[6][11] ;
 wire \fifo.fifo[6][12] ;
 wire \fifo.fifo[6][13] ;
 wire \fifo.fifo[6][14] ;
 wire \fifo.fifo[6][15] ;
 wire \fifo.fifo[6][16] ;
 wire \fifo.fifo[6][17] ;
 wire \fifo.fifo[6][18] ;
 wire \fifo.fifo[6][19] ;
 wire \fifo.fifo[6][1] ;
 wire \fifo.fifo[6][20] ;
 wire \fifo.fifo[6][21] ;
 wire \fifo.fifo[6][22] ;
 wire \fifo.fifo[6][23] ;
 wire \fifo.fifo[6][24] ;
 wire \fifo.fifo[6][25] ;
 wire \fifo.fifo[6][26] ;
 wire \fifo.fifo[6][27] ;
 wire \fifo.fifo[6][28] ;
 wire \fifo.fifo[6][29] ;
 wire \fifo.fifo[6][2] ;
 wire \fifo.fifo[6][30] ;
 wire \fifo.fifo[6][31] ;
 wire \fifo.fifo[6][32] ;
 wire \fifo.fifo[6][33] ;
 wire \fifo.fifo[6][34] ;
 wire \fifo.fifo[6][35] ;
 wire \fifo.fifo[6][36] ;
 wire \fifo.fifo[6][37] ;
 wire \fifo.fifo[6][38] ;
 wire \fifo.fifo[6][39] ;
 wire \fifo.fifo[6][3] ;
 wire \fifo.fifo[6][40] ;
 wire \fifo.fifo[6][41] ;
 wire \fifo.fifo[6][42] ;
 wire \fifo.fifo[6][43] ;
 wire \fifo.fifo[6][44] ;
 wire \fifo.fifo[6][45] ;
 wire \fifo.fifo[6][46] ;
 wire \fifo.fifo[6][47] ;
 wire \fifo.fifo[6][48] ;
 wire \fifo.fifo[6][49] ;
 wire \fifo.fifo[6][4] ;
 wire \fifo.fifo[6][50] ;
 wire \fifo.fifo[6][51] ;
 wire \fifo.fifo[6][52] ;
 wire \fifo.fifo[6][53] ;
 wire \fifo.fifo[6][54] ;
 wire \fifo.fifo[6][55] ;
 wire \fifo.fifo[6][5] ;
 wire \fifo.fifo[6][6] ;
 wire \fifo.fifo[6][7] ;
 wire \fifo.fifo[6][8] ;
 wire \fifo.fifo[6][9] ;
 wire \fifo.fifo[7][0] ;
 wire \fifo.fifo[7][10] ;
 wire \fifo.fifo[7][11] ;
 wire \fifo.fifo[7][12] ;
 wire \fifo.fifo[7][13] ;
 wire \fifo.fifo[7][14] ;
 wire \fifo.fifo[7][15] ;
 wire \fifo.fifo[7][16] ;
 wire \fifo.fifo[7][17] ;
 wire \fifo.fifo[7][18] ;
 wire \fifo.fifo[7][19] ;
 wire \fifo.fifo[7][1] ;
 wire \fifo.fifo[7][20] ;
 wire \fifo.fifo[7][21] ;
 wire \fifo.fifo[7][22] ;
 wire \fifo.fifo[7][23] ;
 wire \fifo.fifo[7][24] ;
 wire \fifo.fifo[7][25] ;
 wire \fifo.fifo[7][26] ;
 wire \fifo.fifo[7][27] ;
 wire \fifo.fifo[7][28] ;
 wire \fifo.fifo[7][29] ;
 wire \fifo.fifo[7][2] ;
 wire \fifo.fifo[7][30] ;
 wire \fifo.fifo[7][31] ;
 wire \fifo.fifo[7][32] ;
 wire \fifo.fifo[7][33] ;
 wire \fifo.fifo[7][34] ;
 wire \fifo.fifo[7][35] ;
 wire \fifo.fifo[7][36] ;
 wire \fifo.fifo[7][37] ;
 wire \fifo.fifo[7][38] ;
 wire \fifo.fifo[7][39] ;
 wire \fifo.fifo[7][3] ;
 wire \fifo.fifo[7][40] ;
 wire \fifo.fifo[7][41] ;
 wire \fifo.fifo[7][42] ;
 wire \fifo.fifo[7][43] ;
 wire \fifo.fifo[7][44] ;
 wire \fifo.fifo[7][45] ;
 wire \fifo.fifo[7][46] ;
 wire \fifo.fifo[7][47] ;
 wire \fifo.fifo[7][48] ;
 wire \fifo.fifo[7][49] ;
 wire \fifo.fifo[7][4] ;
 wire \fifo.fifo[7][50] ;
 wire \fifo.fifo[7][51] ;
 wire \fifo.fifo[7][52] ;
 wire \fifo.fifo[7][53] ;
 wire \fifo.fifo[7][54] ;
 wire \fifo.fifo[7][55] ;
 wire \fifo.fifo[7][5] ;
 wire \fifo.fifo[7][6] ;
 wire \fifo.fifo[7][7] ;
 wire \fifo.fifo[7][8] ;
 wire \fifo.fifo[7][9] ;
 wire \fifo.fifo_empty ;
 wire \fifo.rd_data[0] ;
 wire \fifo.rd_data[10] ;
 wire \fifo.rd_data[11] ;
 wire \fifo.rd_data[12] ;
 wire \fifo.rd_data[13] ;
 wire \fifo.rd_data[14] ;
 wire \fifo.rd_data[15] ;
 wire \fifo.rd_data[16] ;
 wire \fifo.rd_data[17] ;
 wire \fifo.rd_data[18] ;
 wire \fifo.rd_data[19] ;
 wire \fifo.rd_data[1] ;
 wire \fifo.rd_data[20] ;
 wire \fifo.rd_data[21] ;
 wire \fifo.rd_data[22] ;
 wire \fifo.rd_data[23] ;
 wire \fifo.rd_data[24] ;
 wire \fifo.rd_data[25] ;
 wire \fifo.rd_data[26] ;
 wire \fifo.rd_data[27] ;
 wire \fifo.rd_data[28] ;
 wire \fifo.rd_data[29] ;
 wire \fifo.rd_data[2] ;
 wire \fifo.rd_data[30] ;
 wire \fifo.rd_data[31] ;
 wire \fifo.rd_data[32] ;
 wire \fifo.rd_data[33] ;
 wire \fifo.rd_data[34] ;
 wire \fifo.rd_data[35] ;
 wire \fifo.rd_data[36] ;
 wire \fifo.rd_data[37] ;
 wire \fifo.rd_data[38] ;
 wire \fifo.rd_data[39] ;
 wire \fifo.rd_data[3] ;
 wire \fifo.rd_data[40] ;
 wire \fifo.rd_data[41] ;
 wire \fifo.rd_data[42] ;
 wire \fifo.rd_data[43] ;
 wire \fifo.rd_data[44] ;
 wire \fifo.rd_data[45] ;
 wire \fifo.rd_data[46] ;
 wire \fifo.rd_data[47] ;
 wire \fifo.rd_data[48] ;
 wire \fifo.rd_data[49] ;
 wire \fifo.rd_data[4] ;
 wire \fifo.rd_data[50] ;
 wire \fifo.rd_data[51] ;
 wire \fifo.rd_data[52] ;
 wire \fifo.rd_data[53] ;
 wire \fifo.rd_data[54] ;
 wire \fifo.rd_data[55] ;
 wire \fifo.rd_data[5] ;
 wire \fifo.rd_data[6] ;
 wire \fifo.rd_data[7] ;
 wire \fifo.rd_data[8] ;
 wire \fifo.rd_data[9] ;
 wire \fifo.rd_ptr[0] ;
 wire \fifo.rd_ptr[1] ;
 wire \fifo.rd_ptr[2] ;
 wire \fifo.wr_ptr[0] ;
 wire \fifo.wr_ptr[1] ;
 wire \fifo.wr_ptr[2] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \u0.E[10] ;
 wire \u0.E[11] ;
 wire \u0.E[12] ;
 wire \u0.E[15] ;
 wire \u0.E[16] ;
 wire \u0.E[17] ;
 wire \u0.E[18] ;
 wire \u0.E[1] ;
 wire \u0.E[21] ;
 wire \u0.E[22] ;
 wire \u0.E[23] ;
 wire \u0.E[24] ;
 wire \u0.E[27] ;
 wire \u0.E[28] ;
 wire \u0.E[29] ;
 wire \u0.E[2] ;
 wire \u0.E[30] ;
 wire \u0.E[33] ;
 wire \u0.E[34] ;
 wire \u0.E[35] ;
 wire \u0.E[36] ;
 wire \u0.E[39] ;
 wire \u0.E[3] ;
 wire \u0.E[40] ;
 wire \u0.E[41] ;
 wire \u0.E[42] ;
 wire \u0.E[45] ;
 wire \u0.E[46] ;
 wire \u0.E[4] ;
 wire \u0.E[5] ;
 wire \u0.E[6] ;
 wire \u0.E[9] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\u0.E[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_0818_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\fifo.wr_ptr[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_1936_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_1936_));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_8 _2945_ (.A(\counter_inst.count[3] ),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_4 _2946_ (.A(\counter_inst.count[1] ),
    .X(_0659_));
 sky130_fd_sc_hd__clkbuf_4 _2947_ (.A(\counter_inst.count[0] ),
    .X(_0660_));
 sky130_fd_sc_hd__nand4_1 _2948_ (.A(_0658_),
    .B(\counter_inst.count[2] ),
    .C(_0659_),
    .D(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__or2_1 _2949_ (.A(\counter_inst.count[4] ),
    .B(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__nand2_1 _2950_ (.A(net653),
    .B(_0661_),
    .Y(_0663_));
 sky130_fd_sc_hd__a21oi_1 _2951_ (.A1(_0662_),
    .A2(_0663_),
    .B1(net66),
    .Y(_0622_));
 sky130_fd_sc_hd__a31o_1 _2952_ (.A1(\counter_inst.count[2] ),
    .A2(_0659_),
    .A3(_0660_),
    .B1(_0658_),
    .X(_0664_));
 sky130_fd_sc_hd__and3b_1 _2953_ (.A_N(net66),
    .B(_0661_),
    .C(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__clkbuf_1 _2954_ (.A(_0665_),
    .X(_0621_));
 sky130_fd_sc_hd__a21oi_1 _2955_ (.A1(_0659_),
    .A2(_0660_),
    .B1(\counter_inst.count[2] ),
    .Y(_0666_));
 sky130_fd_sc_hd__a31o_1 _2956_ (.A1(\counter_inst.count[2] ),
    .A2(_0659_),
    .A3(_0660_),
    .B1(net66),
    .X(_0667_));
 sky130_fd_sc_hd__nor2_1 _2957_ (.A(_0666_),
    .B(_0667_),
    .Y(_0620_));
 sky130_fd_sc_hd__xnor2_1 _2958_ (.A(_0659_),
    .B(_0660_),
    .Y(_0668_));
 sky130_fd_sc_hd__nor2_1 _2959_ (.A(net66),
    .B(_0668_),
    .Y(_0619_));
 sky130_fd_sc_hd__nor2b_1 _2960_ (.A(net66),
    .B_N(_0662_),
    .Y(_0669_));
 sky130_fd_sc_hd__buf_4 _2961_ (.A(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__xor2_2 _2962_ (.A(\counter_inst.count[3] ),
    .B(_0660_),
    .X(_0671_));
 sky130_fd_sc_hd__xor2_2 _2963_ (.A(_0658_),
    .B(_0659_),
    .X(_0672_));
 sky130_fd_sc_hd__nor2_1 _2964_ (.A(_0671_),
    .B(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__clkbuf_4 _2965_ (.A(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__nor2_1 _2966_ (.A(_0658_),
    .B(\counter_inst.count[2] ),
    .Y(_0675_));
 sky130_fd_sc_hd__and3_1 _2967_ (.A(\counter_inst.count[4] ),
    .B(_0674_),
    .C(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__a211oi_1 _2968_ (.A1(_0670_),
    .A2(_0676_),
    .B1(_0660_),
    .C1(net66),
    .Y(_0618_));
 sky130_fd_sc_hd__buf_4 _2969_ (.A(_0670_),
    .X(_0677_));
 sky130_fd_sc_hd__nor2_1 _2970_ (.A(net66),
    .B(_0662_),
    .Y(_0678_));
 sky130_fd_sc_hd__buf_4 _2971_ (.A(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__a31o_1 _2972_ (.A1(net188),
    .A2(_0677_),
    .A3(_0676_),
    .B1(_0679_),
    .X(_0617_));
 sky130_fd_sc_hd__inv_2 _2973_ (.A(\fifo.wr_ptr[0] ),
    .Y(_0680_));
 sky130_fd_sc_hd__or4_1 _2974_ (.A(net15),
    .B(net14),
    .C(net17),
    .D(net16),
    .X(_0681_));
 sky130_fd_sc_hd__or4_1 _2975_ (.A(net10),
    .B(net9),
    .C(net12),
    .D(net11),
    .X(_0682_));
 sky130_fd_sc_hd__or4_1 _2976_ (.A(net19),
    .B(net18),
    .C(net21),
    .D(net20),
    .X(_0683_));
 sky130_fd_sc_hd__or4_1 _2977_ (.A(net23),
    .B(net22),
    .C(net26),
    .D(net25),
    .X(_0684_));
 sky130_fd_sc_hd__or4_1 _2978_ (.A(_0681_),
    .B(_0682_),
    .C(_0683_),
    .D(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__or4_1 _2979_ (.A(net57),
    .B(net46),
    .C(net63),
    .D(net62),
    .X(_0686_));
 sky130_fd_sc_hd__or4_1 _2980_ (.A(net13),
    .B(net2),
    .C(net35),
    .D(net24),
    .X(_0687_));
 sky130_fd_sc_hd__or4_1 _2981_ (.A(net65),
    .B(net64),
    .C(net4),
    .D(net3),
    .X(_0688_));
 sky130_fd_sc_hd__or4_1 _2982_ (.A(net6),
    .B(net5),
    .C(net8),
    .D(net7),
    .X(_0689_));
 sky130_fd_sc_hd__or4_1 _2983_ (.A(_0686_),
    .B(_0687_),
    .C(_0688_),
    .D(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__or4_1 _2984_ (.A(net32),
    .B(net31),
    .C(net34),
    .D(net33),
    .X(_0691_));
 sky130_fd_sc_hd__or4_2 _2985_ (.A(net28),
    .B(net27),
    .C(net30),
    .D(net29),
    .X(_0692_));
 sky130_fd_sc_hd__or4_1 _2986_ (.A(net37),
    .B(net36),
    .C(net39),
    .D(net38),
    .X(_0693_));
 sky130_fd_sc_hd__or4_2 _2987_ (.A(net41),
    .B(net40),
    .C(net43),
    .D(net42),
    .X(_0694_));
 sky130_fd_sc_hd__or4_2 _2988_ (.A(_0691_),
    .B(_0692_),
    .C(_0693_),
    .D(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__or4_2 _2989_ (.A(net50),
    .B(net49),
    .C(net52),
    .D(net51),
    .X(_0696_));
 sky130_fd_sc_hd__or4_1 _2990_ (.A(net45),
    .B(net44),
    .C(net48),
    .D(net47),
    .X(_0697_));
 sky130_fd_sc_hd__or4_1 _2991_ (.A(net54),
    .B(net53),
    .C(net56),
    .D(net55),
    .X(_0698_));
 sky130_fd_sc_hd__or4_1 _2992_ (.A(net59),
    .B(net58),
    .C(net61),
    .D(net60),
    .X(_0699_));
 sky130_fd_sc_hd__or4_2 _2993_ (.A(_0696_),
    .B(_0697_),
    .C(_0698_),
    .D(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__or4_4 _2994_ (.A(_0685_),
    .B(_0690_),
    .C(_0695_),
    .D(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__clkbuf_4 _2995_ (.A(net118),
    .X(_0702_));
 sky130_fd_sc_hd__clkbuf_4 _2996_ (.A(net111),
    .X(_0703_));
 sky130_fd_sc_hd__or4b_1 _2997_ (.A(_0702_),
    .B(_0703_),
    .C(net120),
    .D_N(net119),
    .X(_0704_));
 sky130_fd_sc_hd__clkbuf_4 _2998_ (.A(net100),
    .X(_0705_));
 sky130_fd_sc_hd__or4b_1 _2999_ (.A(net78),
    .B(_0705_),
    .C(net89),
    .D_N(net67),
    .X(_0706_));
 sky130_fd_sc_hd__or2_4 _3000_ (.A(_0704_),
    .B(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__buf_4 _3001_ (.A(net70),
    .X(_0708_));
 sky130_fd_sc_hd__clkbuf_4 _3002_ (.A(net73),
    .X(_0709_));
 sky130_fd_sc_hd__clkbuf_4 _3003_ (.A(net72),
    .X(_0710_));
 sky130_fd_sc_hd__buf_4 _3004_ (.A(net71),
    .X(_0711_));
 sky130_fd_sc_hd__and4bb_1 _3005_ (.A_N(_0708_),
    .B_N(_0709_),
    .C(_0710_),
    .D(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__clkbuf_4 _3006_ (.A(net121),
    .X(_0713_));
 sky130_fd_sc_hd__buf_2 _3007_ (.A(net122),
    .X(_0714_));
 sky130_fd_sc_hd__buf_4 _3008_ (.A(net69),
    .X(_0715_));
 sky130_fd_sc_hd__and4b_1 _3009_ (.A_N(_0713_),
    .B(_0714_),
    .C(net68),
    .D(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__nand2_2 _3010_ (.A(_0712_),
    .B(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__clkbuf_4 _3011_ (.A(net75),
    .X(_0718_));
 sky130_fd_sc_hd__clkbuf_4 _3012_ (.A(net77),
    .X(_0719_));
 sky130_fd_sc_hd__or4b_1 _3013_ (.A(_0718_),
    .B(_0719_),
    .C(net76),
    .D_N(net74),
    .X(_0720_));
 sky130_fd_sc_hd__clkbuf_4 _3014_ (.A(net79),
    .X(_0721_));
 sky130_fd_sc_hd__clkbuf_4 _3015_ (.A(net82),
    .X(_0722_));
 sky130_fd_sc_hd__clkbuf_4 _3016_ (.A(net81),
    .X(_0723_));
 sky130_fd_sc_hd__clkbuf_4 _3017_ (.A(net80),
    .X(_0724_));
 sky130_fd_sc_hd__or4bb_1 _3018_ (.A(_0721_),
    .B(_0722_),
    .C_N(_0723_),
    .D_N(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__or4_1 _3019_ (.A(_0707_),
    .B(_0717_),
    .C(_0720_),
    .D(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__buf_2 _3020_ (.A(net108),
    .X(_0727_));
 sky130_fd_sc_hd__inv_2 _3021_ (.A(net107),
    .Y(_0728_));
 sky130_fd_sc_hd__clkbuf_4 _3022_ (.A(net105),
    .X(_0729_));
 sky130_fd_sc_hd__clkbuf_4 _3023_ (.A(net106),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_1 _3024_ (.A(_0729_),
    .B(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__clkbuf_4 _3025_ (.A(net104),
    .X(_0732_));
 sky130_fd_sc_hd__clkbuf_4 _3026_ (.A(net103),
    .X(_0733_));
 sky130_fd_sc_hd__buf_2 _3027_ (.A(net102),
    .X(_0734_));
 sky130_fd_sc_hd__or4b_1 _3028_ (.A(net101),
    .B(_0732_),
    .C(_0733_),
    .D_N(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__or4_1 _3029_ (.A(_0727_),
    .B(_0728_),
    .C(_0731_),
    .D(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__clkbuf_4 _3030_ (.A(net110),
    .X(_0737_));
 sky130_fd_sc_hd__clkbuf_4 _3031_ (.A(net109),
    .X(_0738_));
 sky130_fd_sc_hd__buf_2 _3032_ (.A(net113),
    .X(_0739_));
 sky130_fd_sc_hd__or4b_1 _3033_ (.A(_0737_),
    .B(_0738_),
    .C(_0739_),
    .D_N(net112),
    .X(_0740_));
 sky130_fd_sc_hd__buf_2 _3034_ (.A(net115),
    .X(_0741_));
 sky130_fd_sc_hd__buf_2 _3035_ (.A(net116),
    .X(_0742_));
 sky130_fd_sc_hd__buf_2 _3036_ (.A(net114),
    .X(_0743_));
 sky130_fd_sc_hd__or4bb_1 _3037_ (.A(_0741_),
    .B(net117),
    .C_N(_0742_),
    .D_N(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__or3_1 _3038_ (.A(_0736_),
    .B(_0740_),
    .C(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__clkbuf_4 _3039_ (.A(net87),
    .X(_0746_));
 sky130_fd_sc_hd__buf_2 _3040_ (.A(net91),
    .X(_0747_));
 sky130_fd_sc_hd__buf_2 _3041_ (.A(net88),
    .X(_0748_));
 sky130_fd_sc_hd__and4bb_1 _3042_ (.A_N(_0746_),
    .B_N(_0747_),
    .C(net90),
    .D(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__clkbuf_4 _3043_ (.A(net83),
    .X(_0750_));
 sky130_fd_sc_hd__clkbuf_4 _3044_ (.A(net85),
    .X(_0751_));
 sky130_fd_sc_hd__clkbuf_4 _3045_ (.A(net84),
    .X(_0752_));
 sky130_fd_sc_hd__and4bb_1 _3046_ (.A_N(_0750_),
    .B_N(_0751_),
    .C(net86),
    .D(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__nand2_1 _3047_ (.A(_0749_),
    .B(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__clkbuf_4 _3048_ (.A(net92),
    .X(_0755_));
 sky130_fd_sc_hd__buf_4 _3049_ (.A(net93),
    .X(_0756_));
 sky130_fd_sc_hd__buf_4 _3050_ (.A(net94),
    .X(_0757_));
 sky130_fd_sc_hd__clkbuf_4 _3051_ (.A(net95),
    .X(_0758_));
 sky130_fd_sc_hd__nand4_1 _3052_ (.A(_0755_),
    .B(_0756_),
    .C(_0757_),
    .D(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__buf_2 _3053_ (.A(net96),
    .X(_0760_));
 sky130_fd_sc_hd__clkbuf_4 _3054_ (.A(net99),
    .X(_0761_));
 sky130_fd_sc_hd__clkbuf_4 _3055_ (.A(net98),
    .X(_0762_));
 sky130_fd_sc_hd__buf_2 _3056_ (.A(net97),
    .X(_0763_));
 sky130_fd_sc_hd__or4bb_1 _3057_ (.A(_0760_),
    .B(_0761_),
    .C_N(_0762_),
    .D_N(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__or3_1 _3058_ (.A(_0754_),
    .B(_0759_),
    .C(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__or4_4 _3059_ (.A(_0701_),
    .B(_0726_),
    .C(_0745_),
    .D(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__inv_2 _3060_ (.A(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__or3b_1 _3061_ (.A(_0659_),
    .B(net1),
    .C_N(_0660_),
    .X(_0768_));
 sky130_fd_sc_hd__or4b_4 _3062_ (.A(\counter_inst.count[4] ),
    .B(_0767_),
    .C(_0768_),
    .D_N(_0675_),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_1 _3063_ (.A(_0680_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__nand2_1 _3064_ (.A(\fifo.wr_ptr[1] ),
    .B(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__inv_2 _3065_ (.A(\fifo.wr_ptr[2] ),
    .Y(_0772_));
 sky130_fd_sc_hd__and3_1 _3066_ (.A(_0772_),
    .B(\fifo.wr_ptr[1] ),
    .C(_0770_),
    .X(_0773_));
 sky130_fd_sc_hd__buf_6 _3067_ (.A(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__a21o_1 _3068_ (.A1(\fifo.wr_ptr[2] ),
    .A2(_0771_),
    .B1(_0774_),
    .X(_0616_));
 sky130_fd_sc_hd__or2_1 _3069_ (.A(\fifo.wr_ptr[1] ),
    .B(_0770_),
    .X(_0775_));
 sky130_fd_sc_hd__and2_1 _3070_ (.A(_0771_),
    .B(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__clkbuf_1 _3071_ (.A(_0776_),
    .X(_0615_));
 sky130_fd_sc_hd__nor2_1 _3072_ (.A(\fifo.wr_ptr[0] ),
    .B(_0769_),
    .Y(_0777_));
 sky130_fd_sc_hd__and2_1 _3073_ (.A(\fifo.wr_ptr[0] ),
    .B(_0769_),
    .X(_0778_));
 sky130_fd_sc_hd__or2_1 _3074_ (.A(_0777_),
    .B(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__clkbuf_1 _3075_ (.A(_0779_),
    .X(_0614_));
 sky130_fd_sc_hd__inv_2 _3076_ (.A(\fifo.rd_ptr[2] ),
    .Y(_0780_));
 sky130_fd_sc_hd__buf_4 _3077_ (.A(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__buf_4 _3078_ (.A(\fifo.rd_ptr[1] ),
    .X(_0782_));
 sky130_fd_sc_hd__inv_2 _3079_ (.A(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__buf_6 _3080_ (.A(\fifo.rd_ptr[0] ),
    .X(_0784_));
 sky130_fd_sc_hd__buf_4 _3081_ (.A(_0784_),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_1 _3082_ (.A(_0680_),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__o221a_1 _3083_ (.A1(_0772_),
    .A2(\fifo.rd_ptr[2] ),
    .B1(_0783_),
    .B2(\fifo.wr_ptr[1] ),
    .C1(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__inv_2 _3084_ (.A(\fifo.wr_ptr[1] ),
    .Y(_0788_));
 sky130_fd_sc_hd__buf_4 _3085_ (.A(\fifo.rd_ptr[1] ),
    .X(_0789_));
 sky130_fd_sc_hd__o22a_1 _3086_ (.A1(_0788_),
    .A2(_0789_),
    .B1(_0785_),
    .B2(_0680_),
    .X(_0790_));
 sky130_fd_sc_hd__o2111a_1 _3087_ (.A1(\fifo.wr_ptr[2] ),
    .A2(_0781_),
    .B1(_0787_),
    .C1(_0790_),
    .D1(_0658_),
    .X(_0791_));
 sky130_fd_sc_hd__nor3b_1 _3088_ (.A(\counter_inst.count[4] ),
    .B(_0660_),
    .C_N(_0659_),
    .Y(_0792_));
 sky130_fd_sc_hd__and3_1 _3089_ (.A(_0658_),
    .B(\counter_inst.count[2] ),
    .C(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__a21bo_1 _3090_ (.A1(_0767_),
    .A2(_0793_),
    .B1_N(_0769_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2_1 _3091_ (.A0(\fifo.fifo_empty ),
    .A1(_0791_),
    .S(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__clkbuf_1 _3092_ (.A(_0795_),
    .X(_0613_));
 sky130_fd_sc_hd__or4b_1 _3093_ (.A(\counter_inst.count[4] ),
    .B(_0671_),
    .C(_0672_),
    .D_N(_0675_),
    .X(_0796_));
 sky130_fd_sc_hd__clkbuf_4 _3094_ (.A(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__buf_4 _3095_ (.A(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _3096_ (.A0(net61),
    .A1(\R[8] ),
    .S(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__buf_4 _3097_ (.A(_0799_),
    .X(\u0.E[11] ));
 sky130_fd_sc_hd__and2_1 _3098_ (.A(_0678_),
    .B(_0766_),
    .X(_0800_));
 sky130_fd_sc_hd__clkbuf_4 _3099_ (.A(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__a22o_1 _3100_ (.A1(net183),
    .A2(_0677_),
    .B1(\u0.E[11] ),
    .B2(_0801_),
    .X(_0612_));
 sky130_fd_sc_hd__xnor2_1 _3101_ (.A(_0658_),
    .B(_0660_),
    .Y(_0802_));
 sky130_fd_sc_hd__xnor2_1 _3102_ (.A(_0658_),
    .B(_0659_),
    .Y(_0803_));
 sky130_fd_sc_hd__xnor2_4 _3103_ (.A(_0658_),
    .B(\counter_inst.count[2] ),
    .Y(_0804_));
 sky130_fd_sc_hd__and3_1 _3104_ (.A(_0802_),
    .B(_0803_),
    .C(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__clkbuf_4 _3105_ (.A(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__clkbuf_4 _3106_ (.A(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__buf_6 _3107_ (.A(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__xnor2_1 _3108_ (.A(\counter_inst.count[3] ),
    .B(net1),
    .Y(_0809_));
 sky130_fd_sc_hd__buf_2 _3109_ (.A(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__clkbuf_4 _3110_ (.A(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__or2_2 _3111_ (.A(net88),
    .B(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__xor2_2 _3112_ (.A(\counter_inst.count[3] ),
    .B(net1),
    .X(_0813_));
 sky130_fd_sc_hd__clkbuf_4 _3113_ (.A(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__clkbuf_8 _3114_ (.A(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__or2_4 _3115_ (.A(net96),
    .B(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__and3_1 _3116_ (.A(_0671_),
    .B(_0803_),
    .C(_0804_),
    .X(_0817_));
 sky130_fd_sc_hd__clkbuf_4 _3117_ (.A(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__clkbuf_4 _3118_ (.A(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__clkbuf_2 _3119_ (.A(_0813_),
    .X(_0820_));
 sky130_fd_sc_hd__or2_2 _3120_ (.A(net104),
    .B(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__or2_2 _3121_ (.A(net81),
    .B(_0810_),
    .X(_0822_));
 sky130_fd_sc_hd__xor2_2 _3122_ (.A(_0658_),
    .B(\counter_inst.count[2] ),
    .X(_0823_));
 sky130_fd_sc_hd__and3_1 _3123_ (.A(_0671_),
    .B(_0803_),
    .C(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__clkbuf_4 _3124_ (.A(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__clkbuf_4 _3125_ (.A(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__or2_2 _3126_ (.A(net105),
    .B(_0820_),
    .X(_0827_));
 sky130_fd_sc_hd__or2_2 _3127_ (.A(net80),
    .B(_0810_),
    .X(_0828_));
 sky130_fd_sc_hd__and3_1 _3128_ (.A(_0826_),
    .B(_0827_),
    .C(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__and3_1 _3129_ (.A(_0671_),
    .B(_0672_),
    .C(_0804_),
    .X(_0830_));
 sky130_fd_sc_hd__clkbuf_4 _3130_ (.A(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__buf_4 _3131_ (.A(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__buf_2 _3132_ (.A(_0809_),
    .X(_0833_));
 sky130_fd_sc_hd__clkbuf_4 _3133_ (.A(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__or2_2 _3134_ (.A(net110),
    .B(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__clkbuf_4 _3135_ (.A(_0820_),
    .X(_0836_));
 sky130_fd_sc_hd__or2_1 _3136_ (.A(net74),
    .B(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__and3_1 _3137_ (.A(_0832_),
    .B(_0835_),
    .C(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__a311o_1 _3138_ (.A1(_0819_),
    .A2(_0821_),
    .A3(_0822_),
    .B1(_0829_),
    .C1(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__and3_1 _3139_ (.A(_0802_),
    .B(_0672_),
    .C(_0804_),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_4 _3140_ (.A(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__clkbuf_4 _3141_ (.A(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__clkbuf_4 _3142_ (.A(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__or2_1 _3143_ (.A(net121),
    .B(_0833_),
    .X(_0844_));
 sky130_fd_sc_hd__clkbuf_4 _3144_ (.A(net89),
    .X(_0845_));
 sky130_fd_sc_hd__or2_2 _3145_ (.A(_0845_),
    .B(_0836_),
    .X(_0846_));
 sky130_fd_sc_hd__clkbuf_4 _3146_ (.A(net120),
    .X(_0847_));
 sky130_fd_sc_hd__clkbuf_4 _3147_ (.A(_0811_),
    .X(_0848_));
 sky130_fd_sc_hd__clkbuf_4 _3148_ (.A(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__and3_1 _3149_ (.A(_0802_),
    .B(_0672_),
    .C(_0823_),
    .X(_0850_));
 sky130_fd_sc_hd__buf_4 _3150_ (.A(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__clkbuf_4 _3151_ (.A(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__clkbuf_4 _3152_ (.A(_0852_),
    .X(_0853_));
 sky130_fd_sc_hd__or2_2 _3153_ (.A(net91),
    .B(_0836_),
    .X(_0854_));
 sky130_fd_sc_hd__o211a_1 _3154_ (.A1(_0847_),
    .A2(_0849_),
    .B1(_0853_),
    .C1(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__a31o_1 _3155_ (.A1(_0843_),
    .A2(_0844_),
    .A3(_0846_),
    .B1(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__clkbuf_4 _3156_ (.A(net90),
    .X(_0857_));
 sky130_fd_sc_hd__clkbuf_4 _3157_ (.A(_0815_),
    .X(_0858_));
 sky130_fd_sc_hd__clkbuf_4 _3158_ (.A(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__and3_4 _3159_ (.A(_0802_),
    .B(_0803_),
    .C(_0823_),
    .X(_0860_));
 sky130_fd_sc_hd__clkbuf_4 _3160_ (.A(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_4 _3161_ (.A(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__or2_2 _3162_ (.A(net95),
    .B(_0810_),
    .X(_0863_));
 sky130_fd_sc_hd__o211a_1 _3163_ (.A1(_0857_),
    .A2(_0859_),
    .B1(_0862_),
    .C1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__and3_1 _3164_ (.A(_0671_),
    .B(_0672_),
    .C(_0823_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_4 _3165_ (.A(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__clkbuf_4 _3166_ (.A(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__clkbuf_4 _3167_ (.A(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__or2_2 _3168_ (.A(net114),
    .B(_0810_),
    .X(_0869_));
 sky130_fd_sc_hd__or2_1 _3169_ (.A(net106),
    .B(_0820_),
    .X(_0870_));
 sky130_fd_sc_hd__and3_1 _3170_ (.A(_0868_),
    .B(_0869_),
    .C(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__or4_2 _3171_ (.A(_0839_),
    .B(_0856_),
    .C(_0864_),
    .D(_0871_),
    .X(_0872_));
 sky130_fd_sc_hd__a31oi_4 _3172_ (.A1(_0808_),
    .A2(_0812_),
    .A3(_0816_),
    .B1(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(net59),
    .A1(\R[16] ),
    .S(_0797_),
    .X(_0874_));
 sky130_fd_sc_hd__clkbuf_8 _3174_ (.A(_0874_),
    .X(\u0.E[23] ));
 sky130_fd_sc_hd__xnor2_4 _3175_ (.A(_0873_),
    .B(\u0.E[23] ),
    .Y(_0875_));
 sky130_fd_sc_hd__clkbuf_4 _3176_ (.A(_0673_),
    .X(_0876_));
 sky130_fd_sc_hd__clkbuf_4 _3177_ (.A(_0804_),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_2 _3178_ (.A(_0876_),
    .B(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__buf_4 _3179_ (.A(_0878_),
    .X(_0879_));
 sky130_fd_sc_hd__clkbuf_4 _3180_ (.A(net74),
    .X(_0880_));
 sky130_fd_sc_hd__or2_2 _3181_ (.A(_0722_),
    .B(_0836_),
    .X(_0881_));
 sky130_fd_sc_hd__o21a_1 _3182_ (.A1(_0880_),
    .A2(_0849_),
    .B1(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__or2_1 _3183_ (.A(_0879_),
    .B(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__or2_2 _3184_ (.A(net72),
    .B(_0820_),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(net67),
    .A1(_0713_),
    .S(_0815_),
    .X(_0885_));
 sky130_fd_sc_hd__a32o_1 _3186_ (.A1(_0835_),
    .A2(_0852_),
    .A3(_0884_),
    .B1(_0885_),
    .B2(_0826_),
    .X(_0886_));
 sky130_fd_sc_hd__or2_2 _3187_ (.A(net87),
    .B(_0820_),
    .X(_0887_));
 sky130_fd_sc_hd__clkbuf_8 _3188_ (.A(_0833_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(_0714_),
    .A1(net90),
    .S(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_4 _3190_ (.A(_0817_),
    .X(_0890_));
 sky130_fd_sc_hd__clkbuf_4 _3191_ (.A(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__a32o_1 _3192_ (.A1(_0863_),
    .A2(_0867_),
    .A3(_0887_),
    .B1(_0889_),
    .B2(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__buf_4 _3193_ (.A(_0840_),
    .X(_0893_));
 sky130_fd_sc_hd__clkbuf_4 _3194_ (.A(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__or2_2 _3195_ (.A(net112),
    .B(_0833_),
    .X(_0895_));
 sky130_fd_sc_hd__clkbuf_4 _3196_ (.A(_0813_),
    .X(_0896_));
 sky130_fd_sc_hd__buf_4 _3197_ (.A(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(_0747_),
    .A1(_0760_),
    .S(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__buf_4 _3199_ (.A(_0831_),
    .X(_0899_));
 sky130_fd_sc_hd__a32o_1 _3200_ (.A1(_0827_),
    .A2(_0894_),
    .A3(_0895_),
    .B1(_0898_),
    .B2(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__clkbuf_4 _3201_ (.A(_0877_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(_0723_),
    .A1(_0730_),
    .S(_0848_),
    .X(_0902_));
 sky130_fd_sc_hd__o21a_1 _3203_ (.A1(_0901_),
    .A2(_0902_),
    .B1(_0674_),
    .X(_0903_));
 sky130_fd_sc_hd__or4_2 _3204_ (.A(_0886_),
    .B(_0892_),
    .C(_0900_),
    .D(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__buf_6 _3205_ (.A(_0798_),
    .X(_0905_));
 sky130_fd_sc_hd__clkbuf_8 _3206_ (.A(_0797_),
    .X(_0906_));
 sky130_fd_sc_hd__or2b_1 _3207_ (.A(\R[20] ),
    .B_N(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__o21ai_4 _3208_ (.A1(net21),
    .A2(_0905_),
    .B1(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__a21o_2 _3209_ (.A1(_0883_),
    .A2(_0904_),
    .B1(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__nand3_4 _3210_ (.A(_0883_),
    .B(_0904_),
    .C(_0908_),
    .Y(_0910_));
 sky130_fd_sc_hd__mux2_1 _3211_ (.A0(_0845_),
    .A1(net120),
    .S(_0897_),
    .X(_0911_));
 sky130_fd_sc_hd__o21a_1 _3212_ (.A1(_0901_),
    .A2(_0911_),
    .B1(_0674_),
    .X(_0912_));
 sky130_fd_sc_hd__clkbuf_4 _3213_ (.A(_0831_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _3214_ (.A0(net88),
    .A1(_0758_),
    .S(_0897_),
    .X(_0914_));
 sky130_fd_sc_hd__a32o_1 _3215_ (.A1(_0913_),
    .A2(_0821_),
    .A3(_0828_),
    .B1(_0894_),
    .B2(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__or2_2 _3216_ (.A(net113),
    .B(_0810_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _3217_ (.A0(_0709_),
    .A1(_0737_),
    .S(_0897_),
    .X(_0917_));
 sky130_fd_sc_hd__clkbuf_4 _3218_ (.A(_0890_),
    .X(_0918_));
 sky130_fd_sc_hd__a32o_1 _3219_ (.A1(_0827_),
    .A2(_0867_),
    .A3(_0916_),
    .B1(_0917_),
    .B2(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__buf_4 _3220_ (.A(_0825_),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _3221_ (.A0(net90),
    .A1(net98),
    .S(_0897_),
    .X(_0921_));
 sky130_fd_sc_hd__a32o_1 _3222_ (.A1(_0837_),
    .A2(_0920_),
    .A3(_0869_),
    .B1(_0921_),
    .B2(_0852_),
    .X(_0922_));
 sky130_fd_sc_hd__or4_2 _3223_ (.A(_0912_),
    .B(_0915_),
    .C(_0919_),
    .D(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__clkbuf_4 _3224_ (.A(_0813_),
    .X(_0924_));
 sky130_fd_sc_hd__clkbuf_4 _3225_ (.A(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__or2_2 _3226_ (.A(net121),
    .B(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__buf_2 _3227_ (.A(_0810_),
    .X(_0927_));
 sky130_fd_sc_hd__or2_2 _3228_ (.A(net78),
    .B(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__a21o_1 _3229_ (.A1(_0926_),
    .A2(_0928_),
    .B1(_0879_),
    .X(_0929_));
 sky130_fd_sc_hd__buf_4 _3230_ (.A(_0797_),
    .X(_0930_));
 sky130_fd_sc_hd__or2b_1 _3231_ (.A(net730),
    .B_N(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__o21ai_4 _3232_ (.A1(net12),
    .A2(_0905_),
    .B1(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__a21oi_2 _3233_ (.A1(_0923_),
    .A2(_0929_),
    .B1(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__and3_1 _3234_ (.A(_0923_),
    .B(_0929_),
    .C(_0932_),
    .X(_0934_));
 sky130_fd_sc_hd__a211o_1 _3235_ (.A1(_0909_),
    .A2(_0910_),
    .B1(_0933_),
    .C1(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__nand2_4 _3236_ (.A(_0909_),
    .B(_0910_),
    .Y(_0936_));
 sky130_fd_sc_hd__or2_2 _3237_ (.A(net103),
    .B(_0820_),
    .X(_0937_));
 sky130_fd_sc_hd__or2_2 _3238_ (.A(net73),
    .B(_0924_),
    .X(_0938_));
 sky130_fd_sc_hd__and3_1 _3239_ (.A(_0860_),
    .B(_0916_),
    .C(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__clkbuf_4 _3240_ (.A(_0820_),
    .X(_0940_));
 sky130_fd_sc_hd__or2_2 _3241_ (.A(net88),
    .B(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__or2_2 _3242_ (.A(net97),
    .B(_0888_),
    .X(_0942_));
 sky130_fd_sc_hd__clkbuf_4 _3243_ (.A(net78),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(_0943_),
    .A1(net98),
    .S(_0897_),
    .X(_0944_));
 sky130_fd_sc_hd__a32o_1 _3245_ (.A1(_0920_),
    .A2(_0941_),
    .A3(_0942_),
    .B1(_0944_),
    .B2(_0913_),
    .X(_0945_));
 sky130_fd_sc_hd__a311o_1 _3246_ (.A1(_0842_),
    .A2(_0869_),
    .A3(_0937_),
    .B1(_0939_),
    .C1(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_4 _3247_ (.A(_0851_),
    .X(_0947_));
 sky130_fd_sc_hd__or2_2 _3248_ (.A(net82),
    .B(_0833_),
    .X(_0948_));
 sky130_fd_sc_hd__o211a_1 _3249_ (.A1(net120),
    .A2(_0848_),
    .B1(_0918_),
    .C1(_0887_),
    .X(_0949_));
 sky130_fd_sc_hd__or2_2 _3250_ (.A(net122),
    .B(_0834_),
    .X(_0950_));
 sky130_fd_sc_hd__a31o_1 _3251_ (.A1(_0846_),
    .A2(_0867_),
    .A3(_0950_),
    .B1(_0806_),
    .X(_0951_));
 sky130_fd_sc_hd__a311o_1 _3252_ (.A1(_0821_),
    .A2(_0947_),
    .A3(_0948_),
    .B1(_0949_),
    .C1(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__or2_4 _3253_ (.A(_0724_),
    .B(_0925_),
    .X(_0953_));
 sky130_fd_sc_hd__or2_4 _3254_ (.A(_0710_),
    .B(_0888_),
    .X(_0954_));
 sky130_fd_sc_hd__buf_4 _3255_ (.A(_0878_),
    .X(_0955_));
 sky130_fd_sc_hd__a21o_1 _3256_ (.A1(_0953_),
    .A2(_0954_),
    .B1(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__o21a_2 _3257_ (.A1(_0946_),
    .A2(_0952_),
    .B1(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _3258_ (.A0(net4),
    .A1(\R[18] ),
    .S(_0906_),
    .X(_0958_));
 sky130_fd_sc_hd__buf_2 _3259_ (.A(_0958_),
    .X(\u0.E[27] ));
 sky130_fd_sc_hd__xor2_4 _3260_ (.A(_0957_),
    .B(\u0.E[27] ),
    .X(_0959_));
 sky130_fd_sc_hd__xor2_2 _3261_ (.A(_0936_),
    .B(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__or2_4 _3262_ (.A(net89),
    .B(_0834_),
    .X(_0961_));
 sky130_fd_sc_hd__or2_2 _3263_ (.A(net95),
    .B(_0814_),
    .X(_0962_));
 sky130_fd_sc_hd__or2_2 _3264_ (.A(_0732_),
    .B(_0888_),
    .X(_0963_));
 sky130_fd_sc_hd__and3_1 _3265_ (.A(_0826_),
    .B(_0962_),
    .C(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__or2_2 _3266_ (.A(_0743_),
    .B(_0940_),
    .X(_0965_));
 sky130_fd_sc_hd__or2_2 _3267_ (.A(net90),
    .B(_0834_),
    .X(_0966_));
 sky130_fd_sc_hd__and3_1 _3268_ (.A(_0842_),
    .B(_0965_),
    .C(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__a311o_1 _3269_ (.A1(_0862_),
    .A2(_0961_),
    .A3(_0953_),
    .B1(_0964_),
    .C1(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__buf_2 _3270_ (.A(_0810_),
    .X(_0969_));
 sky130_fd_sc_hd__or2_2 _3271_ (.A(_0729_),
    .B(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__or2_2 _3272_ (.A(net98),
    .B(_0940_),
    .X(_0971_));
 sky130_fd_sc_hd__or2_2 _3273_ (.A(net110),
    .B(_0814_),
    .X(_0972_));
 sky130_fd_sc_hd__and3_1 _3274_ (.A(_0947_),
    .B(_0812_),
    .C(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__clkbuf_4 _3275_ (.A(_0866_),
    .X(_0974_));
 sky130_fd_sc_hd__or2_2 _3276_ (.A(net73),
    .B(_0811_),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _3277_ (.A0(net120),
    .A1(net74),
    .S(_0815_),
    .X(_0976_));
 sky130_fd_sc_hd__a32o_1 _3278_ (.A1(_0974_),
    .A2(_0926_),
    .A3(_0975_),
    .B1(_0976_),
    .B2(_0832_),
    .X(_0977_));
 sky130_fd_sc_hd__a311o_1 _3279_ (.A1(_0819_),
    .A2(_0970_),
    .A3(_0971_),
    .B1(_0973_),
    .C1(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__and3_1 _3280_ (.A(_0854_),
    .B(_0807_),
    .C(_0916_),
    .X(_0979_));
 sky130_fd_sc_hd__nor3_4 _3281_ (.A(_0968_),
    .B(_0978_),
    .C(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__mux2_1 _3282_ (.A0(net35),
    .A1(\R[17] ),
    .S(_0905_),
    .X(_0981_));
 sky130_fd_sc_hd__buf_8 _3283_ (.A(_0981_),
    .X(\u0.E[24] ));
 sky130_fd_sc_hd__xnor2_4 _3284_ (.A(_0980_),
    .B(\u0.E[24] ),
    .Y(_0982_));
 sky130_fd_sc_hd__buf_2 _3285_ (.A(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__a21oi_1 _3286_ (.A1(_0935_),
    .A2(_0960_),
    .B1(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__xor2_4 _3287_ (.A(_0980_),
    .B(\u0.E[24] ),
    .X(_0985_));
 sky130_fd_sc_hd__o211a_1 _3288_ (.A1(_0933_),
    .A2(_0934_),
    .B1(_0909_),
    .C1(_0910_),
    .X(_0986_));
 sky130_fd_sc_hd__nor2_1 _3289_ (.A(_0985_),
    .B(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__buf_4 _3290_ (.A(_0810_),
    .X(_0988_));
 sky130_fd_sc_hd__or2_4 _3291_ (.A(net106),
    .B(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_4 _3292_ (.A(_0826_),
    .X(_0990_));
 sky130_fd_sc_hd__or2_2 _3293_ (.A(net78),
    .B(_0820_),
    .X(_0991_));
 sky130_fd_sc_hd__clkbuf_4 _3294_ (.A(_0899_),
    .X(_0992_));
 sky130_fd_sc_hd__or2_2 _3295_ (.A(net67),
    .B(_0820_),
    .X(_0993_));
 sky130_fd_sc_hd__o211a_1 _3296_ (.A1(_0762_),
    .A2(_0849_),
    .B1(_0891_),
    .C1(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__a31o_1 _3297_ (.A1(_0992_),
    .A2(_0887_),
    .A3(_0942_),
    .B1(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__or2_1 _3298_ (.A(net96),
    .B(_0833_),
    .X(_0996_));
 sky130_fd_sc_hd__and3_1 _3299_ (.A(_0974_),
    .B(_0941_),
    .C(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__and3_1 _3300_ (.A(_0861_),
    .B(_0948_),
    .C(_0937_),
    .X(_0998_));
 sky130_fd_sc_hd__and3_1 _3301_ (.A(_0947_),
    .B(_0938_),
    .C(_0895_),
    .X(_0999_));
 sky130_fd_sc_hd__and3_1 _3302_ (.A(_0894_),
    .B(_0916_),
    .C(_0884_),
    .X(_1000_));
 sky130_fd_sc_hd__or4_1 _3303_ (.A(_0997_),
    .B(_0998_),
    .C(_0999_),
    .D(_1000_),
    .X(_1001_));
 sky130_fd_sc_hd__a311o_1 _3304_ (.A1(_0990_),
    .A2(_0950_),
    .A3(_0991_),
    .B1(_0995_),
    .C1(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__a31oi_4 _3305_ (.A1(_0808_),
    .A2(_0965_),
    .A3(_0989_),
    .B1(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__mux2_1 _3306_ (.A0(net30),
    .A1(net720),
    .S(_0930_),
    .X(_1004_));
 sky130_fd_sc_hd__clkbuf_8 _3307_ (.A(_1004_),
    .X(\u0.E[30] ));
 sky130_fd_sc_hd__xor2_4 _3308_ (.A(_1003_),
    .B(\u0.E[30] ),
    .X(_1005_));
 sky130_fd_sc_hd__a21o_1 _3309_ (.A1(_0960_),
    .A2(_0987_),
    .B1(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__a21o_1 _3310_ (.A1(_0923_),
    .A2(_0929_),
    .B1(_0932_),
    .X(_1007_));
 sky130_fd_sc_hd__nand3_2 _3311_ (.A(_0923_),
    .B(_0929_),
    .C(_0932_),
    .Y(_1008_));
 sky130_fd_sc_hd__nand2_2 _3312_ (.A(_1007_),
    .B(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__clkbuf_4 _3313_ (.A(_0959_),
    .X(_1010_));
 sky130_fd_sc_hd__nor2_1 _3314_ (.A(_1009_),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__or3_1 _3315_ (.A(_0983_),
    .B(_0986_),
    .C(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__nand3_1 _3316_ (.A(_1009_),
    .B(_0936_),
    .C(_0959_),
    .Y(_1013_));
 sky130_fd_sc_hd__a211o_1 _3317_ (.A1(_1009_),
    .A2(_0936_),
    .B1(_1010_),
    .C1(_0985_),
    .X(_1014_));
 sky130_fd_sc_hd__and3_1 _3318_ (.A(_1005_),
    .B(_1013_),
    .C(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a2bb2o_1 _3319_ (.A1_N(_0984_),
    .A2_N(_1006_),
    .B1(_1012_),
    .B2(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__o211ai_2 _3320_ (.A1(_0933_),
    .A2(_0934_),
    .B1(_0909_),
    .C1(_0910_),
    .Y(_1017_));
 sky130_fd_sc_hd__and2_1 _3321_ (.A(_0935_),
    .B(_1017_),
    .X(_1018_));
 sky130_fd_sc_hd__xnor2_4 _3322_ (.A(_1003_),
    .B(\u0.E[30] ),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_1 _3323_ (.A(_0982_),
    .B(_0935_),
    .Y(_1020_));
 sky130_fd_sc_hd__a211o_1 _3324_ (.A1(_0983_),
    .A2(_1018_),
    .B1(_1019_),
    .C1(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__nor2_1 _3325_ (.A(_1010_),
    .B(_0986_),
    .Y(_1022_));
 sky130_fd_sc_hd__or3_1 _3326_ (.A(_0982_),
    .B(_1005_),
    .C(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__a22o_1 _3327_ (.A1(_1010_),
    .A2(_0986_),
    .B1(_1021_),
    .B2(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__and3_1 _3328_ (.A(_0935_),
    .B(_0959_),
    .C(_1017_),
    .X(_1025_));
 sky130_fd_sc_hd__o21ai_1 _3329_ (.A1(_1011_),
    .A2(_1025_),
    .B1(_0982_),
    .Y(_1026_));
 sky130_fd_sc_hd__or2_1 _3330_ (.A(_1005_),
    .B(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__a21oi_1 _3331_ (.A1(_1024_),
    .A2(_1027_),
    .B1(_0875_),
    .Y(_1028_));
 sky130_fd_sc_hd__a21o_1 _3332_ (.A1(_0875_),
    .A2(_1016_),
    .B1(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__clkbuf_8 _3333_ (.A(_0905_),
    .X(_1030_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(net60),
    .A1(net257),
    .S(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__xnor2_1 _3335_ (.A(_1029_),
    .B(_1031_),
    .Y(\FP[8] ));
 sky130_fd_sc_hd__a22o_1 _3336_ (.A1(net182),
    .A2(_0677_),
    .B1(_0801_),
    .B2(\FP[8] ),
    .X(_0611_));
 sky130_fd_sc_hd__a22o_1 _3337_ (.A1(net181),
    .A2(_0677_),
    .B1(_0801_),
    .B2(\u0.E[23] ),
    .X(_0610_));
 sky130_fd_sc_hd__nand2_4 _3338_ (.A(_0728_),
    .B(_0836_),
    .Y(_1032_));
 sky130_fd_sc_hd__or2_2 _3339_ (.A(net115),
    .B(_0896_),
    .X(_1033_));
 sky130_fd_sc_hd__or2_4 _3340_ (.A(net70),
    .B(_0927_),
    .X(_1034_));
 sky130_fd_sc_hd__clkbuf_4 _3341_ (.A(_0924_),
    .X(_1035_));
 sky130_fd_sc_hd__or2_4 _3342_ (.A(net118),
    .B(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__or2_2 _3343_ (.A(net94),
    .B(_0940_),
    .X(_1037_));
 sky130_fd_sc_hd__buf_2 _3344_ (.A(net101),
    .X(_1038_));
 sky130_fd_sc_hd__or2_4 _3345_ (.A(_1038_),
    .B(_0888_),
    .X(_1039_));
 sky130_fd_sc_hd__and3_1 _3346_ (.A(_0990_),
    .B(_1037_),
    .C(_1039_),
    .X(_1040_));
 sky130_fd_sc_hd__or2_2 _3347_ (.A(net100),
    .B(_0940_),
    .X(_1041_));
 sky130_fd_sc_hd__or2_2 _3348_ (.A(_0761_),
    .B(_0834_),
    .X(_1042_));
 sky130_fd_sc_hd__and3_1 _3349_ (.A(_0819_),
    .B(_1041_),
    .C(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__a311o_1 _3350_ (.A1(_0868_),
    .A2(_1034_),
    .A3(_1036_),
    .B1(_1040_),
    .C1(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__or2_2 _3351_ (.A(net75),
    .B(_0940_),
    .X(_1045_));
 sky130_fd_sc_hd__or2_1 _3352_ (.A(_0752_),
    .B(_0848_),
    .X(_1046_));
 sky130_fd_sc_hd__and3_1 _3353_ (.A(_0843_),
    .B(_1045_),
    .C(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__buf_4 _3354_ (.A(net119),
    .X(_1048_));
 sky130_fd_sc_hd__or2_2 _3355_ (.A(_0715_),
    .B(_0969_),
    .X(_1049_));
 sky130_fd_sc_hd__o211a_1 _3356_ (.A1(_1048_),
    .A2(_0859_),
    .B1(_1049_),
    .C1(_0992_),
    .X(_1050_));
 sky130_fd_sc_hd__or2_2 _3357_ (.A(_0751_),
    .B(_0888_),
    .X(_1051_));
 sky130_fd_sc_hd__or2_2 _3358_ (.A(net109),
    .B(_0836_),
    .X(_1052_));
 sky130_fd_sc_hd__or2_2 _3359_ (.A(net79),
    .B(_0925_),
    .X(_1053_));
 sky130_fd_sc_hd__or2_2 _3360_ (.A(_0742_),
    .B(_0848_),
    .X(_1054_));
 sky130_fd_sc_hd__and3_1 _3361_ (.A(_0861_),
    .B(_1053_),
    .C(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__a31o_1 _3362_ (.A1(_0853_),
    .A2(_1051_),
    .A3(_1052_),
    .B1(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__or4_1 _3363_ (.A(_1044_),
    .B(_1047_),
    .C(_1050_),
    .D(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__a31o_2 _3364_ (.A1(_0808_),
    .A2(_1032_),
    .A3(_1033_),
    .B1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__xnor2_4 _3365_ (.A(\u0.E[11] ),
    .B(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__or2_2 _3366_ (.A(net68),
    .B(_0988_),
    .X(_1060_));
 sky130_fd_sc_hd__a21o_1 _3367_ (.A1(_1045_),
    .A2(_1060_),
    .B1(_0955_),
    .X(_1061_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(net76),
    .A1(net102),
    .S(_0988_),
    .X(_1062_));
 sky130_fd_sc_hd__o21a_1 _3369_ (.A1(_0877_),
    .A2(_1062_),
    .B1(_0876_),
    .X(_1063_));
 sky130_fd_sc_hd__or2_2 _3370_ (.A(net71),
    .B(_0814_),
    .X(_1064_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(net86),
    .A1(net92),
    .S(_0925_),
    .X(_1065_));
 sky130_fd_sc_hd__a32o_1 _3372_ (.A1(_0893_),
    .A2(_1032_),
    .A3(_1064_),
    .B1(_1065_),
    .B2(_0831_),
    .X(_1066_));
 sky130_fd_sc_hd__or2_2 _3373_ (.A(net85),
    .B(_1035_),
    .X(_1067_));
 sky130_fd_sc_hd__or2_2 _3374_ (.A(_0756_),
    .B(_0969_),
    .X(_1068_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(net100),
    .A1(net83),
    .S(_0811_),
    .X(_1069_));
 sky130_fd_sc_hd__a32o_1 _3376_ (.A1(_0866_),
    .A2(_1067_),
    .A3(_1068_),
    .B1(_1069_),
    .B2(_0890_),
    .X(_1070_));
 sky130_fd_sc_hd__or2_2 _3377_ (.A(net70),
    .B(_0814_),
    .X(_1071_));
 sky130_fd_sc_hd__or2_2 _3378_ (.A(net108),
    .B(_0927_),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _3379_ (.A0(_0703_),
    .A1(net117),
    .S(_0988_),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_4 _3380_ (.A(_0824_),
    .X(_1074_));
 sky130_fd_sc_hd__a32o_1 _3381_ (.A1(_0851_),
    .A2(_1071_),
    .A3(_1072_),
    .B1(_1073_),
    .B2(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__or4_2 _3382_ (.A(_1063_),
    .B(_1066_),
    .C(_1070_),
    .D(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__or2b_1 _3383_ (.A(\R[12] ),
    .B_N(_0798_),
    .X(_1077_));
 sky130_fd_sc_hd__o21ai_4 _3384_ (.A1(net23),
    .A2(_0906_),
    .B1(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__a21o_1 _3385_ (.A1(_1061_),
    .A2(_1076_),
    .B1(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__nand3_2 _3386_ (.A(_1061_),
    .B(_1076_),
    .C(_1078_),
    .Y(_1080_));
 sky130_fd_sc_hd__nand2_4 _3387_ (.A(_1079_),
    .B(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__or2_2 _3388_ (.A(net86),
    .B(_0988_),
    .X(_1082_));
 sky130_fd_sc_hd__a21o_1 _3389_ (.A1(_1037_),
    .A2(_1082_),
    .B1(_0955_),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _3390_ (.A0(net100),
    .A1(net85),
    .S(_0969_),
    .X(_1084_));
 sky130_fd_sc_hd__o21a_1 _3391_ (.A1(_0877_),
    .A2(_1084_),
    .B1(_0876_),
    .X(_1085_));
 sky130_fd_sc_hd__or2_2 _3392_ (.A(net75),
    .B(_0969_),
    .X(_1086_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(net119),
    .A1(net117),
    .S(_0811_),
    .X(_1087_));
 sky130_fd_sc_hd__a32o_1 _3394_ (.A1(_0831_),
    .A2(_1071_),
    .A3(_1086_),
    .B1(_1087_),
    .B2(_0841_),
    .X(_1088_));
 sky130_fd_sc_hd__clkbuf_4 _3395_ (.A(_0865_),
    .X(_1089_));
 sky130_fd_sc_hd__or2_2 _3396_ (.A(net76),
    .B(_0833_),
    .X(_1090_));
 sky130_fd_sc_hd__or2_2 _3397_ (.A(net69),
    .B(_0896_),
    .X(_1091_));
 sky130_fd_sc_hd__mux2_1 _3398_ (.A0(net79),
    .A1(net102),
    .S(_0811_),
    .X(_1092_));
 sky130_fd_sc_hd__a32o_1 _3399_ (.A1(_1089_),
    .A2(_1090_),
    .A3(_1091_),
    .B1(_1092_),
    .B2(_0818_),
    .X(_1093_));
 sky130_fd_sc_hd__or2_2 _3400_ (.A(net101),
    .B(_0814_),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_1 _3401_ (.A0(net92),
    .A1(net116),
    .S(_0988_),
    .X(_1095_));
 sky130_fd_sc_hd__clkbuf_4 _3402_ (.A(_0850_),
    .X(_1096_));
 sky130_fd_sc_hd__a32o_1 _3403_ (.A1(_1074_),
    .A2(_1032_),
    .A3(_1094_),
    .B1(_1095_),
    .B2(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__or4_2 _3404_ (.A(_1085_),
    .B(_1088_),
    .C(_1093_),
    .D(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__or2b_1 _3405_ (.A(\R[11] ),
    .B_N(_0930_),
    .X(_1099_));
 sky130_fd_sc_hd__o21ai_4 _3406_ (.A1(net15),
    .A2(_0905_),
    .B1(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__a21o_1 _3407_ (.A1(_1083_),
    .A2(_1098_),
    .B1(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__nand3_2 _3408_ (.A(_1083_),
    .B(_1098_),
    .C(_1100_),
    .Y(_1102_));
 sky130_fd_sc_hd__and2_2 _3409_ (.A(_1101_),
    .B(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__o211a_1 _3410_ (.A1(net119),
    .A2(_0815_),
    .B1(_1074_),
    .C1(_1034_),
    .X(_1104_));
 sky130_fd_sc_hd__or2_2 _3411_ (.A(net102),
    .B(_0811_),
    .X(_1105_));
 sky130_fd_sc_hd__and3_1 _3412_ (.A(_1089_),
    .B(_1037_),
    .C(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__a311o_1 _3413_ (.A1(_0832_),
    .A2(_1041_),
    .A3(_1039_),
    .B1(_1104_),
    .C1(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__or2_4 _3414_ (.A(net117),
    .B(_0833_),
    .X(_1108_));
 sky130_fd_sc_hd__mux2_1 _3415_ (.A0(net107),
    .A1(net116),
    .S(_1035_),
    .X(_1109_));
 sky130_fd_sc_hd__a32o_1 _3416_ (.A1(_1096_),
    .A2(_1108_),
    .A3(_1053_),
    .B1(_1109_),
    .B2(_0841_),
    .X(_1110_));
 sky130_fd_sc_hd__or2_2 _3417_ (.A(net92),
    .B(_0896_),
    .X(_1111_));
 sky130_fd_sc_hd__and3_1 _3418_ (.A(_0818_),
    .B(_1049_),
    .C(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__a311o_1 _3419_ (.A1(_0861_),
    .A2(_1045_),
    .A3(_1051_),
    .B1(_1110_),
    .C1(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__or2_2 _3420_ (.A(net84),
    .B(_0896_),
    .X(_1114_));
 sky130_fd_sc_hd__and3_1 _3421_ (.A(_0806_),
    .B(_1114_),
    .C(_1090_),
    .X(_1115_));
 sky130_fd_sc_hd__nor3_4 _3422_ (.A(_1107_),
    .B(_1113_),
    .C(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__mux2_1 _3423_ (.A0(net57),
    .A1(\R[9] ),
    .S(_0930_),
    .X(_1117_));
 sky130_fd_sc_hd__buf_4 _3424_ (.A(_1117_),
    .X(\u0.E[12] ));
 sky130_fd_sc_hd__xor2_4 _3425_ (.A(_1116_),
    .B(\u0.E[12] ),
    .X(_1118_));
 sky130_fd_sc_hd__a21o_1 _3426_ (.A1(_1081_),
    .A2(_1103_),
    .B1(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__or2_2 _3427_ (.A(net109),
    .B(_0833_),
    .X(_1120_));
 sky130_fd_sc_hd__or2_2 _3428_ (.A(net116),
    .B(_1035_),
    .X(_1121_));
 sky130_fd_sc_hd__or2_1 _3429_ (.A(net118),
    .B(_0969_),
    .X(_1122_));
 sky130_fd_sc_hd__and3_1 _3430_ (.A(_0841_),
    .B(_1121_),
    .C(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__a31o_1 _3431_ (.A1(_0899_),
    .A2(_1091_),
    .A3(_1120_),
    .B1(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__or2_2 _3432_ (.A(net77),
    .B(_0927_),
    .X(_1125_));
 sky130_fd_sc_hd__o211a_1 _3433_ (.A1(net68),
    .A2(_0815_),
    .B1(_1089_),
    .C1(_1086_),
    .X(_1126_));
 sky130_fd_sc_hd__a31o_1 _3434_ (.A1(_0891_),
    .A2(_1094_),
    .A3(_1125_),
    .B1(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__or2_2 _3435_ (.A(net79),
    .B(_0927_),
    .X(_1128_));
 sky130_fd_sc_hd__or2_2 _3436_ (.A(net99),
    .B(_0814_),
    .X(_1129_));
 sky130_fd_sc_hd__or2_2 _3437_ (.A(net119),
    .B(_0927_),
    .X(_1130_));
 sky130_fd_sc_hd__a31o_1 _3438_ (.A1(_0851_),
    .A2(_1130_),
    .A3(_1033_),
    .B1(_0806_),
    .X(_1131_));
 sky130_fd_sc_hd__or2_2 _3439_ (.A(net94),
    .B(_0811_),
    .X(_1132_));
 sky130_fd_sc_hd__and3_1 _3440_ (.A(_0860_),
    .B(_1114_),
    .C(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__a311o_1 _3441_ (.A1(_0826_),
    .A2(_1128_),
    .A3(_1129_),
    .B1(_1131_),
    .C1(_1133_),
    .X(_1134_));
 sky130_fd_sc_hd__or2_2 _3442_ (.A(net93),
    .B(_0896_),
    .X(_1135_));
 sky130_fd_sc_hd__a21o_1 _3443_ (.A1(_1051_),
    .A2(_1135_),
    .B1(_0955_),
    .X(_1136_));
 sky130_fd_sc_hd__o31a_4 _3444_ (.A1(_1124_),
    .A2(_1127_),
    .A3(_1134_),
    .B1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_1 _3445_ (.A0(net6),
    .A1(\R[10] ),
    .S(_0930_),
    .X(_1138_));
 sky130_fd_sc_hd__buf_4 _3446_ (.A(_1138_),
    .X(\u0.E[15] ));
 sky130_fd_sc_hd__xor2_4 _3447_ (.A(_1137_),
    .B(\u0.E[15] ),
    .X(_1139_));
 sky130_fd_sc_hd__nor2_1 _3448_ (.A(_1081_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__xnor2_4 _3449_ (.A(_1116_),
    .B(\u0.E[12] ),
    .Y(_1141_));
 sky130_fd_sc_hd__xnor2_4 _3450_ (.A(_1137_),
    .B(\u0.E[15] ),
    .Y(_1142_));
 sky130_fd_sc_hd__nor2_1 _3451_ (.A(_1081_),
    .B(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__a22o_1 _3452_ (.A1(_1079_),
    .A2(_1080_),
    .B1(_1101_),
    .B2(_1102_),
    .X(_1144_));
 sky130_fd_sc_hd__or3b_1 _3453_ (.A(_1141_),
    .B(_1143_),
    .C_N(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__o21a_1 _3454_ (.A1(_1119_),
    .A2(_1140_),
    .B1(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__nor2_1 _3455_ (.A(_1103_),
    .B(_1139_),
    .Y(_1147_));
 sky130_fd_sc_hd__o211ai_1 _3456_ (.A1(_1119_),
    .A2(_1147_),
    .B1(_1059_),
    .C1(_1145_),
    .Y(_1148_));
 sky130_fd_sc_hd__o21ai_1 _3457_ (.A1(_1059_),
    .A2(_1146_),
    .B1(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__xnor2_2 _3458_ (.A(_1081_),
    .B(_1139_),
    .Y(_1150_));
 sky130_fd_sc_hd__nand2_2 _3459_ (.A(_1101_),
    .B(_1102_),
    .Y(_1151_));
 sky130_fd_sc_hd__nor2_1 _3460_ (.A(_1151_),
    .B(_1139_),
    .Y(_1152_));
 sky130_fd_sc_hd__or2_1 _3461_ (.A(_1150_),
    .B(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__nand2_1 _3462_ (.A(_1118_),
    .B(_1103_),
    .Y(_1154_));
 sky130_fd_sc_hd__mux2_1 _3463_ (.A0(_1143_),
    .A1(_1153_),
    .S(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__nand4_2 _3464_ (.A(_1079_),
    .B(_1080_),
    .C(_1101_),
    .D(_1102_),
    .Y(_1156_));
 sky130_fd_sc_hd__a21oi_2 _3465_ (.A1(_1144_),
    .A2(_1156_),
    .B1(_1142_),
    .Y(_1157_));
 sky130_fd_sc_hd__a21o_1 _3466_ (.A1(_1151_),
    .A2(_1142_),
    .B1(_1141_),
    .X(_1158_));
 sky130_fd_sc_hd__nor2_1 _3467_ (.A(_1157_),
    .B(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__o21ai_1 _3468_ (.A1(_1147_),
    .A2(_1143_),
    .B1(_1141_),
    .Y(_1160_));
 sky130_fd_sc_hd__nand2_1 _3469_ (.A(_1059_),
    .B(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__o22a_1 _3470_ (.A1(_1059_),
    .A2(_1155_),
    .B1(_1159_),
    .B2(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__and3_1 _3471_ (.A(_1074_),
    .B(_1091_),
    .C(_1086_),
    .X(_1163_));
 sky130_fd_sc_hd__and3_1 _3472_ (.A(_0818_),
    .B(_1071_),
    .C(_1120_),
    .X(_1164_));
 sky130_fd_sc_hd__a311o_1 _3473_ (.A1(_0832_),
    .A2(_1128_),
    .A3(_1094_),
    .B1(_1163_),
    .C1(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__and3_1 _3474_ (.A(_0974_),
    .B(_1032_),
    .C(_1129_),
    .X(_1166_));
 sky130_fd_sc_hd__and3_1 _3475_ (.A(_0861_),
    .B(_1130_),
    .C(_1121_),
    .X(_1167_));
 sky130_fd_sc_hd__or2_1 _3476_ (.A(net100),
    .B(_0927_),
    .X(_1168_));
 sky130_fd_sc_hd__and3_1 _3477_ (.A(_0852_),
    .B(_1114_),
    .C(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__a31o_1 _3478_ (.A1(_0842_),
    .A2(_1067_),
    .A3(_1132_),
    .B1(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__or4_1 _3479_ (.A(_1165_),
    .B(_1166_),
    .C(_1167_),
    .D(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__a31o_2 _3480_ (.A1(_0807_),
    .A2(_1108_),
    .A3(_1036_),
    .B1(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__mux2_1 _3481_ (.A0(net32),
    .A1(\R[13] ),
    .S(_0798_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_4 _3482_ (.A(_1173_),
    .X(\u0.E[18] ));
 sky130_fd_sc_hd__xor2_4 _3483_ (.A(_1172_),
    .B(\u0.E[18] ),
    .X(_1174_));
 sky130_fd_sc_hd__mux2_1 _3484_ (.A0(_1149_),
    .A1(_1162_),
    .S(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__mux2_1 _3485_ (.A0(net58),
    .A1(\L[16] ),
    .S(_1030_),
    .X(_1176_));
 sky130_fd_sc_hd__xor2_2 _3486_ (.A(_1175_),
    .B(_1176_),
    .X(\FP[16] ));
 sky130_fd_sc_hd__a22o_1 _3487_ (.A1(net180),
    .A2(_0677_),
    .B1(_0801_),
    .B2(\FP[16] ),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(net56),
    .A1(net189),
    .S(_0797_),
    .X(_1177_));
 sky130_fd_sc_hd__buf_4 _3489_ (.A(_1177_),
    .X(\u0.E[35] ));
 sky130_fd_sc_hd__a22o_1 _3490_ (.A1(net178),
    .A2(_0677_),
    .B1(_0801_),
    .B2(\u0.E[35] ),
    .X(_0608_));
 sky130_fd_sc_hd__and3_1 _3491_ (.A(_1142_),
    .B(_1144_),
    .C(_1156_),
    .X(_1178_));
 sky130_fd_sc_hd__nor2_1 _3492_ (.A(_1103_),
    .B(_1142_),
    .Y(_1179_));
 sky130_fd_sc_hd__or3_2 _3493_ (.A(_1118_),
    .B(_1157_),
    .C(_1178_),
    .X(_1180_));
 sky130_fd_sc_hd__o31a_1 _3494_ (.A1(_1141_),
    .A2(_1178_),
    .A3(_1179_),
    .B1(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__or3_1 _3495_ (.A(_1081_),
    .B(_1103_),
    .C(_1142_),
    .X(_1182_));
 sky130_fd_sc_hd__or3b_1 _3496_ (.A(_1140_),
    .B(_1158_),
    .C_N(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__nand2_1 _3497_ (.A(_1180_),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__a21o_1 _3498_ (.A1(_1144_),
    .A2(_1156_),
    .B1(_1141_),
    .X(_1185_));
 sky130_fd_sc_hd__nand2_1 _3499_ (.A(_1180_),
    .B(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__or2_1 _3500_ (.A(_1139_),
    .B(_1156_),
    .X(_1187_));
 sky130_fd_sc_hd__and2b_1 _3501_ (.A_N(_1119_),
    .B(_1150_),
    .X(_1188_));
 sky130_fd_sc_hd__a31o_1 _3502_ (.A1(_1118_),
    .A2(_1144_),
    .A3(_1187_),
    .B1(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__mux4_1 _3503_ (.A0(_1181_),
    .A1(_1184_),
    .A2(_1186_),
    .A3(_1189_),
    .S0(_1059_),
    .S1(_1174_),
    .X(_1190_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(net55),
    .A1(\L[24] ),
    .S(_1030_),
    .X(_1191_));
 sky130_fd_sc_hd__xnor2_1 _3505_ (.A(_1190_),
    .B(_1191_),
    .Y(\FP[24] ));
 sky130_fd_sc_hd__a22o_1 _3506_ (.A1(net690),
    .A2(_0677_),
    .B1(_0801_),
    .B2(\FP[24] ),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(net54),
    .A1(\R[32] ),
    .S(_0798_),
    .X(_1192_));
 sky130_fd_sc_hd__clkbuf_4 _3508_ (.A(_1192_),
    .X(\u0.E[1] ));
 sky130_fd_sc_hd__a22o_1 _3509_ (.A1(net176),
    .A2(_0677_),
    .B1(_0801_),
    .B2(\u0.E[1] ),
    .X(_0606_));
 sky130_fd_sc_hd__or2_2 _3510_ (.A(net91),
    .B(_0969_),
    .X(_1193_));
 sky130_fd_sc_hd__and3_1 _3511_ (.A(_0826_),
    .B(_0895_),
    .C(_0937_),
    .X(_1194_));
 sky130_fd_sc_hd__and3_1 _3512_ (.A(_0918_),
    .B(_0870_),
    .C(_0916_),
    .X(_1195_));
 sky130_fd_sc_hd__a311o_1 _3513_ (.A1(_0992_),
    .A2(_0884_),
    .A3(_0948_),
    .B1(_1194_),
    .C1(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__and3_1 _3514_ (.A(_0822_),
    .B(_0868_),
    .C(_0938_),
    .X(_1197_));
 sky130_fd_sc_hd__and3_1 _3515_ (.A(_0862_),
    .B(_0950_),
    .C(_0887_),
    .X(_1198_));
 sky130_fd_sc_hd__and3_1 _3516_ (.A(_0947_),
    .B(_0996_),
    .C(_0991_),
    .X(_1199_));
 sky130_fd_sc_hd__a31o_1 _3517_ (.A1(_0843_),
    .A2(_0993_),
    .A3(_0942_),
    .B1(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__or4_1 _3518_ (.A(_1196_),
    .B(_1197_),
    .C(_1198_),
    .D(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__a31o_2 _3519_ (.A1(_0808_),
    .A2(_0971_),
    .A3(_1193_),
    .B1(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__mux2_1 _3520_ (.A0(net28),
    .A1(\R[29] ),
    .S(_0906_),
    .X(_1203_));
 sky130_fd_sc_hd__buf_4 _3521_ (.A(_1203_),
    .X(\u0.E[42] ));
 sky130_fd_sc_hd__xor2_4 _3522_ (.A(_1202_),
    .B(\u0.E[42] ),
    .X(_1204_));
 sky130_fd_sc_hd__inv_2 _3523_ (.A(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__and3_1 _3524_ (.A(_0899_),
    .B(_0870_),
    .C(_0895_),
    .X(_1206_));
 sky130_fd_sc_hd__and3_1 _3525_ (.A(_0891_),
    .B(_0827_),
    .C(_0948_),
    .X(_1207_));
 sky130_fd_sc_hd__a311o_1 _3526_ (.A1(_0842_),
    .A2(_0854_),
    .A3(_0950_),
    .B1(_1206_),
    .C1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__and3_1 _3527_ (.A(_0844_),
    .B(_1096_),
    .C(_0887_),
    .X(_1209_));
 sky130_fd_sc_hd__and3_1 _3528_ (.A(_0835_),
    .B(_1089_),
    .C(_0937_),
    .X(_1210_));
 sky130_fd_sc_hd__and3_1 _3529_ (.A(_0860_),
    .B(_0993_),
    .C(_0996_),
    .X(_1211_));
 sky130_fd_sc_hd__and3_1 _3530_ (.A(_0822_),
    .B(_0920_),
    .C(_0884_),
    .X(_1212_));
 sky130_fd_sc_hd__or4_1 _3531_ (.A(_1209_),
    .B(_1210_),
    .C(_1211_),
    .D(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__or2_2 _3532_ (.A(net97),
    .B(_0925_),
    .X(_1214_));
 sky130_fd_sc_hd__and3_1 _3533_ (.A(_0807_),
    .B(_0966_),
    .C(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__nor3_2 _3534_ (.A(_1208_),
    .B(_1213_),
    .C(_1215_),
    .Y(_1216_));
 sky130_fd_sc_hd__mux2_1 _3535_ (.A0(net13),
    .A1(\R[25] ),
    .S(_0930_),
    .X(_1217_));
 sky130_fd_sc_hd__buf_2 _3536_ (.A(_1217_),
    .X(\u0.E[36] ));
 sky130_fd_sc_hd__xnor2_4 _3537_ (.A(_1216_),
    .B(\u0.E[36] ),
    .Y(_1218_));
 sky130_fd_sc_hd__buf_2 _3538_ (.A(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__or2_2 _3539_ (.A(net122),
    .B(_0925_),
    .X(_1220_));
 sky130_fd_sc_hd__or2_2 _3540_ (.A(net87),
    .B(_0988_),
    .X(_1221_));
 sky130_fd_sc_hd__mux2_1 _3541_ (.A0(net67),
    .A1(net81),
    .S(_0848_),
    .X(_1222_));
 sky130_fd_sc_hd__a32o_1 _3542_ (.A1(_0918_),
    .A2(_0972_),
    .A3(_1221_),
    .B1(_1222_),
    .B2(_0899_),
    .X(_1223_));
 sky130_fd_sc_hd__and3_1 _3543_ (.A(_0974_),
    .B(_0966_),
    .C(_0881_),
    .X(_1224_));
 sky130_fd_sc_hd__a311o_1 _3544_ (.A1(_0853_),
    .A2(_0970_),
    .A3(_1220_),
    .B1(_1223_),
    .C1(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__a21o_1 _3545_ (.A1(_0816_),
    .A2(_0989_),
    .B1(_0901_),
    .X(_1226_));
 sky130_fd_sc_hd__buf_2 _3546_ (.A(net112),
    .X(_1227_));
 sky130_fd_sc_hd__o211a_1 _3547_ (.A1(_1227_),
    .A2(_0858_),
    .B1(_0826_),
    .C1(_1193_),
    .X(_1228_));
 sky130_fd_sc_hd__and3_1 _3548_ (.A(_0894_),
    .B(_0926_),
    .C(_0954_),
    .X(_1229_));
 sky130_fd_sc_hd__a211o_1 _3549_ (.A1(_0674_),
    .A2(_1226_),
    .B1(_1228_),
    .C1(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__a21o_1 _3550_ (.A1(_0863_),
    .A2(_0937_),
    .B1(_0879_),
    .X(_1231_));
 sky130_fd_sc_hd__o21ai_4 _3551_ (.A1(_1225_),
    .A2(_1230_),
    .B1(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(net19),
    .A1(\R[28] ),
    .S(_0906_),
    .X(_1233_));
 sky130_fd_sc_hd__buf_4 _3553_ (.A(_1233_),
    .X(\u0.E[41] ));
 sky130_fd_sc_hd__xnor2_4 _3554_ (.A(_1232_),
    .B(\u0.E[41] ),
    .Y(_1234_));
 sky130_fd_sc_hd__buf_2 _3555_ (.A(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__o211a_1 _3556_ (.A1(net98),
    .A2(_0848_),
    .B1(_0854_),
    .C1(_0867_),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(net120),
    .A1(net90),
    .S(_0834_),
    .X(_1237_));
 sky130_fd_sc_hd__a32o_1 _3558_ (.A1(_0837_),
    .A2(_0828_),
    .A3(_0860_),
    .B1(_1237_),
    .B2(_0920_),
    .X(_1238_));
 sky130_fd_sc_hd__a311o_1 _3559_ (.A1(_0827_),
    .A2(_0947_),
    .A3(_0869_),
    .B1(_1236_),
    .C1(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__and3_1 _3560_ (.A(_0818_),
    .B(_0844_),
    .C(_0941_),
    .X(_1240_));
 sky130_fd_sc_hd__a31o_1 _3561_ (.A1(_0913_),
    .A2(_0846_),
    .A3(_0863_),
    .B1(_0806_),
    .X(_1241_));
 sky130_fd_sc_hd__a311o_1 _3562_ (.A1(_0835_),
    .A2(_0821_),
    .A3(_0842_),
    .B1(_1240_),
    .C1(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__or2_1 _3563_ (.A(net81),
    .B(_0925_),
    .X(_1243_));
 sky130_fd_sc_hd__a21o_1 _3564_ (.A1(_0975_),
    .A2(_1243_),
    .B1(_0955_),
    .X(_1244_));
 sky130_fd_sc_hd__o21a_4 _3565_ (.A1(_1239_),
    .A2(_1242_),
    .B1(_1244_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _3566_ (.A0(net65),
    .A1(\R[26] ),
    .S(_0930_),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_4 _3567_ (.A(_1246_),
    .X(\u0.E[39] ));
 sky130_fd_sc_hd__xor2_4 _3568_ (.A(_1245_),
    .B(\u0.E[39] ),
    .X(_1247_));
 sky130_fd_sc_hd__or2_2 _3569_ (.A(net120),
    .B(_0897_),
    .X(_1248_));
 sky130_fd_sc_hd__and3_1 _3570_ (.A(_0918_),
    .B(_1248_),
    .C(_0989_),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_1 _3571_ (.A0(net121),
    .A1(net74),
    .S(_0815_),
    .X(_1250_));
 sky130_fd_sc_hd__a32o_1 _3572_ (.A1(_0867_),
    .A2(_0816_),
    .A3(_0963_),
    .B1(_1250_),
    .B2(_0826_),
    .X(_1251_));
 sky130_fd_sc_hd__a311o_1 _3573_ (.A1(_0842_),
    .A2(_0953_),
    .A3(_1193_),
    .B1(_1249_),
    .C1(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__a21o_1 _3574_ (.A1(_0966_),
    .A2(_0972_),
    .B1(_0901_),
    .X(_1253_));
 sky130_fd_sc_hd__and3_1 _3575_ (.A(_0852_),
    .B(_0961_),
    .C(_1243_),
    .X(_1254_));
 sky130_fd_sc_hd__and3_1 _3576_ (.A(_0899_),
    .B(_0962_),
    .C(_0970_),
    .X(_1255_));
 sky130_fd_sc_hd__a211o_1 _3577_ (.A1(_0674_),
    .A2(_1253_),
    .B1(_1254_),
    .C1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__a21o_1 _3578_ (.A1(_0869_),
    .A2(_0993_),
    .B1(_0879_),
    .X(_1257_));
 sky130_fd_sc_hd__o21ai_4 _3579_ (.A1(_1252_),
    .A2(_1256_),
    .B1(_1257_),
    .Y(_1258_));
 sky130_fd_sc_hd__mux2_1 _3580_ (.A0(net10),
    .A1(\R[27] ),
    .S(_0906_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_4 _3581_ (.A(_1259_),
    .X(\u0.E[40] ));
 sky130_fd_sc_hd__xor2_4 _3582_ (.A(_1258_),
    .B(\u0.E[40] ),
    .X(_1260_));
 sky130_fd_sc_hd__xnor2_2 _3583_ (.A(_1247_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__xor2_1 _3584_ (.A(_1235_),
    .B(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__xnor2_1 _3585_ (.A(_1234_),
    .B(_1247_),
    .Y(_1263_));
 sky130_fd_sc_hd__or2_1 _3586_ (.A(_1218_),
    .B(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__a21boi_1 _3587_ (.A1(_1219_),
    .A2(_1262_),
    .B1_N(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__xnor2_4 _3588_ (.A(_1245_),
    .B(\u0.E[39] ),
    .Y(_1266_));
 sky130_fd_sc_hd__xnor2_2 _3589_ (.A(_1258_),
    .B(\u0.E[40] ),
    .Y(_1267_));
 sky130_fd_sc_hd__and3b_1 _3590_ (.A_N(_1234_),
    .B(_1266_),
    .C(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__inv_2 _3591_ (.A(_1218_),
    .Y(_1269_));
 sky130_fd_sc_hd__nand2_2 _3592_ (.A(_1234_),
    .B(_1260_),
    .Y(_1270_));
 sky130_fd_sc_hd__or3b_1 _3593_ (.A(_1268_),
    .B(_1269_),
    .C_N(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__o211ai_1 _3594_ (.A1(_1266_),
    .A2(_1260_),
    .B1(_1269_),
    .C1(_1263_),
    .Y(_1272_));
 sky130_fd_sc_hd__a21o_1 _3595_ (.A1(_1271_),
    .A2(_1272_),
    .B1(_1204_),
    .X(_1273_));
 sky130_fd_sc_hd__o21ai_1 _3596_ (.A1(_1205_),
    .A2(_1265_),
    .B1(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__xnor2_1 _3597_ (.A(_1234_),
    .B(_1260_),
    .Y(_1275_));
 sky130_fd_sc_hd__a21o_1 _3598_ (.A1(_1235_),
    .A2(_1266_),
    .B1(_1218_),
    .X(_1276_));
 sky130_fd_sc_hd__nor2_1 _3599_ (.A(_1235_),
    .B(_1260_),
    .Y(_1277_));
 sky130_fd_sc_hd__o2bb2a_1 _3600_ (.A1_N(_1219_),
    .A2_N(_1275_),
    .B1(_1276_),
    .B2(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__o21a_1 _3601_ (.A1(_1235_),
    .A2(_1261_),
    .B1(_1270_),
    .X(_1279_));
 sky130_fd_sc_hd__o21a_1 _3602_ (.A1(_1234_),
    .A2(_1260_),
    .B1(_1247_),
    .X(_1280_));
 sky130_fd_sc_hd__o21ai_1 _3603_ (.A1(_1268_),
    .A2(_1280_),
    .B1(_1218_),
    .Y(_1281_));
 sky130_fd_sc_hd__o211a_1 _3604_ (.A1(_1219_),
    .A2(_1279_),
    .B1(_1281_),
    .C1(_1205_),
    .X(_1282_));
 sky130_fd_sc_hd__a21oi_1 _3605_ (.A1(_1204_),
    .A2(_1278_),
    .B1(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__or2_2 _3606_ (.A(_0739_),
    .B(_0836_),
    .X(_1284_));
 sky130_fd_sc_hd__and3_1 _3607_ (.A(_0992_),
    .B(_0975_),
    .C(_1214_),
    .X(_1285_));
 sky130_fd_sc_hd__a31o_1 _3608_ (.A1(_0862_),
    .A2(_0928_),
    .A3(_1284_),
    .B1(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__and3_1 _3609_ (.A(_0819_),
    .B(_0963_),
    .C(_1220_),
    .X(_1287_));
 sky130_fd_sc_hd__a31o_1 _3610_ (.A1(_0843_),
    .A2(_0812_),
    .A3(_0881_),
    .B1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__or2_2 _3611_ (.A(_0733_),
    .B(_0811_),
    .X(_1289_));
 sky130_fd_sc_hd__and3_1 _3612_ (.A(_0990_),
    .B(_0971_),
    .C(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__a311o_1 _3613_ (.A1(_0868_),
    .A2(_1248_),
    .A3(_0954_),
    .B1(_1288_),
    .C1(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__a311o_2 _3614_ (.A1(_0853_),
    .A2(_0965_),
    .A3(_1221_),
    .B1(_1286_),
    .C1(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__a31oi_4 _3615_ (.A1(_0846_),
    .A2(_0808_),
    .A3(_0895_),
    .B1(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__xnor2_4 _3616_ (.A(\u0.E[35] ),
    .B(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__mux2_2 _3617_ (.A0(_1274_),
    .A1(_1283_),
    .S(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_1 _3618_ (.A0(net53),
    .A1(\L[32] ),
    .S(_1030_),
    .X(_1296_));
 sky130_fd_sc_hd__xnor2_2 _3619_ (.A(_1295_),
    .B(_1296_),
    .Y(\FP[32] ));
 sky130_fd_sc_hd__a22o_1 _3620_ (.A1(net175),
    .A2(_0677_),
    .B1(_0801_),
    .B2(\FP[32] ),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _3621_ (.A0(net52),
    .A1(\R[7] ),
    .S(_0797_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_2 _3622_ (.A(_1297_),
    .X(\u0.E[10] ));
 sky130_fd_sc_hd__or4_1 _3623_ (.A(_0707_),
    .B(_0717_),
    .C(_0720_),
    .D(_0725_),
    .X(_1298_));
 sky130_fd_sc_hd__or3_1 _3624_ (.A(_0736_),
    .B(_0740_),
    .C(_0744_),
    .X(_1299_));
 sky130_fd_sc_hd__or3_1 _3625_ (.A(_0754_),
    .B(_0759_),
    .C(_0764_),
    .X(_1300_));
 sky130_fd_sc_hd__or4_4 _3626_ (.A(_0701_),
    .B(_1298_),
    .C(_1299_),
    .D(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__buf_4 _3627_ (.A(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__buf_4 _3628_ (.A(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _3629_ (.A0(net668),
    .A1(\u0.E[10] ),
    .S(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__a22o_1 _3630_ (.A1(net718),
    .A2(_0677_),
    .B1(_0679_),
    .B2(_1304_),
    .X(_0604_));
 sky130_fd_sc_hd__buf_4 _3631_ (.A(_0678_),
    .X(_1305_));
 sky130_fd_sc_hd__mux2_1 _3632_ (.A0(_1266_),
    .A1(_1280_),
    .S(_1270_),
    .X(_1306_));
 sky130_fd_sc_hd__a21bo_1 _3633_ (.A1(_1269_),
    .A2(_1306_),
    .B1_N(_1271_),
    .X(_1307_));
 sky130_fd_sc_hd__nand2_1 _3634_ (.A(_1266_),
    .B(_1218_),
    .Y(_1308_));
 sky130_fd_sc_hd__a31o_1 _3635_ (.A1(_1266_),
    .A2(_1218_),
    .A3(_1270_),
    .B1(_1204_),
    .X(_1309_));
 sky130_fd_sc_hd__a21oi_1 _3636_ (.A1(_1306_),
    .A2(_1308_),
    .B1(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__a211oi_1 _3637_ (.A1(_1204_),
    .A2(_1307_),
    .B1(_1310_),
    .C1(_1294_),
    .Y(_1311_));
 sky130_fd_sc_hd__o211a_1 _3638_ (.A1(_1219_),
    .A2(_1262_),
    .B1(_1281_),
    .C1(_1204_),
    .X(_1312_));
 sky130_fd_sc_hd__o21a_1 _3639_ (.A1(_1310_),
    .A2(_1312_),
    .B1(_1294_),
    .X(_1313_));
 sky130_fd_sc_hd__mux2_1 _3640_ (.A0(net51),
    .A1(\L[7] ),
    .S(_1030_),
    .X(_1314_));
 sky130_fd_sc_hd__or3_1 _3641_ (.A(_1311_),
    .B(_1313_),
    .C(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__o21ai_1 _3642_ (.A1(_1311_),
    .A2(_1313_),
    .B1(_1314_),
    .Y(_1316_));
 sky130_fd_sc_hd__a21o_1 _3643_ (.A1(_1315_),
    .A2(_1316_),
    .B1(_0767_),
    .X(_1317_));
 sky130_fd_sc_hd__or2_4 _3644_ (.A(\fifo.rd_data[54] ),
    .B(_1303_),
    .X(_1318_));
 sky130_fd_sc_hd__a32o_1 _3645_ (.A1(_1305_),
    .A2(_1317_),
    .A3(_1318_),
    .B1(_0670_),
    .B2(net173),
    .X(_0603_));
 sky130_fd_sc_hd__clkbuf_4 _3646_ (.A(_0670_),
    .X(_1319_));
 sky130_fd_sc_hd__or2b_1 _3647_ (.A(net713),
    .B_N(_0798_),
    .X(_1320_));
 sky130_fd_sc_hd__o21ai_2 _3648_ (.A1(net50),
    .A2(_0906_),
    .B1(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__inv_2 _3649_ (.A(_1321_),
    .Y(\u0.E[22] ));
 sky130_fd_sc_hd__mux2_1 _3650_ (.A0(net275),
    .A1(\u0.E[22] ),
    .S(_1303_),
    .X(_1322_));
 sky130_fd_sc_hd__a22o_1 _3651_ (.A1(net172),
    .A2(_1319_),
    .B1(_0679_),
    .B2(_1322_),
    .X(_0602_));
 sky130_fd_sc_hd__and3_1 _3652_ (.A(_0947_),
    .B(_0971_),
    .C(_0954_),
    .X(_1323_));
 sky130_fd_sc_hd__and3_1 _3653_ (.A(_0899_),
    .B(_0928_),
    .C(_0881_),
    .X(_1324_));
 sky130_fd_sc_hd__a311o_1 _3654_ (.A1(_0990_),
    .A2(_1221_),
    .A3(_1284_),
    .B1(_1323_),
    .C1(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_1 _3655_ (.A0(_0748_),
    .A1(net112),
    .S(_0848_),
    .X(_1326_));
 sky130_fd_sc_hd__a32o_1 _3656_ (.A1(_0861_),
    .A2(_1214_),
    .A3(_1289_),
    .B1(_1326_),
    .B2(_0891_),
    .X(_1327_));
 sky130_fd_sc_hd__o211a_1 _3657_ (.A1(net67),
    .A2(_0849_),
    .B1(_0974_),
    .C1(_0965_),
    .X(_1328_));
 sky130_fd_sc_hd__a311o_1 _3658_ (.A1(_0843_),
    .A2(_0975_),
    .A3(_1220_),
    .B1(_1327_),
    .C1(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__and3_1 _3659_ (.A(_0821_),
    .B(_0807_),
    .C(_0996_),
    .X(_1330_));
 sky130_fd_sc_hd__nor3_4 _3660_ (.A(_1325_),
    .B(_1329_),
    .C(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__xnor2_4 _3661_ (.A(\u0.E[42] ),
    .B(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__buf_2 _3662_ (.A(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__and3_1 _3663_ (.A(_0893_),
    .B(_1221_),
    .C(_1243_),
    .X(_1334_));
 sky130_fd_sc_hd__and3_1 _3664_ (.A(_0890_),
    .B(_0926_),
    .C(_1289_),
    .X(_1335_));
 sky130_fd_sc_hd__and3_1 _3665_ (.A(_0825_),
    .B(_0989_),
    .C(_1220_),
    .X(_1336_));
 sky130_fd_sc_hd__and3_1 _3666_ (.A(_0866_),
    .B(_0970_),
    .C(_1214_),
    .X(_1337_));
 sky130_fd_sc_hd__or4_2 _3667_ (.A(_1334_),
    .B(_1335_),
    .C(_1336_),
    .D(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__mux2_1 _3668_ (.A0(net67),
    .A1(net112),
    .S(_0834_),
    .X(_1339_));
 sky130_fd_sc_hd__o21a_1 _3669_ (.A1(_0877_),
    .A2(_1339_),
    .B1(_0876_),
    .X(_1340_));
 sky130_fd_sc_hd__and3_1 _3670_ (.A(_1096_),
    .B(_0881_),
    .C(_1193_),
    .X(_1341_));
 sky130_fd_sc_hd__a311o_1 _3671_ (.A1(_0832_),
    .A2(_0816_),
    .A3(_0954_),
    .B1(_1340_),
    .C1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__a21o_1 _3672_ (.A1(_0835_),
    .A2(_0991_),
    .B1(_0955_),
    .X(_1343_));
 sky130_fd_sc_hd__o21ai_4 _3673_ (.A1(_1338_),
    .A2(_1342_),
    .B1(_1343_),
    .Y(_1344_));
 sky130_fd_sc_hd__mux2_1 _3674_ (.A0(net45),
    .A1(\R[31] ),
    .S(_0930_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_4 _3675_ (.A(_1345_),
    .X(\u0.E[46] ));
 sky130_fd_sc_hd__xnor2_4 _3676_ (.A(_1344_),
    .B(\u0.E[46] ),
    .Y(_1346_));
 sky130_fd_sc_hd__clkbuf_4 _3677_ (.A(net67),
    .X(_1347_));
 sky130_fd_sc_hd__o21a_1 _3678_ (.A1(_1347_),
    .A2(_0849_),
    .B1(_1248_),
    .X(_1348_));
 sky130_fd_sc_hd__and3_1 _3679_ (.A(_0821_),
    .B(_1089_),
    .C(_0895_),
    .X(_1349_));
 sky130_fd_sc_hd__mux2_2 _3680_ (.A0(_0746_),
    .A1(net98),
    .S(_0940_),
    .X(_1350_));
 sky130_fd_sc_hd__a32o_1 _3681_ (.A1(_0913_),
    .A2(_0916_),
    .A3(_0937_),
    .B1(_1350_),
    .B2(_0894_),
    .X(_1351_));
 sky130_fd_sc_hd__a311o_1 _3682_ (.A1(_0891_),
    .A2(_0869_),
    .A3(_0884_),
    .B1(_1349_),
    .C1(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__a21o_1 _3683_ (.A1(_0991_),
    .A2(_0942_),
    .B1(_0901_),
    .X(_1353_));
 sky130_fd_sc_hd__and3_1 _3684_ (.A(_0920_),
    .B(_0938_),
    .C(_0948_),
    .X(_1354_));
 sky130_fd_sc_hd__and3_1 _3685_ (.A(_0852_),
    .B(_0941_),
    .C(_0950_),
    .X(_1355_));
 sky130_fd_sc_hd__a211o_1 _3686_ (.A1(_0674_),
    .A2(_1353_),
    .B1(_1354_),
    .C1(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__o22ai_4 _3687_ (.A1(_0879_),
    .A2(_1348_),
    .B1(_1352_),
    .B2(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__xor2_4 _3688_ (.A(\u0.E[1] ),
    .B(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__and3_1 _3689_ (.A(_0866_),
    .B(_0972_),
    .C(_0928_),
    .X(_1359_));
 sky130_fd_sc_hd__and3_1 _3690_ (.A(_0851_),
    .B(_0962_),
    .C(_0975_),
    .X(_1360_));
 sky130_fd_sc_hd__o211a_1 _3691_ (.A1(net74),
    .A2(_0848_),
    .B1(_0893_),
    .C1(_0971_),
    .X(_1361_));
 sky130_fd_sc_hd__and3_1 _3692_ (.A(_0825_),
    .B(_0812_),
    .C(_0953_),
    .X(_1362_));
 sky130_fd_sc_hd__or4_2 _3693_ (.A(_1359_),
    .B(_1360_),
    .C(_1361_),
    .D(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__a21o_1 _3694_ (.A1(_0963_),
    .A2(_1248_),
    .B1(_0901_),
    .X(_1364_));
 sky130_fd_sc_hd__and3_1 _3695_ (.A(_0913_),
    .B(_0965_),
    .C(_0961_),
    .X(_1365_));
 sky130_fd_sc_hd__and3_1 _3696_ (.A(_0818_),
    .B(_0966_),
    .C(_1284_),
    .X(_1366_));
 sky130_fd_sc_hd__a211o_1 _3697_ (.A1(_0674_),
    .A2(_1364_),
    .B1(_1365_),
    .C1(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__a21o_1 _3698_ (.A1(_0827_),
    .A2(_0942_),
    .B1(_0955_),
    .X(_1368_));
 sky130_fd_sc_hd__o21ai_4 _3699_ (.A1(_1363_),
    .A2(_1367_),
    .B1(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__mux2_1 _3700_ (.A0(net37),
    .A1(net716),
    .S(_0798_),
    .X(_1370_));
 sky130_fd_sc_hd__buf_2 _3701_ (.A(_1370_),
    .X(\u0.E[45] ));
 sky130_fd_sc_hd__xnor2_4 _3702_ (.A(_1369_),
    .B(\u0.E[45] ),
    .Y(_1371_));
 sky130_fd_sc_hd__buf_2 _3703_ (.A(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__o211a_1 _3704_ (.A1(net74),
    .A2(_0849_),
    .B1(_0974_),
    .C1(_1220_),
    .X(_1373_));
 sky130_fd_sc_hd__and3_1 _3705_ (.A(_0826_),
    .B(_0816_),
    .C(_0970_),
    .X(_1374_));
 sky130_fd_sc_hd__a311o_1 _3706_ (.A1(_0992_),
    .A2(_0926_),
    .A3(_0989_),
    .B1(_1373_),
    .C1(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__and3_1 _3707_ (.A(_0918_),
    .B(_0962_),
    .C(_0954_),
    .X(_1376_));
 sky130_fd_sc_hd__and3_1 _3708_ (.A(_0861_),
    .B(_1243_),
    .C(_1193_),
    .X(_1377_));
 sky130_fd_sc_hd__o211a_1 _3709_ (.A1(net112),
    .A2(_0858_),
    .B1(_0852_),
    .C1(_0966_),
    .X(_1378_));
 sky130_fd_sc_hd__o211a_1 _3710_ (.A1(net67),
    .A2(_0849_),
    .B1(_0894_),
    .C1(_0972_),
    .X(_1379_));
 sky130_fd_sc_hd__or4_2 _3711_ (.A(_1376_),
    .B(_1377_),
    .C(_1378_),
    .D(_1379_),
    .X(_1380_));
 sky130_fd_sc_hd__and3_1 _3712_ (.A(_0828_),
    .B(_0807_),
    .C(_0887_),
    .X(_1381_));
 sky130_fd_sc_hd__nor3_4 _3713_ (.A(_1375_),
    .B(_1380_),
    .C(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__mux2_1 _3714_ (.A0(net63),
    .A1(\R[1] ),
    .S(_0906_),
    .X(_1383_));
 sky130_fd_sc_hd__buf_4 _3715_ (.A(_1383_),
    .X(\u0.E[2] ));
 sky130_fd_sc_hd__xnor2_4 _3716_ (.A(_1382_),
    .B(\u0.E[2] ),
    .Y(_1384_));
 sky130_fd_sc_hd__mux2_1 _3717_ (.A0(_1358_),
    .A1(_1372_),
    .S(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__buf_2 _3718_ (.A(_1358_),
    .X(_1386_));
 sky130_fd_sc_hd__nand2_1 _3719_ (.A(_1386_),
    .B(_1372_),
    .Y(_1387_));
 sky130_fd_sc_hd__o21ai_1 _3720_ (.A1(_1346_),
    .A2(_1385_),
    .B1(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__o21ba_1 _3721_ (.A1(_1346_),
    .A2(_1386_),
    .B1_N(_1332_),
    .X(_1389_));
 sky130_fd_sc_hd__a22o_1 _3722_ (.A1(_1333_),
    .A2(_1388_),
    .B1(_1389_),
    .B2(_1387_),
    .X(_1390_));
 sky130_fd_sc_hd__inv_2 _3723_ (.A(_1384_),
    .Y(_1391_));
 sky130_fd_sc_hd__o21ai_2 _3724_ (.A1(_1358_),
    .A2(_1371_),
    .B1(_1332_),
    .Y(_1392_));
 sky130_fd_sc_hd__xnor2_1 _3725_ (.A(_1346_),
    .B(_1371_),
    .Y(_1393_));
 sky130_fd_sc_hd__nand2_1 _3726_ (.A(_1392_),
    .B(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__or2_1 _3727_ (.A(_1392_),
    .B(_1393_),
    .X(_1395_));
 sky130_fd_sc_hd__or2_1 _3728_ (.A(_1346_),
    .B(_1358_),
    .X(_1396_));
 sky130_fd_sc_hd__nor2_1 _3729_ (.A(_1386_),
    .B(_1372_),
    .Y(_1397_));
 sky130_fd_sc_hd__xor2_4 _3730_ (.A(_1344_),
    .B(\u0.E[46] ),
    .X(_1398_));
 sky130_fd_sc_hd__a221o_1 _3731_ (.A1(_1396_),
    .A2(_1372_),
    .B1(_1397_),
    .B2(_1398_),
    .C1(_1333_),
    .X(_1399_));
 sky130_fd_sc_hd__o21a_1 _3732_ (.A1(_1398_),
    .A2(_1372_),
    .B1(_1333_),
    .X(_1400_));
 sky130_fd_sc_hd__a21oi_1 _3733_ (.A1(_1396_),
    .A2(_1400_),
    .B1(_1391_),
    .Y(_1401_));
 sky130_fd_sc_hd__a32o_1 _3734_ (.A1(_1391_),
    .A2(_1394_),
    .A3(_1395_),
    .B1(_1399_),
    .B2(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__and3_1 _3735_ (.A(_0992_),
    .B(_0812_),
    .C(_1284_),
    .X(_1403_));
 sky130_fd_sc_hd__a31o_1 _3736_ (.A1(_0819_),
    .A2(_0961_),
    .A3(_0881_),
    .B1(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__and3_1 _3737_ (.A(_0843_),
    .B(_0963_),
    .C(_1214_),
    .X(_1405_));
 sky130_fd_sc_hd__and3_1 _3738_ (.A(_0947_),
    .B(_1248_),
    .C(_1289_),
    .X(_1406_));
 sky130_fd_sc_hd__a31o_1 _3739_ (.A1(_0868_),
    .A2(_0953_),
    .A3(_1221_),
    .B1(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__a311o_1 _3740_ (.A1(_0862_),
    .A2(_0971_),
    .A3(_0975_),
    .B1(_1405_),
    .C1(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__a311o_1 _3741_ (.A1(_0990_),
    .A2(_0965_),
    .A3(_0928_),
    .B1(_1404_),
    .C1(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__a31o_2 _3742_ (.A1(_0837_),
    .A2(_0808_),
    .A3(_0950_),
    .B1(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__xor2_4 _3743_ (.A(\u0.E[41] ),
    .B(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__mux2_2 _3744_ (.A0(_1390_),
    .A1(_1402_),
    .S(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__clkbuf_8 _3745_ (.A(_0905_),
    .X(_1413_));
 sky130_fd_sc_hd__mux2_1 _3746_ (.A0(net49),
    .A1(\L[15] ),
    .S(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__xnor2_2 _3747_ (.A(_1412_),
    .B(_1414_),
    .Y(\FP[15] ));
 sky130_fd_sc_hd__mux2_1 _3748_ (.A0(net346),
    .A1(\FP[15] ),
    .S(_1303_),
    .X(_1415_));
 sky130_fd_sc_hd__a22o_1 _3749_ (.A1(net708),
    .A2(_1319_),
    .B1(_0679_),
    .B2(_1415_),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _3750_ (.A0(net48),
    .A1(\R[23] ),
    .S(_0797_),
    .X(_1416_));
 sky130_fd_sc_hd__clkbuf_2 _3751_ (.A(_1416_),
    .X(\u0.E[34] ));
 sky130_fd_sc_hd__mux2_1 _3752_ (.A0(\fifo.rd_data[51] ),
    .A1(\u0.E[34] ),
    .S(_1303_),
    .X(_1417_));
 sky130_fd_sc_hd__a22o_1 _3753_ (.A1(net170),
    .A2(_1319_),
    .B1(_0679_),
    .B2(_1417_),
    .X(_0600_));
 sky130_fd_sc_hd__or2_4 _3754_ (.A(net111),
    .B(_1035_),
    .X(_1418_));
 sky130_fd_sc_hd__or2_2 _3755_ (.A(net71),
    .B(_0927_),
    .X(_1419_));
 sky130_fd_sc_hd__and3_1 _3756_ (.A(_0825_),
    .B(_1111_),
    .C(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__and3_1 _3757_ (.A(_0890_),
    .B(_1034_),
    .C(_1135_),
    .X(_1421_));
 sky130_fd_sc_hd__a311o_1 _3758_ (.A1(_0899_),
    .A2(_1105_),
    .A3(_1418_),
    .B1(_1420_),
    .C1(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__or2_2 _3759_ (.A(net108),
    .B(_0896_),
    .X(_1423_));
 sky130_fd_sc_hd__mux2_1 _3760_ (.A0(net76),
    .A1(net86),
    .S(_0896_),
    .X(_1424_));
 sky130_fd_sc_hd__a32o_1 _3761_ (.A1(_0893_),
    .A2(_1108_),
    .A3(_1423_),
    .B1(_1424_),
    .B2(_0860_),
    .X(_1425_));
 sky130_fd_sc_hd__buf_2 _3762_ (.A(net107),
    .X(_1426_));
 sky130_fd_sc_hd__or2_2 _3763_ (.A(net83),
    .B(_0988_),
    .X(_1427_));
 sky130_fd_sc_hd__o211a_1 _3764_ (.A1(_1426_),
    .A2(_0815_),
    .B1(_0851_),
    .C1(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__a311o_1 _3765_ (.A1(_0974_),
    .A2(_1041_),
    .A3(_1060_),
    .B1(_1425_),
    .C1(_1428_),
    .X(_1429_));
 sky130_fd_sc_hd__nand3_1 _3766_ (.A(_0806_),
    .B(_1067_),
    .C(_1125_),
    .Y(_1430_));
 sky130_fd_sc_hd__or3b_4 _3767_ (.A(_1422_),
    .B(_1429_),
    .C_N(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_1 _3768_ (.A0(net8),
    .A1(\R[2] ),
    .S(_0798_),
    .X(_1432_));
 sky130_fd_sc_hd__buf_2 _3769_ (.A(_1432_),
    .X(\u0.E[3] ));
 sky130_fd_sc_hd__xor2_4 _3770_ (.A(_1431_),
    .B(\u0.E[3] ),
    .X(_1433_));
 sky130_fd_sc_hd__buf_2 _3771_ (.A(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_1 _3772_ (.A0(net83),
    .A1(net92),
    .S(_0814_),
    .X(_1435_));
 sky130_fd_sc_hd__a32o_1 _3773_ (.A1(_0831_),
    .A2(_1090_),
    .A3(_1064_),
    .B1(_1435_),
    .B2(_0893_),
    .X(_1436_));
 sky130_fd_sc_hd__or2_1 _3774_ (.A(net102),
    .B(_0925_),
    .X(_1437_));
 sky130_fd_sc_hd__mux2_1 _3775_ (.A0(net93),
    .A1(net117),
    .S(_0927_),
    .X(_1438_));
 sky130_fd_sc_hd__a32o_1 _3776_ (.A1(_0825_),
    .A2(_1072_),
    .A3(_1437_),
    .B1(_1438_),
    .B2(_0851_),
    .X(_1439_));
 sky130_fd_sc_hd__mux2_1 _3777_ (.A0(net68),
    .A1(net107),
    .S(_0814_),
    .X(_1440_));
 sky130_fd_sc_hd__a32o_1 _3778_ (.A1(_0866_),
    .A2(_1071_),
    .A3(_1125_),
    .B1(_1440_),
    .B2(_0890_),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_1 _3779_ (.A0(net111),
    .A1(net86),
    .S(_0811_),
    .X(_1442_));
 sky130_fd_sc_hd__o21a_1 _3780_ (.A1(_0877_),
    .A2(_1442_),
    .B1(_0876_),
    .X(_1443_));
 sky130_fd_sc_hd__or4_1 _3781_ (.A(_1436_),
    .B(_1439_),
    .C(_1441_),
    .D(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__or2_1 _3782_ (.A(net115),
    .B(_0888_),
    .X(_1445_));
 sky130_fd_sc_hd__a21o_1 _3783_ (.A1(_1041_),
    .A2(_1445_),
    .B1(_0955_),
    .X(_1446_));
 sky130_fd_sc_hd__or2b_1 _3784_ (.A(net728),
    .B_N(_0798_),
    .X(_1447_));
 sky130_fd_sc_hd__o21ai_4 _3785_ (.A1(net17),
    .A2(_0906_),
    .B1(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__a21o_1 _3786_ (.A1(_1444_),
    .A2(_1446_),
    .B1(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__nand3_2 _3787_ (.A(_1444_),
    .B(_1446_),
    .C(_1448_),
    .Y(_1450_));
 sky130_fd_sc_hd__nand2_1 _3788_ (.A(_1449_),
    .B(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__nand2_1 _3789_ (.A(_1434_),
    .B(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hd__mux2_1 _3790_ (.A0(net109),
    .A1(net115),
    .S(_1035_),
    .X(_1453_));
 sky130_fd_sc_hd__a32o_1 _3791_ (.A1(_0841_),
    .A2(_1037_),
    .A3(_1060_),
    .B1(_1453_),
    .B2(_0831_),
    .X(_1454_));
 sky130_fd_sc_hd__mux2_1 _3792_ (.A0(net77),
    .A1(net84),
    .S(_0925_),
    .X(_1455_));
 sky130_fd_sc_hd__a32o_1 _3793_ (.A1(_0851_),
    .A2(_1049_),
    .A3(_1135_),
    .B1(_1455_),
    .B2(_1074_),
    .X(_1456_));
 sky130_fd_sc_hd__mux2_1 _3794_ (.A0(net108),
    .A1(net116),
    .S(_0925_),
    .X(_1457_));
 sky130_fd_sc_hd__a32o_1 _3795_ (.A1(_0890_),
    .A2(_1053_),
    .A3(_1427_),
    .B1(_1457_),
    .B2(_1089_),
    .X(_1458_));
 sky130_fd_sc_hd__mux2_1 _3796_ (.A0(_0702_),
    .A1(net99),
    .S(_1035_),
    .X(_1459_));
 sky130_fd_sc_hd__o21a_1 _3797_ (.A1(_0877_),
    .A2(_1459_),
    .B1(_0876_),
    .X(_1460_));
 sky130_fd_sc_hd__or4_4 _3798_ (.A(_1454_),
    .B(_1456_),
    .C(_1458_),
    .D(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__a21o_1 _3799_ (.A1(_1064_),
    .A2(_1130_),
    .B1(_0955_),
    .X(_1462_));
 sky130_fd_sc_hd__or2b_1 _3800_ (.A(\R[4] ),
    .B_N(_0930_),
    .X(_1463_));
 sky130_fd_sc_hd__o21ai_4 _3801_ (.A1(net26),
    .A2(_0905_),
    .B1(_1463_),
    .Y(_1464_));
 sky130_fd_sc_hd__a21o_2 _3802_ (.A1(_1461_),
    .A2(_1462_),
    .B1(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__nand3_4 _3803_ (.A(_1461_),
    .B(_1462_),
    .C(_1464_),
    .Y(_1466_));
 sky130_fd_sc_hd__a22o_1 _3804_ (.A1(_1449_),
    .A2(_1450_),
    .B1(_1465_),
    .B2(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__nand4_4 _3805_ (.A(_1449_),
    .B(_1450_),
    .C(_1465_),
    .D(_1466_),
    .Y(_1468_));
 sky130_fd_sc_hd__a21o_1 _3806_ (.A1(_1467_),
    .A2(_1468_),
    .B1(_1433_),
    .X(_1469_));
 sky130_fd_sc_hd__and3_1 _3807_ (.A(_0974_),
    .B(_1053_),
    .C(_1082_),
    .X(_1470_));
 sky130_fd_sc_hd__o211a_1 _3808_ (.A1(_1426_),
    .A2(_0858_),
    .B1(_1051_),
    .C1(_0832_),
    .X(_1471_));
 sky130_fd_sc_hd__a311o_1 _3809_ (.A1(_0990_),
    .A2(_1045_),
    .A3(_1108_),
    .B1(_1470_),
    .C1(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__mux2_1 _3810_ (.A0(net76),
    .A1(net116),
    .S(_0815_),
    .X(_1473_));
 sky130_fd_sc_hd__a32o_1 _3811_ (.A1(_0861_),
    .A2(_1041_),
    .A3(_1034_),
    .B1(_1473_),
    .B2(_0891_),
    .X(_1474_));
 sky130_fd_sc_hd__o211a_1 _3812_ (.A1(net119),
    .A2(_0858_),
    .B1(_0947_),
    .C1(_1105_),
    .X(_1475_));
 sky130_fd_sc_hd__a311o_1 _3813_ (.A1(_0843_),
    .A2(_1039_),
    .A3(_1111_),
    .B1(_1474_),
    .C1(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__or2_1 _3814_ (.A(net111),
    .B(_0927_),
    .X(_1477_));
 sky130_fd_sc_hd__and3_1 _3815_ (.A(_0807_),
    .B(_1477_),
    .C(_1091_),
    .X(_1478_));
 sky130_fd_sc_hd__nor3_4 _3816_ (.A(_1472_),
    .B(_1476_),
    .C(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__xnor2_4 _3817_ (.A(\u0.E[2] ),
    .B(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__a21o_1 _3818_ (.A1(_1452_),
    .A2(_1469_),
    .B1(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__xor2_2 _3819_ (.A(\u0.E[2] ),
    .B(_1479_),
    .X(_1482_));
 sky130_fd_sc_hd__buf_2 _3820_ (.A(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__and4_1 _3821_ (.A(_1433_),
    .B(_1451_),
    .C(_1465_),
    .D(_1466_),
    .X(_1484_));
 sky130_fd_sc_hd__and2_1 _3822_ (.A(_1449_),
    .B(_1450_),
    .X(_1485_));
 sky130_fd_sc_hd__buf_2 _3823_ (.A(_1485_),
    .X(_1486_));
 sky130_fd_sc_hd__nand2_4 _3824_ (.A(_1465_),
    .B(_1466_),
    .Y(_1487_));
 sky130_fd_sc_hd__o21ba_1 _3825_ (.A1(_1486_),
    .A2(_1487_),
    .B1_N(_1433_),
    .X(_1488_));
 sky130_fd_sc_hd__and3_1 _3826_ (.A(_1096_),
    .B(_1042_),
    .C(_1418_),
    .X(_1489_));
 sky130_fd_sc_hd__or2_1 _3827_ (.A(net77),
    .B(_1035_),
    .X(_1490_));
 sky130_fd_sc_hd__and3_1 _3828_ (.A(_0913_),
    .B(_1490_),
    .C(_1427_),
    .X(_1491_));
 sky130_fd_sc_hd__a311o_1 _3829_ (.A1(_0891_),
    .A2(_1082_),
    .A3(_1052_),
    .B1(_1489_),
    .C1(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__clkbuf_4 _3830_ (.A(net76),
    .X(_1493_));
 sky130_fd_sc_hd__o211a_1 _3831_ (.A1(_1493_),
    .A2(_0858_),
    .B1(_0868_),
    .C1(_1046_),
    .X(_1494_));
 sky130_fd_sc_hd__and3_1 _3832_ (.A(_0861_),
    .B(_1060_),
    .C(_1135_),
    .X(_1495_));
 sky130_fd_sc_hd__and3_1 _3833_ (.A(_0920_),
    .B(_1423_),
    .C(_1445_),
    .X(_1496_));
 sky130_fd_sc_hd__a31o_1 _3834_ (.A1(_0842_),
    .A2(_1036_),
    .A3(_1419_),
    .B1(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__or4_1 _3835_ (.A(_1492_),
    .B(_1494_),
    .C(_1495_),
    .D(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__a31o_1 _3836_ (.A1(_0808_),
    .A2(_1437_),
    .A3(_1132_),
    .B1(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_1 _3837_ (.A0(net34),
    .A1(\R[5] ),
    .S(_0906_),
    .X(_1500_));
 sky130_fd_sc_hd__buf_2 _3838_ (.A(_1500_),
    .X(\u0.E[6] ));
 sky130_fd_sc_hd__xor2_2 _3839_ (.A(_1499_),
    .B(\u0.E[6] ),
    .X(_1501_));
 sky130_fd_sc_hd__o31a_1 _3840_ (.A1(_1483_),
    .A2(_1484_),
    .A3(_1488_),
    .B1(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__nand2_1 _3841_ (.A(_1434_),
    .B(_1467_),
    .Y(_1503_));
 sky130_fd_sc_hd__a31o_1 _3842_ (.A1(_1483_),
    .A2(_1468_),
    .A3(_1503_),
    .B1(_1501_),
    .X(_1504_));
 sky130_fd_sc_hd__xor2_1 _3843_ (.A(_1433_),
    .B(_1467_),
    .X(_1505_));
 sky130_fd_sc_hd__nor2_1 _3844_ (.A(_1483_),
    .B(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__o2bb2a_1 _3845_ (.A1_N(_1481_),
    .A2_N(_1502_),
    .B1(_1504_),
    .B2(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__or2_1 _3846_ (.A(_1485_),
    .B(_1487_),
    .X(_1508_));
 sky130_fd_sc_hd__nand2_2 _3847_ (.A(_1433_),
    .B(_1487_),
    .Y(_1509_));
 sky130_fd_sc_hd__a21oi_1 _3848_ (.A1(_1434_),
    .A2(_1486_),
    .B1(_1482_),
    .Y(_1510_));
 sky130_fd_sc_hd__a32o_1 _3849_ (.A1(_1483_),
    .A2(_1508_),
    .A3(_1509_),
    .B1(_1510_),
    .B2(_1469_),
    .X(_1511_));
 sky130_fd_sc_hd__or2_1 _3850_ (.A(_1433_),
    .B(_1468_),
    .X(_1512_));
 sky130_fd_sc_hd__a21oi_1 _3851_ (.A1(_1434_),
    .A2(_1486_),
    .B1(_1480_),
    .Y(_1513_));
 sky130_fd_sc_hd__nand2_1 _3852_ (.A(_1467_),
    .B(_1468_),
    .Y(_1514_));
 sky130_fd_sc_hd__a32oi_1 _3853_ (.A1(_1480_),
    .A2(_1509_),
    .A3(_1512_),
    .B1(_1513_),
    .B2(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__clkbuf_4 _3854_ (.A(_1501_),
    .X(_1516_));
 sky130_fd_sc_hd__mux2_1 _3855_ (.A0(_1511_),
    .A1(_1515_),
    .S(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__buf_4 _3856_ (.A(net68),
    .X(_1518_));
 sky130_fd_sc_hd__o211a_1 _3857_ (.A1(_1518_),
    .A2(_0859_),
    .B1(_0853_),
    .C1(_1128_),
    .X(_1519_));
 sky130_fd_sc_hd__and3_1 _3858_ (.A(_0832_),
    .B(_1114_),
    .C(_1122_),
    .X(_1520_));
 sky130_fd_sc_hd__a311o_1 _3859_ (.A1(_0819_),
    .A2(_1068_),
    .A3(_1121_),
    .B1(_1519_),
    .C1(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__or2_1 _3860_ (.A(_0750_),
    .B(_0858_),
    .X(_1522_));
 sky130_fd_sc_hd__and3_1 _3861_ (.A(_0868_),
    .B(_1522_),
    .C(_1130_),
    .X(_1523_));
 sky130_fd_sc_hd__and3_1 _3862_ (.A(_0862_),
    .B(_1120_),
    .C(_1129_),
    .X(_1524_));
 sky130_fd_sc_hd__and3_1 _3863_ (.A(_0990_),
    .B(_1132_),
    .C(_1033_),
    .X(_1525_));
 sky130_fd_sc_hd__a31o_1 _3864_ (.A1(_0843_),
    .A2(_1091_),
    .A3(_1125_),
    .B1(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__or4_2 _3865_ (.A(_1521_),
    .B(_1523_),
    .C(_1524_),
    .D(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__a31oi_4 _3866_ (.A1(_0808_),
    .A2(_1039_),
    .A3(_1423_),
    .B1(_1527_),
    .Y(_1528_));
 sky130_fd_sc_hd__xnor2_2 _3867_ (.A(\u0.E[1] ),
    .B(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__mux2_1 _3868_ (.A0(_1507_),
    .A1(_1517_),
    .S(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _3869_ (.A0(net47),
    .A1(net703),
    .S(_1413_),
    .X(_1531_));
 sky130_fd_sc_hd__xnor2_1 _3870_ (.A(_1530_),
    .B(_1531_),
    .Y(\FP[23] ));
 sky130_fd_sc_hd__mux2_1 _3871_ (.A0(\fifo.rd_data[50] ),
    .A1(\FP[23] ),
    .S(_1303_),
    .X(_1532_));
 sky130_fd_sc_hd__a22o_1 _3872_ (.A1(net169),
    .A2(_1319_),
    .B1(_0679_),
    .B2(_1532_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _3873_ (.A0(\fifo.rd_data[49] ),
    .A1(\u0.E[46] ),
    .S(_1303_),
    .X(_1533_));
 sky130_fd_sc_hd__a22o_1 _3874_ (.A1(net719),
    .A2(_1319_),
    .B1(_0679_),
    .B2(_1533_),
    .X(_0598_));
 sky130_fd_sc_hd__inv_2 _3875_ (.A(_1529_),
    .Y(_1534_));
 sky130_fd_sc_hd__and3_2 _3876_ (.A(_1433_),
    .B(_1467_),
    .C(_1468_),
    .X(_1535_));
 sky130_fd_sc_hd__nor2_1 _3877_ (.A(_1434_),
    .B(_1486_),
    .Y(_1536_));
 sky130_fd_sc_hd__nor2_1 _3878_ (.A(_1433_),
    .B(_1487_),
    .Y(_1537_));
 sky130_fd_sc_hd__a21oi_2 _3879_ (.A1(_1486_),
    .A2(_1487_),
    .B1(_1482_),
    .Y(_1538_));
 sky130_fd_sc_hd__a21oi_1 _3880_ (.A1(_1509_),
    .A2(_1538_),
    .B1(_1516_),
    .Y(_1539_));
 sky130_fd_sc_hd__o41a_1 _3881_ (.A1(_1480_),
    .A2(_1535_),
    .A3(_1536_),
    .A4(_1537_),
    .B1(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__nand2_1 _3882_ (.A(_1434_),
    .B(_1468_),
    .Y(_1541_));
 sky130_fd_sc_hd__and3_1 _3883_ (.A(_1483_),
    .B(_1512_),
    .C(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__o21a_1 _3884_ (.A1(_1506_),
    .A2(_1542_),
    .B1(_1516_),
    .X(_1543_));
 sky130_fd_sc_hd__or3_1 _3885_ (.A(_1538_),
    .B(_1535_),
    .C(_1536_),
    .X(_1544_));
 sky130_fd_sc_hd__o21ai_1 _3886_ (.A1(_1535_),
    .A2(_1536_),
    .B1(_1538_),
    .Y(_1545_));
 sky130_fd_sc_hd__a21oi_1 _3887_ (.A1(_1544_),
    .A2(_1545_),
    .B1(_1516_),
    .Y(_1546_));
 sky130_fd_sc_hd__o2bb2a_1 _3888_ (.A1_N(_1469_),
    .A2_N(_1513_),
    .B1(_1505_),
    .B2(_1483_),
    .X(_1547_));
 sky130_fd_sc_hd__a21o_1 _3889_ (.A1(_1516_),
    .A2(_1547_),
    .B1(_1529_),
    .X(_1548_));
 sky130_fd_sc_hd__o32a_2 _3890_ (.A1(_1534_),
    .A2(_1540_),
    .A3(_1543_),
    .B1(_1546_),
    .B2(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__mux2_2 _3891_ (.A0(net44),
    .A1(\L[31] ),
    .S(_1413_),
    .X(_1550_));
 sky130_fd_sc_hd__xnor2_4 _3892_ (.A(_1549_),
    .B(_1550_),
    .Y(\FP[31] ));
 sky130_fd_sc_hd__mux2_1 _3893_ (.A0(net465),
    .A1(\FP[31] ),
    .S(_1303_),
    .X(_1551_));
 sky130_fd_sc_hd__a22o_1 _3894_ (.A1(net166),
    .A2(_1319_),
    .B1(_0679_),
    .B2(_1551_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _3895_ (.A0(net43),
    .A1(\R[6] ),
    .S(_0930_),
    .X(_1552_));
 sky130_fd_sc_hd__buf_4 _3896_ (.A(_1552_),
    .X(\u0.E[9] ));
 sky130_fd_sc_hd__mux2_1 _3897_ (.A0(net418),
    .A1(\u0.E[9] ),
    .S(_1303_),
    .X(_1553_));
 sky130_fd_sc_hd__a22o_1 _3898_ (.A1(net689),
    .A2(_1319_),
    .B1(_0679_),
    .B2(_1553_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _3899_ (.A0(_1151_),
    .A1(_1139_),
    .S(_1081_),
    .X(_1554_));
 sky130_fd_sc_hd__xnor2_1 _3900_ (.A(_1174_),
    .B(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__xnor2_1 _3901_ (.A(_1141_),
    .B(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__nor2_1 _3902_ (.A(_1157_),
    .B(_1178_),
    .Y(_1557_));
 sky130_fd_sc_hd__o21a_1 _3903_ (.A1(_1152_),
    .A2(_1157_),
    .B1(_1141_),
    .X(_1558_));
 sky130_fd_sc_hd__a211oi_1 _3904_ (.A1(_1118_),
    .A2(_1557_),
    .B1(_1558_),
    .C1(_1174_),
    .Y(_1559_));
 sky130_fd_sc_hd__nand2_1 _3905_ (.A(_1118_),
    .B(_1150_),
    .Y(_1560_));
 sky130_fd_sc_hd__o31a_1 _3906_ (.A1(_1118_),
    .A2(_1140_),
    .A3(_1179_),
    .B1(_1174_),
    .X(_1561_));
 sky130_fd_sc_hd__a21o_1 _3907_ (.A1(_1560_),
    .A2(_1561_),
    .B1(_1059_),
    .X(_1562_));
 sky130_fd_sc_hd__o2bb2a_1 _3908_ (.A1_N(_1059_),
    .A2_N(_1556_),
    .B1(_1559_),
    .B2(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__mux2_1 _3909_ (.A0(net42),
    .A1(net509),
    .S(_1413_),
    .X(_1564_));
 sky130_fd_sc_hd__xnor2_1 _3910_ (.A(_1563_),
    .B(_1564_),
    .Y(\FP[6] ));
 sky130_fd_sc_hd__buf_4 _3911_ (.A(_1302_),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_1 _3912_ (.A0(net231),
    .A1(\FP[6] ),
    .S(_1565_),
    .X(_1566_));
 sky130_fd_sc_hd__a22o_1 _3913_ (.A1(net164),
    .A2(_1319_),
    .B1(_0679_),
    .B2(_1566_),
    .X(_0595_));
 sky130_fd_sc_hd__clkbuf_4 _3914_ (.A(_1305_),
    .X(_1567_));
 sky130_fd_sc_hd__mux2_1 _3915_ (.A0(net41),
    .A1(\R[14] ),
    .S(_0798_),
    .X(_1568_));
 sky130_fd_sc_hd__buf_2 _3916_ (.A(_1568_),
    .X(\u0.E[21] ));
 sky130_fd_sc_hd__mux2_1 _3917_ (.A0(net422),
    .A1(\u0.E[21] ),
    .S(_1565_),
    .X(_1569_));
 sky130_fd_sc_hd__a22o_1 _3918_ (.A1(net163),
    .A2(_1319_),
    .B1(_1567_),
    .B2(_1569_),
    .X(_0594_));
 sky130_fd_sc_hd__xor2_2 _3919_ (.A(_0873_),
    .B(\u0.E[23] ),
    .X(_1570_));
 sky130_fd_sc_hd__o21ba_1 _3920_ (.A1(_1009_),
    .A2(_0936_),
    .B1_N(_0959_),
    .X(_1571_));
 sky130_fd_sc_hd__nor2_1 _3921_ (.A(_1025_),
    .B(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__o21ai_2 _3922_ (.A1(_0936_),
    .A2(_1010_),
    .B1(_0982_),
    .Y(_1573_));
 sky130_fd_sc_hd__o221a_1 _3923_ (.A1(_0983_),
    .A2(_1572_),
    .B1(_1573_),
    .B2(_1018_),
    .C1(_1005_),
    .X(_1574_));
 sky130_fd_sc_hd__a21o_1 _3924_ (.A1(_1007_),
    .A2(_1008_),
    .B1(_0959_),
    .X(_1575_));
 sky130_fd_sc_hd__or2b_1 _3925_ (.A(_1025_),
    .B_N(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__nand2_1 _3926_ (.A(_0936_),
    .B(_1010_),
    .Y(_1577_));
 sky130_fd_sc_hd__a31o_1 _3927_ (.A1(_0985_),
    .A2(_1577_),
    .A3(_1575_),
    .B1(_1005_),
    .X(_1578_));
 sky130_fd_sc_hd__a21oi_1 _3928_ (.A1(_0983_),
    .A2(_1576_),
    .B1(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__inv_2 _3929_ (.A(_1013_),
    .Y(_1580_));
 sky130_fd_sc_hd__o21a_1 _3930_ (.A1(_1010_),
    .A2(_1018_),
    .B1(_1013_),
    .X(_1581_));
 sky130_fd_sc_hd__o221a_1 _3931_ (.A1(_1580_),
    .A2(_1573_),
    .B1(_1581_),
    .B2(_0983_),
    .C1(_1019_),
    .X(_1582_));
 sky130_fd_sc_hd__a21oi_1 _3932_ (.A1(_0985_),
    .A2(_1009_),
    .B1(_0960_),
    .Y(_1583_));
 sky130_fd_sc_hd__a31o_1 _3933_ (.A1(_0985_),
    .A2(_1009_),
    .A3(_0960_),
    .B1(_1019_),
    .X(_1584_));
 sky130_fd_sc_hd__o21ai_1 _3934_ (.A1(_1583_),
    .A2(_1584_),
    .B1(_1570_),
    .Y(_1585_));
 sky130_fd_sc_hd__o32a_2 _3935_ (.A1(_1570_),
    .A2(_1574_),
    .A3(_1579_),
    .B1(_1582_),
    .B2(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__mux2_1 _3936_ (.A0(net40),
    .A1(net673),
    .S(_1030_),
    .X(_1587_));
 sky130_fd_sc_hd__xor2_1 _3937_ (.A(_1586_),
    .B(_1587_),
    .X(\FP[14] ));
 sky130_fd_sc_hd__mux2_1 _3938_ (.A0(net232),
    .A1(\FP[14] ),
    .S(_1565_),
    .X(_1588_));
 sky130_fd_sc_hd__a22o_1 _3939_ (.A1(net162),
    .A2(_1319_),
    .B1(_1567_),
    .B2(_1588_),
    .X(_0593_));
 sky130_fd_sc_hd__buf_4 _3940_ (.A(_0670_),
    .X(_1589_));
 sky130_fd_sc_hd__mux2_1 _3941_ (.A0(net39),
    .A1(\R[22] ),
    .S(_0797_),
    .X(_1590_));
 sky130_fd_sc_hd__clkbuf_8 _3942_ (.A(_1590_),
    .X(\u0.E[33] ));
 sky130_fd_sc_hd__mux2_1 _3943_ (.A0(net436),
    .A1(\u0.E[33] ),
    .S(_1565_),
    .X(_1591_));
 sky130_fd_sc_hd__a22o_1 _3944_ (.A1(net161),
    .A2(_1589_),
    .B1(_1567_),
    .B2(_1591_),
    .X(_0592_));
 sky130_fd_sc_hd__or2_1 _3945_ (.A(_1235_),
    .B(_1266_),
    .X(_1592_));
 sky130_fd_sc_hd__a21bo_1 _3946_ (.A1(_1235_),
    .A2(_1261_),
    .B1_N(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__nor2_1 _3947_ (.A(_1219_),
    .B(_1261_),
    .Y(_1594_));
 sky130_fd_sc_hd__a21oi_1 _3948_ (.A1(_1219_),
    .A2(_1593_),
    .B1(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__a211oi_1 _3949_ (.A1(_1235_),
    .A2(_1247_),
    .B1(_1277_),
    .C1(_1219_),
    .Y(_1596_));
 sky130_fd_sc_hd__a211o_1 _3950_ (.A1(_1219_),
    .A2(_1593_),
    .B1(_1596_),
    .C1(_1204_),
    .X(_1597_));
 sky130_fd_sc_hd__o211a_1 _3951_ (.A1(_1205_),
    .A2(_1595_),
    .B1(_1597_),
    .C1(_1294_),
    .X(_1598_));
 sky130_fd_sc_hd__nor3_1 _3952_ (.A(_1235_),
    .B(_1267_),
    .C(_1218_),
    .Y(_1599_));
 sky130_fd_sc_hd__a21oi_1 _3953_ (.A1(_1219_),
    .A2(_1275_),
    .B1(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__xnor2_1 _3954_ (.A(_1266_),
    .B(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__a21o_1 _3955_ (.A1(_1592_),
    .A2(_1308_),
    .B1(_1260_),
    .X(_1602_));
 sky130_fd_sc_hd__o211a_1 _3956_ (.A1(_1267_),
    .A2(_1219_),
    .B1(_1204_),
    .C1(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__a211oi_1 _3957_ (.A1(_1205_),
    .A2(_1601_),
    .B1(_1603_),
    .C1(_1294_),
    .Y(_1604_));
 sky130_fd_sc_hd__mux2_1 _3958_ (.A0(net38),
    .A1(net710),
    .S(_1030_),
    .X(_1605_));
 sky130_fd_sc_hd__or3_1 _3959_ (.A(_1598_),
    .B(_1604_),
    .C(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__o21ai_1 _3960_ (.A1(_1598_),
    .A2(_1604_),
    .B1(_1605_),
    .Y(_1607_));
 sky130_fd_sc_hd__nand3_1 _3961_ (.A(_0766_),
    .B(_1606_),
    .C(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__or2_1 _3962_ (.A(\fifo.rd_data[42] ),
    .B(_1303_),
    .X(_1609_));
 sky130_fd_sc_hd__a32o_1 _3963_ (.A1(_1305_),
    .A2(_1608_),
    .A3(_1609_),
    .B1(_0670_),
    .B2(net160),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _3964_ (.A0(net701),
    .A1(\u0.E[45] ),
    .S(_1565_),
    .X(_1610_));
 sky130_fd_sc_hd__a22o_1 _3965_ (.A1(net159),
    .A2(_1589_),
    .B1(_1567_),
    .B2(_1610_),
    .X(_0590_));
 sky130_fd_sc_hd__nand2_1 _3966_ (.A(_1141_),
    .B(_1150_),
    .Y(_1611_));
 sky130_fd_sc_hd__or3b_1 _3967_ (.A(_1141_),
    .B(_1151_),
    .C_N(_1081_),
    .X(_1612_));
 sky130_fd_sc_hd__and3b_1 _3968_ (.A_N(_1174_),
    .B(_1182_),
    .C(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__nand2_1 _3969_ (.A(_1141_),
    .B(_1151_),
    .Y(_1614_));
 sky130_fd_sc_hd__nand2_1 _3970_ (.A(_1157_),
    .B(_1614_),
    .Y(_1615_));
 sky130_fd_sc_hd__nand2_1 _3971_ (.A(_1081_),
    .B(_1142_),
    .Y(_1616_));
 sky130_fd_sc_hd__o221a_1 _3972_ (.A1(_1151_),
    .A2(_1616_),
    .B1(_1157_),
    .B2(_1614_),
    .C1(_1174_),
    .X(_1617_));
 sky130_fd_sc_hd__a22o_1 _3973_ (.A1(_1611_),
    .A2(_1613_),
    .B1(_1615_),
    .B2(_1617_),
    .X(_1618_));
 sky130_fd_sc_hd__o2bb2a_1 _3974_ (.A1_N(_1154_),
    .A2_N(_1150_),
    .B1(_1616_),
    .B2(_1151_),
    .X(_1619_));
 sky130_fd_sc_hd__and3_1 _3975_ (.A(_1081_),
    .B(_1103_),
    .C(_1139_),
    .X(_1620_));
 sky130_fd_sc_hd__o31a_1 _3976_ (.A1(_1140_),
    .A2(_1158_),
    .A3(_1620_),
    .B1(_1174_),
    .X(_1621_));
 sky130_fd_sc_hd__a2bb2o_1 _3977_ (.A1_N(_1174_),
    .A2_N(_1619_),
    .B1(_1621_),
    .B2(_1180_),
    .X(_1622_));
 sky130_fd_sc_hd__mux2_1 _3978_ (.A0(_1618_),
    .A1(_1622_),
    .S(_1059_),
    .X(_1623_));
 sky130_fd_sc_hd__buf_4 _3979_ (.A(_0905_),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(net36),
    .A1(net518),
    .S(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__xnor2_1 _3981_ (.A(_1623_),
    .B(_1625_),
    .Y(\FP[30] ));
 sky130_fd_sc_hd__mux2_1 _3982_ (.A0(\fifo.rd_data[40] ),
    .A1(\FP[30] ),
    .S(_1565_),
    .X(_1626_));
 sky130_fd_sc_hd__a22o_1 _3983_ (.A1(net158),
    .A2(_1589_),
    .B1(_1567_),
    .B2(_1626_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _3984_ (.A0(net731),
    .A1(\u0.E[6] ),
    .S(_1565_),
    .X(_1627_));
 sky130_fd_sc_hd__a22o_1 _3985_ (.A1(net156),
    .A2(_1589_),
    .B1(_1567_),
    .B2(_1627_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _3986_ (.A0(net33),
    .A1(net702),
    .S(_1413_),
    .X(_1628_));
 sky130_fd_sc_hd__nand3_1 _3987_ (.A(_1398_),
    .B(_1386_),
    .C(_1372_),
    .Y(_1629_));
 sky130_fd_sc_hd__a21o_1 _3988_ (.A1(_1398_),
    .A2(_1358_),
    .B1(_1372_),
    .X(_1630_));
 sky130_fd_sc_hd__o21ai_1 _3989_ (.A1(_1398_),
    .A2(_1386_),
    .B1(_1333_),
    .Y(_1631_));
 sky130_fd_sc_hd__a21o_1 _3990_ (.A1(_1629_),
    .A2(_1630_),
    .B1(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__nand3_1 _3991_ (.A(_1629_),
    .B(_1631_),
    .C(_1630_),
    .Y(_1633_));
 sky130_fd_sc_hd__a211o_1 _3992_ (.A1(_1398_),
    .A2(_1371_),
    .B1(_1332_),
    .C1(_1358_),
    .X(_1634_));
 sky130_fd_sc_hd__o211a_1 _3993_ (.A1(_1333_),
    .A2(_1629_),
    .B1(_1634_),
    .C1(_1391_),
    .X(_1635_));
 sky130_fd_sc_hd__a21oi_1 _3994_ (.A1(_1346_),
    .A2(_1386_),
    .B1(_1372_),
    .Y(_1636_));
 sky130_fd_sc_hd__and3_1 _3995_ (.A(_1346_),
    .B(_1358_),
    .C(_1371_),
    .X(_1637_));
 sky130_fd_sc_hd__or3b_1 _3996_ (.A(_1636_),
    .B(_1637_),
    .C_N(_1333_),
    .X(_1638_));
 sky130_fd_sc_hd__a32o_1 _3997_ (.A1(_1384_),
    .A2(_1632_),
    .A3(_1633_),
    .B1(_1635_),
    .B2(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__a21oi_1 _3998_ (.A1(_1386_),
    .A2(_1372_),
    .B1(_1346_),
    .Y(_1640_));
 sky130_fd_sc_hd__o21a_1 _3999_ (.A1(_1637_),
    .A2(_1640_),
    .B1(_1333_),
    .X(_1641_));
 sky130_fd_sc_hd__a21o_1 _4000_ (.A1(_1387_),
    .A2(_1389_),
    .B1(_1384_),
    .X(_1642_));
 sky130_fd_sc_hd__o21ai_1 _4001_ (.A1(_1398_),
    .A2(_1386_),
    .B1(_1372_),
    .Y(_1643_));
 sky130_fd_sc_hd__or3_1 _4002_ (.A(_1398_),
    .B(_1358_),
    .C(_1371_),
    .X(_1644_));
 sky130_fd_sc_hd__o21ba_1 _4003_ (.A1(_1358_),
    .A2(_1371_),
    .B1_N(_1332_),
    .X(_1645_));
 sky130_fd_sc_hd__nand2_1 _4004_ (.A(_1398_),
    .B(_1386_),
    .Y(_1646_));
 sky130_fd_sc_hd__a32o_1 _4005_ (.A1(_1333_),
    .A2(_1643_),
    .A3(_1644_),
    .B1(_1645_),
    .B2(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__a2bb2o_1 _4006_ (.A1_N(_1641_),
    .A2_N(_1642_),
    .B1(_1647_),
    .B2(_1384_),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_1 _4007_ (.A0(_1639_),
    .A1(_1648_),
    .S(_1411_),
    .X(_1649_));
 sky130_fd_sc_hd__xor2_1 _4008_ (.A(_1628_),
    .B(_1649_),
    .X(\FP[5] ));
 sky130_fd_sc_hd__mux2_1 _4009_ (.A0(\fifo.rd_data[38] ),
    .A1(\FP[5] ),
    .S(_1565_),
    .X(_1650_));
 sky130_fd_sc_hd__a22o_1 _4010_ (.A1(net692),
    .A2(_1589_),
    .B1(_1567_),
    .B2(_1650_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _4011_ (.A0(\fifo.rd_data[37] ),
    .A1(\u0.E[18] ),
    .S(_1565_),
    .X(_1651_));
 sky130_fd_sc_hd__a22o_1 _4012_ (.A1(net695),
    .A2(_1589_),
    .B1(_1567_),
    .B2(_1651_),
    .X(_0586_));
 sky130_fd_sc_hd__and3_1 _4013_ (.A(_1074_),
    .B(_1105_),
    .C(_1041_),
    .X(_1652_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(net119),
    .A1(_0711_),
    .S(_0836_),
    .X(_1653_));
 sky130_fd_sc_hd__a32o_1 _4015_ (.A1(_0818_),
    .A2(_1039_),
    .A3(_1418_),
    .B1(_1653_),
    .B2(_0867_),
    .X(_1654_));
 sky130_fd_sc_hd__a311o_1 _4016_ (.A1(_0947_),
    .A2(_1045_),
    .A3(_1082_),
    .B1(_1652_),
    .C1(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__mux2_1 _4017_ (.A0(net107),
    .A1(net117),
    .S(_0836_),
    .X(_1656_));
 sky130_fd_sc_hd__o21a_1 _4018_ (.A1(_0901_),
    .A2(_1656_),
    .B1(_0876_),
    .X(_1657_));
 sky130_fd_sc_hd__o211a_1 _4019_ (.A1(_1493_),
    .A2(_0858_),
    .B1(_0894_),
    .C1(_1051_),
    .X(_1658_));
 sky130_fd_sc_hd__a311o_1 _4020_ (.A1(_0832_),
    .A2(_1034_),
    .A3(_1111_),
    .B1(_1657_),
    .C1(_1658_),
    .X(_1659_));
 sky130_fd_sc_hd__a21o_1 _4021_ (.A1(_1072_),
    .A2(_1121_),
    .B1(_0879_),
    .X(_1660_));
 sky130_fd_sc_hd__o21ai_4 _4022_ (.A1(_1655_),
    .A2(_1659_),
    .B1(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__xor2_4 _4023_ (.A(\u0.E[9] ),
    .B(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__a21o_1 _4024_ (.A1(_1105_),
    .A2(_1052_),
    .B1(_0879_),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _4025_ (.A0(net75),
    .A1(net101),
    .S(_0969_),
    .X(_1664_));
 sky130_fd_sc_hd__o21a_1 _4026_ (.A1(_0877_),
    .A2(_1664_),
    .B1(_0876_),
    .X(_1665_));
 sky130_fd_sc_hd__or2_1 _4027_ (.A(net92),
    .B(_0834_),
    .X(_1666_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(_0757_),
    .A1(net117),
    .S(_0969_),
    .X(_1667_));
 sky130_fd_sc_hd__a32o_1 _4029_ (.A1(_1089_),
    .A2(_1114_),
    .A3(_1666_),
    .B1(_1667_),
    .B2(_0818_),
    .X(_1668_));
 sky130_fd_sc_hd__mux2_1 _4030_ (.A0(_0705_),
    .A1(net116),
    .S(_0969_),
    .X(_1669_));
 sky130_fd_sc_hd__a32o_1 _4031_ (.A1(_1096_),
    .A2(_1032_),
    .A3(_1091_),
    .B1(_1669_),
    .B2(_1074_),
    .X(_1670_));
 sky130_fd_sc_hd__mux2_1 _4032_ (.A0(_0708_),
    .A1(net79),
    .S(_0940_),
    .X(_1671_));
 sky130_fd_sc_hd__a32o_1 _4033_ (.A1(_0831_),
    .A2(_1067_),
    .A3(_1130_),
    .B1(_1671_),
    .B2(_0841_),
    .X(_1672_));
 sky130_fd_sc_hd__or4_2 _4034_ (.A(_1665_),
    .B(_1668_),
    .C(_1670_),
    .D(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__a21boi_4 _4035_ (.A1(_1663_),
    .A2(_1673_),
    .B1_N(\u0.E[10] ),
    .Y(_1674_));
 sky130_fd_sc_hd__and3b_2 _4036_ (.A_N(\u0.E[10] ),
    .B(_1663_),
    .C(_1673_),
    .X(_1675_));
 sky130_fd_sc_hd__a21o_1 _4037_ (.A1(_1666_),
    .A2(_1129_),
    .B1(_0879_),
    .X(_1676_));
 sky130_fd_sc_hd__mux2_1 _4038_ (.A0(net119),
    .A1(_1038_),
    .S(_0836_),
    .X(_1677_));
 sky130_fd_sc_hd__o21a_1 _4039_ (.A1(_0901_),
    .A2(_1677_),
    .B1(_0674_),
    .X(_1678_));
 sky130_fd_sc_hd__mux2_1 _4040_ (.A0(net84),
    .A1(net107),
    .S(_0834_),
    .X(_1679_));
 sky130_fd_sc_hd__a32o_1 _4041_ (.A1(_1089_),
    .A2(_1108_),
    .A3(_1052_),
    .B1(_1679_),
    .B2(_0918_),
    .X(_1680_));
 sky130_fd_sc_hd__mux2_1 _4042_ (.A0(net79),
    .A1(net85),
    .S(_0940_),
    .X(_1681_));
 sky130_fd_sc_hd__a32o_1 _4043_ (.A1(_1096_),
    .A2(_1037_),
    .A3(_1034_),
    .B1(_1681_),
    .B2(_0920_),
    .X(_1682_));
 sky130_fd_sc_hd__mux2_1 _4044_ (.A0(_0718_),
    .A1(net116),
    .S(_0940_),
    .X(_1683_));
 sky130_fd_sc_hd__a32o_1 _4045_ (.A1(_0841_),
    .A2(_1041_),
    .A3(_1049_),
    .B1(_1683_),
    .B2(_0913_),
    .X(_1684_));
 sky130_fd_sc_hd__or4_4 _4046_ (.A(_1678_),
    .B(_1680_),
    .C(_1682_),
    .D(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__a21o_2 _4047_ (.A1(_1676_),
    .A2(_1685_),
    .B1(\u0.E[11] ),
    .X(_1686_));
 sky130_fd_sc_hd__nand3_4 _4048_ (.A(\u0.E[11] ),
    .B(_1676_),
    .C(_1685_),
    .Y(_1687_));
 sky130_fd_sc_hd__or4bb_1 _4049_ (.A(_1674_),
    .B(_1675_),
    .C_N(_1686_),
    .D_N(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__o21a_1 _4050_ (.A1(_1048_),
    .A2(_0859_),
    .B1(_1427_),
    .X(_1689_));
 sky130_fd_sc_hd__and3_1 _4051_ (.A(_1096_),
    .B(_1067_),
    .C(_1477_),
    .X(_1690_));
 sky130_fd_sc_hd__and3_1 _4052_ (.A(_1074_),
    .B(_1090_),
    .C(_1071_),
    .X(_1691_));
 sky130_fd_sc_hd__and3_1 _4053_ (.A(_1089_),
    .B(_1072_),
    .C(_1094_),
    .X(_1692_));
 sky130_fd_sc_hd__and3_1 _4054_ (.A(_0818_),
    .B(_1064_),
    .C(_1086_),
    .X(_1693_));
 sky130_fd_sc_hd__or4_1 _4055_ (.A(_1690_),
    .B(_1691_),
    .C(_1692_),
    .D(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__mux2_1 _4056_ (.A0(_0755_),
    .A1(net117),
    .S(_0888_),
    .X(_1695_));
 sky130_fd_sc_hd__o21a_1 _4057_ (.A1(_0901_),
    .A2(_1695_),
    .B1(_0674_),
    .X(_1696_));
 sky130_fd_sc_hd__o211a_1 _4058_ (.A1(net86),
    .A2(_0858_),
    .B1(_0894_),
    .C1(_1168_),
    .X(_1697_));
 sky130_fd_sc_hd__a311o_1 _4059_ (.A1(_0832_),
    .A2(_1437_),
    .A3(_1032_),
    .B1(_1696_),
    .C1(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__o22a_1 _4060_ (.A1(_0879_),
    .A2(_1689_),
    .B1(_1694_),
    .B2(_1698_),
    .X(_1699_));
 sky130_fd_sc_hd__xnor2_2 _4061_ (.A(\u0.E[6] ),
    .B(_1699_),
    .Y(_1700_));
 sky130_fd_sc_hd__buf_2 _4062_ (.A(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__a21boi_1 _4063_ (.A1(_1662_),
    .A2(_1688_),
    .B1_N(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__o21ai_1 _4064_ (.A1(_1662_),
    .A2(_1688_),
    .B1(_1702_),
    .Y(_1703_));
 sky130_fd_sc_hd__o211ai_4 _4065_ (.A1(_1674_),
    .A2(_1675_),
    .B1(_1686_),
    .C1(_1687_),
    .Y(_1704_));
 sky130_fd_sc_hd__a211o_2 _4066_ (.A1(_1686_),
    .A2(_1687_),
    .B1(_1674_),
    .C1(_1675_),
    .X(_1705_));
 sky130_fd_sc_hd__xnor2_4 _4067_ (.A(\u0.E[9] ),
    .B(_1661_),
    .Y(_1706_));
 sky130_fd_sc_hd__a21o_1 _4068_ (.A1(_1704_),
    .A2(_1705_),
    .B1(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__o211a_1 _4069_ (.A1(_1674_),
    .A2(_1675_),
    .B1(_1686_),
    .C1(_1687_),
    .X(_1708_));
 sky130_fd_sc_hd__or3b_1 _4070_ (.A(_1662_),
    .B(_1708_),
    .C_N(_1705_),
    .X(_1709_));
 sky130_fd_sc_hd__a21o_1 _4071_ (.A1(_1707_),
    .A2(_1709_),
    .B1(_1701_),
    .X(_1710_));
 sky130_fd_sc_hd__and3_1 _4072_ (.A(_0947_),
    .B(_1086_),
    .C(_1129_),
    .X(_1711_));
 sky130_fd_sc_hd__and3_1 _4073_ (.A(_0899_),
    .B(_1121_),
    .C(_1132_),
    .X(_1712_));
 sky130_fd_sc_hd__and3_1 _4074_ (.A(_0891_),
    .B(_1067_),
    .C(_1122_),
    .X(_1713_));
 sky130_fd_sc_hd__and3_1 _4075_ (.A(_0866_),
    .B(_1168_),
    .C(_1033_),
    .X(_1714_));
 sky130_fd_sc_hd__and3_1 _4076_ (.A(_0860_),
    .B(_1128_),
    .C(_1091_),
    .X(_1715_));
 sky130_fd_sc_hd__and3_1 _4077_ (.A(_0825_),
    .B(_1114_),
    .C(_1130_),
    .X(_1716_));
 sky130_fd_sc_hd__and3_1 _4078_ (.A(_0893_),
    .B(_1094_),
    .C(_1120_),
    .X(_1717_));
 sky130_fd_sc_hd__or4_1 _4079_ (.A(_1714_),
    .B(_1715_),
    .C(_1716_),
    .D(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__or4_1 _4080_ (.A(_1711_),
    .B(_1712_),
    .C(_1713_),
    .D(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__a31o_1 _4081_ (.A1(_0807_),
    .A2(_1034_),
    .A3(_1490_),
    .B1(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__xnor2_2 _4082_ (.A(\u0.E[12] ),
    .B(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__buf_2 _4083_ (.A(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__a21o_1 _4084_ (.A1(_1703_),
    .A2(_1710_),
    .B1(_1722_),
    .X(_1723_));
 sky130_fd_sc_hd__inv_2 _4085_ (.A(_1464_),
    .Y(\u0.E[5] ));
 sky130_fd_sc_hd__and3_1 _4086_ (.A(_0853_),
    .B(_1046_),
    .C(_1423_),
    .X(_1724_));
 sky130_fd_sc_hd__and3_1 _4087_ (.A(_0819_),
    .B(_1037_),
    .C(_1419_),
    .X(_1725_));
 sky130_fd_sc_hd__a311o_1 _4088_ (.A1(_0992_),
    .A2(_1060_),
    .A3(_1036_),
    .B1(_1724_),
    .C1(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__and3_1 _4089_ (.A(_0862_),
    .B(_1490_),
    .C(_1445_),
    .X(_1727_));
 sky130_fd_sc_hd__and3_1 _4090_ (.A(_0990_),
    .B(_1135_),
    .C(_1042_),
    .X(_1728_));
 sky130_fd_sc_hd__a31o_1 _4091_ (.A1(_0843_),
    .A2(_1052_),
    .A3(_1427_),
    .B1(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__a311o_1 _4092_ (.A1(_0868_),
    .A2(_1049_),
    .A3(_1418_),
    .B1(_1727_),
    .C1(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__clkbuf_4 _4093_ (.A(net86),
    .X(_1731_));
 sky130_fd_sc_hd__o211a_1 _4094_ (.A1(_1731_),
    .A2(_0859_),
    .B1(_0807_),
    .C1(_1128_),
    .X(_1732_));
 sky130_fd_sc_hd__or3_4 _4095_ (.A(_1726_),
    .B(_1730_),
    .C(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__xnor2_4 _4096_ (.A(\u0.E[5] ),
    .B(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _4097_ (.A(_1704_),
    .B(_1705_),
    .Y(_1735_));
 sky130_fd_sc_hd__o211ai_1 _4098_ (.A1(_1701_),
    .A2(_1735_),
    .B1(_1703_),
    .C1(_1722_),
    .Y(_1736_));
 sky130_fd_sc_hd__nand2_2 _4099_ (.A(_1686_),
    .B(_1687_),
    .Y(_1737_));
 sky130_fd_sc_hd__a21oi_1 _4100_ (.A1(_1706_),
    .A2(_1737_),
    .B1(_1700_),
    .Y(_1738_));
 sky130_fd_sc_hd__nand2_1 _4101_ (.A(_1706_),
    .B(_1737_),
    .Y(_1739_));
 sky130_fd_sc_hd__nor2_2 _4102_ (.A(_1674_),
    .B(_1675_),
    .Y(_1740_));
 sky130_fd_sc_hd__nor2_1 _4103_ (.A(_1701_),
    .B(_1740_),
    .Y(_1741_));
 sky130_fd_sc_hd__a21oi_1 _4104_ (.A1(_1704_),
    .A2(_1739_),
    .B1(_1741_),
    .Y(_1742_));
 sky130_fd_sc_hd__a311o_1 _4105_ (.A1(_1704_),
    .A2(_1705_),
    .A3(_1738_),
    .B1(_1742_),
    .C1(_1722_),
    .X(_1743_));
 sky130_fd_sc_hd__xnor2_2 _4106_ (.A(_1662_),
    .B(_1737_),
    .Y(_1744_));
 sky130_fd_sc_hd__or2b_1 _4107_ (.A(_1741_),
    .B_N(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__or3_1 _4108_ (.A(_1701_),
    .B(_1740_),
    .C(_1744_),
    .X(_1746_));
 sky130_fd_sc_hd__a31oi_1 _4109_ (.A1(_1722_),
    .A2(_1745_),
    .A3(_1746_),
    .B1(_1734_),
    .Y(_1747_));
 sky130_fd_sc_hd__a32o_1 _4110_ (.A1(_1723_),
    .A2(_1734_),
    .A3(_1736_),
    .B1(_1743_),
    .B2(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__mux2_1 _4111_ (.A0(net31),
    .A1(net729),
    .S(_1624_),
    .X(_1749_));
 sky130_fd_sc_hd__xnor2_2 _4112_ (.A(_1748_),
    .B(_1749_),
    .Y(\FP[13] ));
 sky130_fd_sc_hd__mux2_1 _4113_ (.A0(\fifo.rd_data[36] ),
    .A1(\FP[13] ),
    .S(_1565_),
    .X(_1750_));
 sky130_fd_sc_hd__a22o_1 _4114_ (.A1(net153),
    .A2(_1589_),
    .B1(_1567_),
    .B2(_1750_),
    .X(_0585_));
 sky130_fd_sc_hd__buf_4 _4115_ (.A(_1302_),
    .X(_1751_));
 sky130_fd_sc_hd__mux2_2 _4116_ (.A0(\fifo.rd_data[35] ),
    .A1(\u0.E[30] ),
    .S(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__a22o_1 _4117_ (.A1(net152),
    .A2(_1589_),
    .B1(_1567_),
    .B2(_1752_),
    .X(_0584_));
 sky130_fd_sc_hd__buf_4 _4118_ (.A(_1305_),
    .X(_1753_));
 sky130_fd_sc_hd__or2_1 _4119_ (.A(_1384_),
    .B(_1647_),
    .X(_1754_));
 sky130_fd_sc_hd__or2_1 _4120_ (.A(_1392_),
    .B(_1637_),
    .X(_1755_));
 sky130_fd_sc_hd__a21o_1 _4121_ (.A1(_1634_),
    .A2(_1755_),
    .B1(_1391_),
    .X(_1756_));
 sky130_fd_sc_hd__a21o_1 _4122_ (.A1(_1632_),
    .A2(_1633_),
    .B1(_1384_),
    .X(_1757_));
 sky130_fd_sc_hd__a211o_1 _4123_ (.A1(_1346_),
    .A2(_1386_),
    .B1(_1333_),
    .C1(_1640_),
    .X(_1758_));
 sky130_fd_sc_hd__a31oi_1 _4124_ (.A1(_1384_),
    .A2(_1755_),
    .A3(_1758_),
    .B1(_1411_),
    .Y(_1759_));
 sky130_fd_sc_hd__a32o_2 _4125_ (.A1(_1411_),
    .A2(_1754_),
    .A3(_1756_),
    .B1(_1757_),
    .B2(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__mux2_1 _4126_ (.A0(net29),
    .A1(\L[21] ),
    .S(_1624_),
    .X(_1761_));
 sky130_fd_sc_hd__xnor2_2 _4127_ (.A(_1760_),
    .B(_1761_),
    .Y(\FP[21] ));
 sky130_fd_sc_hd__mux2_1 _4128_ (.A0(net202),
    .A1(\FP[21] ),
    .S(_1751_),
    .X(_1762_));
 sky130_fd_sc_hd__a22o_1 _4129_ (.A1(net705),
    .A2(_1589_),
    .B1(_1753_),
    .B2(_1762_),
    .X(_0583_));
 sky130_fd_sc_hd__mux2_1 _4130_ (.A0(net394),
    .A1(\u0.E[42] ),
    .S(_1751_),
    .X(_1763_));
 sky130_fd_sc_hd__a22o_1 _4131_ (.A1(net150),
    .A2(_1589_),
    .B1(_1753_),
    .B2(_1763_),
    .X(_0582_));
 sky130_fd_sc_hd__buf_4 _4132_ (.A(_0670_),
    .X(_1764_));
 sky130_fd_sc_hd__a21o_1 _4133_ (.A1(_0962_),
    .A2(_1221_),
    .B1(_0878_),
    .X(_1765_));
 sky130_fd_sc_hd__mux2_1 _4134_ (.A0(net89),
    .A1(net97),
    .S(_0924_),
    .X(_1766_));
 sky130_fd_sc_hd__a32o_1 _4135_ (.A1(_0821_),
    .A2(_0824_),
    .A3(_0916_),
    .B1(_1766_),
    .B2(_0851_),
    .X(_1767_));
 sky130_fd_sc_hd__mux2_1 _4136_ (.A0(net74),
    .A1(net82),
    .S(_0924_),
    .X(_1768_));
 sky130_fd_sc_hd__a32o_1 _4137_ (.A1(_0817_),
    .A2(_0828_),
    .A3(_0937_),
    .B1(_1768_),
    .B2(_0866_),
    .X(_1769_));
 sky130_fd_sc_hd__mux2_1 _4138_ (.A0(net78),
    .A1(net120),
    .S(_0924_),
    .X(_1770_));
 sky130_fd_sc_hd__a32o_1 _4139_ (.A1(_0830_),
    .A2(_0869_),
    .A3(_0938_),
    .B1(_1770_),
    .B2(_0840_),
    .X(_1771_));
 sky130_fd_sc_hd__mux2_1 _4140_ (.A0(net88),
    .A1(net98),
    .S(_0924_),
    .X(_1772_));
 sky130_fd_sc_hd__o21a_1 _4141_ (.A1(_0804_),
    .A2(_1772_),
    .B1(_0673_),
    .X(_1773_));
 sky130_fd_sc_hd__or4_2 _4142_ (.A(_1767_),
    .B(_1769_),
    .C(_1771_),
    .D(_1773_),
    .X(_1774_));
 sky130_fd_sc_hd__a21oi_4 _4143_ (.A1(_1765_),
    .A2(_1774_),
    .B1(\u0.E[35] ),
    .Y(_1775_));
 sky130_fd_sc_hd__and3_2 _4144_ (.A(\u0.E[35] ),
    .B(_1765_),
    .C(_1774_),
    .X(_1776_));
 sky130_fd_sc_hd__nor2_2 _4145_ (.A(_1775_),
    .B(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__mux2_1 _4146_ (.A0(net121),
    .A1(net91),
    .S(_0810_),
    .X(_1778_));
 sky130_fd_sc_hd__o21a_1 _4147_ (.A1(_0804_),
    .A2(_1778_),
    .B1(_0673_),
    .X(_1779_));
 sky130_fd_sc_hd__mux2_1 _4148_ (.A0(net90),
    .A1(net96),
    .S(_0924_),
    .X(_1780_));
 sky130_fd_sc_hd__a32o_1 _4149_ (.A1(_0830_),
    .A2(_0822_),
    .A3(_0827_),
    .B1(_0893_),
    .B2(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(net74),
    .A1(net112),
    .S(_0924_),
    .X(_1782_));
 sky130_fd_sc_hd__a32o_1 _4151_ (.A1(_0828_),
    .A2(_0865_),
    .A3(_0884_),
    .B1(_1782_),
    .B2(_0890_),
    .X(_1783_));
 sky130_fd_sc_hd__mux2_1 _4152_ (.A0(net106),
    .A1(net110),
    .S(_0924_),
    .X(_1784_));
 sky130_fd_sc_hd__a32o_1 _4153_ (.A1(_0850_),
    .A2(_0863_),
    .A3(_0993_),
    .B1(_1784_),
    .B2(_0825_),
    .X(_1785_));
 sky130_fd_sc_hd__or4_2 _4154_ (.A(_1779_),
    .B(_1781_),
    .C(_1783_),
    .D(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__a21o_1 _4155_ (.A1(_0961_),
    .A2(_1220_),
    .B1(_0878_),
    .X(_1787_));
 sky130_fd_sc_hd__a21oi_2 _4156_ (.A1(_1786_),
    .A2(_1787_),
    .B1(\u0.E[34] ),
    .Y(_1788_));
 sky130_fd_sc_hd__and3_2 _4157_ (.A(\u0.E[34] ),
    .B(_1786_),
    .C(_1787_),
    .X(_1789_));
 sky130_fd_sc_hd__or2_1 _4158_ (.A(_1788_),
    .B(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__and3_1 _4159_ (.A(_0844_),
    .B(_0866_),
    .C(_0991_),
    .X(_1791_));
 sky130_fd_sc_hd__a31o_1 _4160_ (.A1(_0822_),
    .A2(_1096_),
    .A3(_0937_),
    .B1(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__and3_1 _4161_ (.A(_0893_),
    .B(_0870_),
    .C(_0948_),
    .X(_1793_));
 sky130_fd_sc_hd__a31o_1 _4162_ (.A1(_0918_),
    .A2(_0854_),
    .A3(_0942_),
    .B1(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__and3_1 _4163_ (.A(_0860_),
    .B(_0884_),
    .C(_0895_),
    .X(_1795_));
 sky130_fd_sc_hd__a31o_1 _4164_ (.A1(_0825_),
    .A2(_0887_),
    .A3(_0996_),
    .B1(_0806_),
    .X(_1796_));
 sky130_fd_sc_hd__a311o_1 _4165_ (.A1(_0913_),
    .A2(_0993_),
    .A3(_0950_),
    .B1(_1795_),
    .C1(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__a21o_1 _4166_ (.A1(_0970_),
    .A2(_1284_),
    .B1(_0878_),
    .X(_1798_));
 sky130_fd_sc_hd__o31a_4 _4167_ (.A1(_1792_),
    .A2(_1794_),
    .A3(_1797_),
    .B1(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__xnor2_4 _4168_ (.A(\u0.E[33] ),
    .B(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__or3_1 _4169_ (.A(_1777_),
    .B(_1790_),
    .C(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__buf_2 _4170_ (.A(_1790_),
    .X(_1802_));
 sky130_fd_sc_hd__o21ai_1 _4171_ (.A1(_1777_),
    .A2(_1802_),
    .B1(_1800_),
    .Y(_1803_));
 sky130_fd_sc_hd__and2_1 _4172_ (.A(_1777_),
    .B(_1790_),
    .X(_1804_));
 sky130_fd_sc_hd__a21o_1 _4173_ (.A1(_1801_),
    .A2(_1803_),
    .B1(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__or2_1 _4174_ (.A(_1777_),
    .B(_1802_),
    .X(_1806_));
 sky130_fd_sc_hd__and3_1 _4175_ (.A(_0861_),
    .B(_0812_),
    .C(_0965_),
    .X(_1807_));
 sky130_fd_sc_hd__and3_1 _4176_ (.A(_0867_),
    .B(_0962_),
    .C(_1289_),
    .X(_1808_));
 sky130_fd_sc_hd__a311o_1 _4177_ (.A1(_0853_),
    .A2(_0953_),
    .A3(_0928_),
    .B1(_1807_),
    .C1(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__and3_1 _4178_ (.A(_0920_),
    .B(_1248_),
    .C(_0975_),
    .X(_1810_));
 sky130_fd_sc_hd__mux2_1 _4179_ (.A0(net74),
    .A1(_0763_),
    .S(_0888_),
    .X(_1811_));
 sky130_fd_sc_hd__a32o_1 _4180_ (.A1(_0899_),
    .A2(_0963_),
    .A3(_0971_),
    .B1(_1811_),
    .B2(_0918_),
    .X(_1812_));
 sky130_fd_sc_hd__a311o_1 _4181_ (.A1(_0842_),
    .A2(_0961_),
    .A3(_1284_),
    .B1(_1810_),
    .C1(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__o211a_1 _4182_ (.A1(_0857_),
    .A2(_0859_),
    .B1(_0806_),
    .C1(_0948_),
    .X(_1814_));
 sky130_fd_sc_hd__nor3_1 _4183_ (.A(_1809_),
    .B(_1813_),
    .C(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__xor2_1 _4184_ (.A(\u0.E[36] ),
    .B(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__clkbuf_4 _4185_ (.A(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__and3_1 _4186_ (.A(_0867_),
    .B(_0971_),
    .C(_0989_),
    .X(_1818_));
 sky130_fd_sc_hd__and3_1 _4187_ (.A(_0920_),
    .B(_0954_),
    .C(_1214_),
    .X(_1819_));
 sky130_fd_sc_hd__a311o_1 _4188_ (.A1(_0832_),
    .A2(_1220_),
    .A3(_1289_),
    .B1(_1818_),
    .C1(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__mux2_1 _4189_ (.A0(_0943_),
    .A1(net112),
    .S(_0834_),
    .X(_1821_));
 sky130_fd_sc_hd__a32o_1 _4190_ (.A1(_0860_),
    .A2(_0881_),
    .A3(_1221_),
    .B1(_1821_),
    .B2(_0894_),
    .X(_1822_));
 sky130_fd_sc_hd__o211a_1 _4191_ (.A1(net67),
    .A2(_0848_),
    .B1(_0852_),
    .C1(_1284_),
    .X(_1823_));
 sky130_fd_sc_hd__a311o_1 _4192_ (.A1(_0891_),
    .A2(_0816_),
    .A3(_0975_),
    .B1(_1822_),
    .C1(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__and3_1 _4193_ (.A(_0822_),
    .B(_0806_),
    .C(_0941_),
    .X(_1825_));
 sky130_fd_sc_hd__nor3_4 _4194_ (.A(_1820_),
    .B(_1824_),
    .C(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__xor2_2 _4195_ (.A(\u0.E[30] ),
    .B(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__xnor2_1 _4196_ (.A(_1817_),
    .B(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__inv_2 _4197_ (.A(_1816_),
    .Y(_1829_));
 sky130_fd_sc_hd__o2bb2a_1 _4198_ (.A1_N(_1806_),
    .A2_N(_1828_),
    .B1(_1829_),
    .B2(_1802_),
    .X(_1830_));
 sky130_fd_sc_hd__nor2_1 _4199_ (.A(_1805_),
    .B(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__o211a_1 _4200_ (.A1(_0880_),
    .A2(_0849_),
    .B1(_0853_),
    .C1(_0816_),
    .X(_1832_));
 sky130_fd_sc_hd__o211a_1 _4201_ (.A1(_1347_),
    .A2(_0849_),
    .B1(_0819_),
    .C1(_0953_),
    .X(_1833_));
 sky130_fd_sc_hd__a311o_1 _4202_ (.A1(_0992_),
    .A2(_0972_),
    .A3(_1193_),
    .B1(_1832_),
    .C1(_1833_),
    .X(_1834_));
 sky130_fd_sc_hd__o211a_1 _4203_ (.A1(_1227_),
    .A2(_0859_),
    .B1(_0868_),
    .C1(_0961_),
    .X(_1835_));
 sky130_fd_sc_hd__and3_1 _4204_ (.A(_0990_),
    .B(_0966_),
    .C(_1243_),
    .X(_1836_));
 sky130_fd_sc_hd__a31o_1 _4205_ (.A1(_0843_),
    .A2(_0962_),
    .A3(_0989_),
    .B1(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__a311o_1 _4206_ (.A1(_0862_),
    .A2(_0970_),
    .A3(_0926_),
    .B1(_1835_),
    .C1(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__o211a_1 _4207_ (.A1(_0847_),
    .A2(_0849_),
    .B1(_0807_),
    .C1(_0884_),
    .X(_1839_));
 sky130_fd_sc_hd__nor3_2 _4208_ (.A(_1834_),
    .B(_1838_),
    .C(_1839_),
    .Y(_1840_));
 sky130_fd_sc_hd__xnor2_4 _4209_ (.A(_0908_),
    .B(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__inv_2 _4210_ (.A(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__a21o_1 _4211_ (.A1(_1805_),
    .A2(_1830_),
    .B1(_1842_),
    .X(_1843_));
 sky130_fd_sc_hd__o22a_1 _4212_ (.A1(_1775_),
    .A2(_1776_),
    .B1(_1788_),
    .B2(_1789_),
    .X(_1844_));
 sky130_fd_sc_hd__or4_4 _4213_ (.A(_1775_),
    .B(_1776_),
    .C(_1788_),
    .D(_1789_),
    .X(_1845_));
 sky130_fd_sc_hd__or3b_1 _4214_ (.A(_1800_),
    .B(_1844_),
    .C_N(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4215_ (.A(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__or2_1 _4216_ (.A(_1775_),
    .B(_1776_),
    .X(_1848_));
 sky130_fd_sc_hd__nand2_1 _4217_ (.A(_1848_),
    .B(_1800_),
    .Y(_1849_));
 sky130_fd_sc_hd__buf_2 _4218_ (.A(_1827_),
    .X(_1850_));
 sky130_fd_sc_hd__a21oi_1 _4219_ (.A1(_1847_),
    .A2(_1849_),
    .B1(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__o22ai_4 _4220_ (.A1(_1775_),
    .A2(_1776_),
    .B1(_1788_),
    .B2(_1789_),
    .Y(_1852_));
 sky130_fd_sc_hd__xor2_4 _4221_ (.A(\u0.E[33] ),
    .B(_1799_),
    .X(_1853_));
 sky130_fd_sc_hd__a21o_1 _4222_ (.A1(_1852_),
    .A2(_1845_),
    .B1(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__and3_1 _4223_ (.A(_1850_),
    .B(_1847_),
    .C(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__a21oi_1 _4224_ (.A1(_1777_),
    .A2(_1853_),
    .B1(_1850_),
    .Y(_1856_));
 sky130_fd_sc_hd__a21o_1 _4225_ (.A1(_1777_),
    .A2(_1853_),
    .B1(_1844_),
    .X(_1857_));
 sky130_fd_sc_hd__a221o_1 _4226_ (.A1(_1849_),
    .A2(_1856_),
    .B1(_1857_),
    .B2(_1850_),
    .C1(_1829_),
    .X(_1858_));
 sky130_fd_sc_hd__o31ai_1 _4227_ (.A1(_1817_),
    .A2(_1851_),
    .A3(_1855_),
    .B1(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__o22a_1 _4228_ (.A1(_1831_),
    .A2(_1843_),
    .B1(_1859_),
    .B2(_1841_),
    .X(_1860_));
 sky130_fd_sc_hd__mux2_1 _4229_ (.A0(net27),
    .A1(net685),
    .S(_1030_),
    .X(_1861_));
 sky130_fd_sc_hd__xor2_1 _4230_ (.A(_1860_),
    .B(_1861_),
    .X(\FP[29] ));
 sky130_fd_sc_hd__mux2_1 _4231_ (.A0(\fifo.rd_data[32] ),
    .A1(\FP[29] ),
    .S(_1751_),
    .X(_1862_));
 sky130_fd_sc_hd__a22o_1 _4232_ (.A1(net149),
    .A2(_1764_),
    .B1(_1753_),
    .B2(_1862_),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _4233_ (.A0(net683),
    .A1(\u0.E[5] ),
    .S(_1751_),
    .X(_1863_));
 sky130_fd_sc_hd__a22o_1 _4234_ (.A1(net694),
    .A2(_1764_),
    .B1(_1753_),
    .B2(_1863_),
    .X(_0580_));
 sky130_fd_sc_hd__nor2_1 _4235_ (.A(_1853_),
    .B(_1827_),
    .Y(_1864_));
 sky130_fd_sc_hd__xnor2_4 _4236_ (.A(\u0.E[30] ),
    .B(_1826_),
    .Y(_1865_));
 sky130_fd_sc_hd__a21oi_1 _4237_ (.A1(_1777_),
    .A2(_1802_),
    .B1(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__nor2_1 _4238_ (.A(_1802_),
    .B(_1800_),
    .Y(_1867_));
 sky130_fd_sc_hd__a221o_1 _4239_ (.A1(_1802_),
    .A2(_1864_),
    .B1(_1866_),
    .B2(_1849_),
    .C1(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__o21ai_1 _4240_ (.A1(_1802_),
    .A2(_1865_),
    .B1(_1800_),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_1 _4241_ (.A(_1852_),
    .B(_1845_),
    .Y(_1870_));
 sky130_fd_sc_hd__a221o_1 _4242_ (.A1(_1845_),
    .A2(_1864_),
    .B1(_1869_),
    .B2(_1870_),
    .C1(_1829_),
    .X(_1871_));
 sky130_fd_sc_hd__a21bo_1 _4243_ (.A1(_1829_),
    .A2(_1868_),
    .B1_N(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(_1864_),
    .A1(_1850_),
    .S(_1804_),
    .X(_1873_));
 sky130_fd_sc_hd__nand2_1 _4245_ (.A(_1817_),
    .B(_1847_),
    .Y(_1874_));
 sky130_fd_sc_hd__a21oi_1 _4246_ (.A1(_1802_),
    .A2(_1800_),
    .B1(_1865_),
    .Y(_1875_));
 sky130_fd_sc_hd__or2_1 _4247_ (.A(_1802_),
    .B(_1853_),
    .X(_1876_));
 sky130_fd_sc_hd__a221o_1 _4248_ (.A1(_1847_),
    .A2(_1875_),
    .B1(_1876_),
    .B2(_1856_),
    .C1(_1817_),
    .X(_1877_));
 sky130_fd_sc_hd__o21ai_1 _4249_ (.A1(_1873_),
    .A2(_1874_),
    .B1(_1877_),
    .Y(_1878_));
 sky130_fd_sc_hd__mux2_1 _4250_ (.A0(_1872_),
    .A1(_1878_),
    .S(_1841_),
    .X(_1879_));
 sky130_fd_sc_hd__mux2_1 _4251_ (.A0(net25),
    .A1(\L[4] ),
    .S(_1030_),
    .X(_1880_));
 sky130_fd_sc_hd__xor2_2 _4252_ (.A(_1879_),
    .B(_1880_),
    .X(\FP[4] ));
 sky130_fd_sc_hd__mux2_1 _4253_ (.A0(net669),
    .A1(\FP[4] ),
    .S(_1751_),
    .X(_1881_));
 sky130_fd_sc_hd__a22o_1 _4254_ (.A1(net147),
    .A2(_1764_),
    .B1(_1753_),
    .B2(_1881_),
    .X(_0579_));
 sky130_fd_sc_hd__inv_2 _4255_ (.A(_1078_),
    .Y(\u0.E[17] ));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(\fifo.rd_data[29] ),
    .A1(\u0.E[17] ),
    .S(_1751_),
    .X(_1882_));
 sky130_fd_sc_hd__a22o_1 _4257_ (.A1(net145),
    .A2(_1764_),
    .B1(_1753_),
    .B2(_1882_),
    .X(_0578_));
 sky130_fd_sc_hd__a221o_1 _4258_ (.A1(_1235_),
    .A2(_1266_),
    .B1(_1270_),
    .B2(_1280_),
    .C1(_1269_),
    .X(_1883_));
 sky130_fd_sc_hd__a21o_1 _4259_ (.A1(_1264_),
    .A2(_1883_),
    .B1(_1205_),
    .X(_1884_));
 sky130_fd_sc_hd__and3_1 _4260_ (.A(_1235_),
    .B(_1266_),
    .C(_1267_),
    .X(_1885_));
 sky130_fd_sc_hd__a2111o_1 _4261_ (.A1(_1218_),
    .A2(_1263_),
    .B1(_1599_),
    .C1(_1885_),
    .D1(_1205_),
    .X(_1886_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(_1275_),
    .A1(_1263_),
    .S(_1218_),
    .X(_1887_));
 sky130_fd_sc_hd__a21oi_1 _4263_ (.A1(_1205_),
    .A2(_1887_),
    .B1(_1294_),
    .Y(_1888_));
 sky130_fd_sc_hd__a32o_1 _4264_ (.A1(_1294_),
    .A2(_1273_),
    .A3(_1884_),
    .B1(_1886_),
    .B2(_1888_),
    .X(_1889_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(net22),
    .A1(\L[12] ),
    .S(_1030_),
    .X(_1890_));
 sky130_fd_sc_hd__xor2_2 _4266_ (.A(_1889_),
    .B(_1890_),
    .X(\FP[12] ));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(net672),
    .A1(\FP[12] ),
    .S(_1751_),
    .X(_1891_));
 sky130_fd_sc_hd__a22o_1 _4268_ (.A1(net725),
    .A2(_1764_),
    .B1(_1753_),
    .B2(_1891_),
    .X(_0577_));
 sky130_fd_sc_hd__inv_2 _4269_ (.A(_0908_),
    .Y(\u0.E[29] ));
 sky130_fd_sc_hd__mux2_1 _4270_ (.A0(net279),
    .A1(\u0.E[29] ),
    .S(_1751_),
    .X(_1892_));
 sky130_fd_sc_hd__a22o_1 _4271_ (.A1(net143),
    .A2(_1764_),
    .B1(_1753_),
    .B2(_1892_),
    .X(_0576_));
 sky130_fd_sc_hd__and3_1 _4272_ (.A(_0862_),
    .B(_1122_),
    .C(_1033_),
    .X(_1893_));
 sky130_fd_sc_hd__a31o_1 _4273_ (.A1(_0992_),
    .A2(_1129_),
    .A3(_1125_),
    .B1(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__and3_1 _4274_ (.A(_0842_),
    .B(_1114_),
    .C(_1068_),
    .X(_1895_));
 sky130_fd_sc_hd__a31o_1 _4275_ (.A1(_0819_),
    .A2(_1072_),
    .A3(_1091_),
    .B1(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__o211a_1 _4276_ (.A1(_1518_),
    .A2(_0859_),
    .B1(_0990_),
    .C1(_1120_),
    .X(_1897_));
 sky130_fd_sc_hd__a311o_1 _4277_ (.A1(_0868_),
    .A2(_1064_),
    .A3(_1128_),
    .B1(_1896_),
    .C1(_1897_),
    .X(_1898_));
 sky130_fd_sc_hd__a311o_1 _4278_ (.A1(_0853_),
    .A2(_1522_),
    .A3(_1132_),
    .B1(_1894_),
    .C1(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__a31oi_4 _4279_ (.A1(_0808_),
    .A2(_1054_),
    .A3(_1418_),
    .B1(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__xnor2_4 _4280_ (.A(\u0.E[17] ),
    .B(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__a21o_1 _4281_ (.A1(_1111_),
    .A2(_1046_),
    .B1(_0878_),
    .X(_1902_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(net83),
    .A1(net93),
    .S(_0814_),
    .X(_1903_));
 sky130_fd_sc_hd__o21a_1 _4283_ (.A1(_0877_),
    .A2(_1903_),
    .B1(_0876_),
    .X(_1904_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(net102),
    .A1(net109),
    .S(_0896_),
    .X(_1905_));
 sky130_fd_sc_hd__a32o_1 _4285_ (.A1(_0890_),
    .A2(_1090_),
    .A3(_1129_),
    .B1(_1905_),
    .B2(_0866_),
    .X(_1906_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(net118),
    .A1(net86),
    .S(_0833_),
    .X(_1907_));
 sky130_fd_sc_hd__a32o_1 _4287_ (.A1(_0825_),
    .A2(_1064_),
    .A3(_1125_),
    .B1(_1907_),
    .B2(_0851_),
    .X(_1908_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(net68),
    .A1(net108),
    .S(_0896_),
    .X(_1909_));
 sky130_fd_sc_hd__a32o_1 _4289_ (.A1(_0893_),
    .A2(_1477_),
    .A3(_1033_),
    .B1(_1909_),
    .B2(_0831_),
    .X(_1910_));
 sky130_fd_sc_hd__or4_1 _4290_ (.A(_1904_),
    .B(_1906_),
    .C(_1908_),
    .D(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__a21o_1 _4291_ (.A1(_1902_),
    .A2(_1911_),
    .B1(_1321_),
    .X(_1912_));
 sky130_fd_sc_hd__nand3_2 _4292_ (.A(_1321_),
    .B(_1902_),
    .C(_1911_),
    .Y(_1913_));
 sky130_fd_sc_hd__nand2_1 _4293_ (.A(_1912_),
    .B(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hd__a21o_1 _4294_ (.A1(_1068_),
    .A2(_1094_),
    .B1(_0955_),
    .X(_1915_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(net92),
    .A1(_0734_),
    .S(_1035_),
    .X(_1916_));
 sky130_fd_sc_hd__o21a_1 _4296_ (.A1(_0877_),
    .A2(_1916_),
    .B1(_0876_),
    .X(_1917_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(net85),
    .A1(_0727_),
    .S(_0988_),
    .X(_1918_));
 sky130_fd_sc_hd__a32o_1 _4298_ (.A1(_1089_),
    .A2(_1045_),
    .A3(_1427_),
    .B1(_1918_),
    .B2(_0818_),
    .X(_1919_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(net86),
    .A1(net107),
    .S(_0988_),
    .X(_1920_));
 sky130_fd_sc_hd__a32o_1 _4300_ (.A1(_1096_),
    .A2(_1041_),
    .A3(_1419_),
    .B1(_1920_),
    .B2(_1074_),
    .X(_1921_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(net76),
    .A1(net117),
    .S(_1035_),
    .X(_1922_));
 sky130_fd_sc_hd__a32o_1 _4302_ (.A1(_0841_),
    .A2(_1034_),
    .A3(_1418_),
    .B1(_1922_),
    .B2(_0831_),
    .X(_1923_));
 sky130_fd_sc_hd__or4_4 _4303_ (.A(_1917_),
    .B(_1919_),
    .C(_1921_),
    .D(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__a21oi_2 _4304_ (.A1(_1915_),
    .A2(_1924_),
    .B1(\u0.E[23] ),
    .Y(_1925_));
 sky130_fd_sc_hd__and3_1 _4305_ (.A(\u0.E[23] ),
    .B(_1915_),
    .C(_1924_),
    .X(_1926_));
 sky130_fd_sc_hd__a21o_1 _4306_ (.A1(_1522_),
    .A2(_1086_),
    .B1(_0879_),
    .X(_1927_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(net84),
    .A1(_0738_),
    .S(_0888_),
    .X(_1928_));
 sky130_fd_sc_hd__o21a_1 _4308_ (.A1(_0901_),
    .A2(_1928_),
    .B1(_0674_),
    .X(_1929_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(net119),
    .A1(net68),
    .S(_0897_),
    .X(_1930_));
 sky130_fd_sc_hd__a32o_1 _4310_ (.A1(_0867_),
    .A2(_1039_),
    .A3(_1135_),
    .B1(_1930_),
    .B2(_0918_),
    .X(_1931_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(_0719_),
    .A1(net116),
    .S(_0897_),
    .X(_1932_));
 sky130_fd_sc_hd__a32o_1 _4312_ (.A1(_0920_),
    .A2(_1049_),
    .A3(_1036_),
    .B1(_1932_),
    .B2(_0852_),
    .X(_1933_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(_0721_),
    .A1(_0741_),
    .S(_0897_),
    .X(_1934_));
 sky130_fd_sc_hd__a32o_1 _4314_ (.A1(_0913_),
    .A2(_1037_),
    .A3(_1042_),
    .B1(_1934_),
    .B2(_0894_),
    .X(_1935_));
 sky130_fd_sc_hd__or4_4 _4315_ (.A(_1929_),
    .B(_1931_),
    .C(_1933_),
    .D(_1935_),
    .X(_1936_));
 sky130_fd_sc_hd__a21o_1 _4316_ (.A1(_1927_),
    .A2(_1936_),
    .B1(\u0.E[21] ),
    .X(_1937_));
 sky130_fd_sc_hd__nand3_2 _4317_ (.A(\u0.E[21] ),
    .B(_1927_),
    .C(_1936_),
    .Y(_1938_));
 sky130_fd_sc_hd__o211a_1 _4318_ (.A1(_1925_),
    .A2(_1926_),
    .B1(_1937_),
    .C1(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__a21o_1 _4319_ (.A1(_1915_),
    .A2(_1924_),
    .B1(\u0.E[23] ),
    .X(_1940_));
 sky130_fd_sc_hd__nand3_1 _4320_ (.A(\u0.E[23] ),
    .B(_1915_),
    .C(_1924_),
    .Y(_1941_));
 sky130_fd_sc_hd__a22o_1 _4321_ (.A1(_1912_),
    .A2(_1913_),
    .B1(_1940_),
    .B2(_1941_),
    .X(_1942_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(_1937_),
    .B(_1938_),
    .Y(_1943_));
 sky130_fd_sc_hd__a22o_1 _4323_ (.A1(_1914_),
    .A2(_1939_),
    .B1(_1942_),
    .B2(_1943_),
    .X(_1944_));
 sky130_fd_sc_hd__and4_1 _4324_ (.A(_1912_),
    .B(_1913_),
    .C(_1940_),
    .D(_1941_),
    .X(_1945_));
 sky130_fd_sc_hd__and3_1 _4325_ (.A(_0913_),
    .B(_1135_),
    .C(_1419_),
    .X(_1946_));
 sky130_fd_sc_hd__o211a_1 _4326_ (.A1(net76),
    .A2(_0815_),
    .B1(_0852_),
    .C1(_1445_),
    .X(_1947_));
 sky130_fd_sc_hd__a311o_1 _4327_ (.A1(_0974_),
    .A2(_1111_),
    .A3(_1042_),
    .B1(_1946_),
    .C1(_1947_),
    .X(_1948_));
 sky130_fd_sc_hd__and3_1 _4328_ (.A(_0860_),
    .B(_1423_),
    .C(_1427_),
    .X(_1949_));
 sky130_fd_sc_hd__and3_1 _4329_ (.A(_0890_),
    .B(_1105_),
    .C(_1036_),
    .X(_1950_));
 sky130_fd_sc_hd__and3_1 _4330_ (.A(_0841_),
    .B(_1082_),
    .C(_1490_),
    .X(_1951_));
 sky130_fd_sc_hd__and3_1 _4331_ (.A(_1074_),
    .B(_1060_),
    .C(_1418_),
    .X(_1952_));
 sky130_fd_sc_hd__or4_1 _4332_ (.A(_1949_),
    .B(_1950_),
    .C(_1951_),
    .D(_1952_),
    .X(_1953_));
 sky130_fd_sc_hd__clkbuf_4 _4333_ (.A(net117),
    .X(_1954_));
 sky130_fd_sc_hd__o211a_1 _4334_ (.A1(_1954_),
    .A2(_0858_),
    .B1(_0806_),
    .C1(_1120_),
    .X(_1955_));
 sky130_fd_sc_hd__nor3_1 _4335_ (.A(_1948_),
    .B(_1953_),
    .C(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__xnor2_2 _4336_ (.A(\u0.E[18] ),
    .B(_1956_),
    .Y(_1957_));
 sky130_fd_sc_hd__and2b_1 _4337_ (.A_N(_1945_),
    .B(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__nand2_1 _4338_ (.A(_1940_),
    .B(_1941_),
    .Y(_1959_));
 sky130_fd_sc_hd__or2b_1 _4339_ (.A(_1959_),
    .B_N(_1943_),
    .X(_1960_));
 sky130_fd_sc_hd__buf_2 _4340_ (.A(_1957_),
    .X(_1961_));
 sky130_fd_sc_hd__a21oi_1 _4341_ (.A1(_1914_),
    .A2(_1939_),
    .B1(_1961_),
    .Y(_1962_));
 sky130_fd_sc_hd__a22o_1 _4342_ (.A1(_1944_),
    .A2(_1958_),
    .B1(_1960_),
    .B2(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__a211oi_4 _4343_ (.A1(_1937_),
    .A2(_1938_),
    .B1(_1925_),
    .C1(_1926_),
    .Y(_1964_));
 sky130_fd_sc_hd__and2_1 _4344_ (.A(_1912_),
    .B(_1913_),
    .X(_1965_));
 sky130_fd_sc_hd__clkbuf_2 _4345_ (.A(_1965_),
    .X(_1966_));
 sky130_fd_sc_hd__a2bb2o_1 _4346_ (.A1_N(_1945_),
    .A2_N(_1943_),
    .B1(_1964_),
    .B2(_1966_),
    .X(_1967_));
 sky130_fd_sc_hd__a211o_1 _4347_ (.A1(_1912_),
    .A2(_1913_),
    .B1(_1925_),
    .C1(_1926_),
    .X(_1968_));
 sky130_fd_sc_hd__a21boi_2 _4348_ (.A1(_1966_),
    .A2(_1959_),
    .B1_N(_1961_),
    .Y(_1969_));
 sky130_fd_sc_hd__a2bb2o_1 _4349_ (.A1_N(_1961_),
    .A2_N(_1967_),
    .B1(_1968_),
    .B2(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__and3_1 _4350_ (.A(_0853_),
    .B(_1090_),
    .C(_1094_),
    .X(_1971_));
 sky130_fd_sc_hd__o211a_1 _4351_ (.A1(_1954_),
    .A2(_0859_),
    .B1(_1168_),
    .C1(_0992_),
    .X(_1972_));
 sky130_fd_sc_hd__o211a_1 _4352_ (.A1(_1731_),
    .A2(_0859_),
    .B1(_0819_),
    .C1(_1130_),
    .X(_1973_));
 sky130_fd_sc_hd__and3_1 _4353_ (.A(_0974_),
    .B(_1477_),
    .C(_1121_),
    .X(_1974_));
 sky130_fd_sc_hd__and3_1 _4354_ (.A(_0841_),
    .B(_1437_),
    .C(_1086_),
    .X(_1975_));
 sky130_fd_sc_hd__a31o_1 _4355_ (.A1(_0826_),
    .A2(_1666_),
    .A3(_1067_),
    .B1(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__a311o_1 _4356_ (.A1(_0862_),
    .A2(_1071_),
    .A3(_1032_),
    .B1(_1974_),
    .C1(_1976_),
    .X(_1977_));
 sky130_fd_sc_hd__or4_2 _4357_ (.A(_1971_),
    .B(_1972_),
    .C(_1973_),
    .D(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__a31oi_4 _4358_ (.A1(_0808_),
    .A2(_1053_),
    .A3(_1419_),
    .B1(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__xor2_4 _4359_ (.A(\u0.E[24] ),
    .B(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__mux2_1 _4360_ (.A0(_1963_),
    .A1(_1970_),
    .S(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__xnor2_4 _4361_ (.A(\u0.E[24] ),
    .B(_1979_),
    .Y(_1982_));
 sky130_fd_sc_hd__a21o_1 _4362_ (.A1(_1966_),
    .A2(_1964_),
    .B1(_1961_),
    .X(_1983_));
 sky130_fd_sc_hd__nor2_1 _4363_ (.A(_1966_),
    .B(_1964_),
    .Y(_1984_));
 sky130_fd_sc_hd__a2bb2o_1 _4364_ (.A1_N(_1983_),
    .A2_N(_1984_),
    .B1(_1961_),
    .B2(_1944_),
    .X(_1985_));
 sky130_fd_sc_hd__nand2_1 _4365_ (.A(_1982_),
    .B(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__nand2_1 _4366_ (.A(_1943_),
    .B(_1968_),
    .Y(_1987_));
 sky130_fd_sc_hd__nor2_1 _4367_ (.A(_1939_),
    .B(_1961_),
    .Y(_1988_));
 sky130_fd_sc_hd__a22o_1 _4368_ (.A1(_1969_),
    .A2(_1987_),
    .B1(_1988_),
    .B2(_1968_),
    .X(_1989_));
 sky130_fd_sc_hd__a21oi_1 _4369_ (.A1(_1980_),
    .A2(_1989_),
    .B1(_1901_),
    .Y(_1990_));
 sky130_fd_sc_hd__a22o_1 _4370_ (.A1(_1901_),
    .A2(_1981_),
    .B1(_1986_),
    .B2(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__mux2_1 _4371_ (.A0(net20),
    .A1(net190),
    .S(_1624_),
    .X(_1992_));
 sky130_fd_sc_hd__xnor2_1 _4372_ (.A(_1991_),
    .B(_1992_),
    .Y(\FP[20] ));
 sky130_fd_sc_hd__mux2_1 _4373_ (.A0(net194),
    .A1(\FP[20] ),
    .S(_1751_),
    .X(_1993_));
 sky130_fd_sc_hd__a22o_1 _4374_ (.A1(net142),
    .A2(_1764_),
    .B1(_1753_),
    .B2(_1993_),
    .X(_0575_));
 sky130_fd_sc_hd__clkbuf_4 _4375_ (.A(_1302_),
    .X(_1994_));
 sky130_fd_sc_hd__mux2_1 _4376_ (.A0(net712),
    .A1(\u0.E[41] ),
    .S(_1994_),
    .X(_1995_));
 sky130_fd_sc_hd__a22o_1 _4377_ (.A1(net141),
    .A2(_1764_),
    .B1(_1753_),
    .B2(_1995_),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_4 _4378_ (.A(_1305_),
    .X(_1996_));
 sky130_fd_sc_hd__xnor2_1 _4379_ (.A(_1700_),
    .B(_1705_),
    .Y(_1997_));
 sky130_fd_sc_hd__o21a_1 _4380_ (.A1(_1706_),
    .A2(_1997_),
    .B1(_1709_),
    .X(_1998_));
 sky130_fd_sc_hd__nor2_1 _4381_ (.A(_1722_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__inv_2 _4382_ (.A(_1721_),
    .Y(_2000_));
 sky130_fd_sc_hd__inv_2 _4383_ (.A(_1701_),
    .Y(_2001_));
 sky130_fd_sc_hd__and3_1 _4384_ (.A(_1700_),
    .B(_1704_),
    .C(_1705_),
    .X(_2002_));
 sky130_fd_sc_hd__a21oi_1 _4385_ (.A1(_2001_),
    .A2(_1744_),
    .B1(_2002_),
    .Y(_2003_));
 sky130_fd_sc_hd__o21ai_1 _4386_ (.A1(_2000_),
    .A2(_2003_),
    .B1(_1734_),
    .Y(_2004_));
 sky130_fd_sc_hd__a21oi_1 _4387_ (.A1(_1688_),
    .A2(_1738_),
    .B1(_2002_),
    .Y(_2005_));
 sky130_fd_sc_hd__mux2_1 _4388_ (.A0(_1998_),
    .A1(_2005_),
    .S(_1722_),
    .X(_2006_));
 sky130_fd_sc_hd__o22a_1 _4389_ (.A1(_1999_),
    .A2(_2004_),
    .B1(_2006_),
    .B2(_1734_),
    .X(_2007_));
 sky130_fd_sc_hd__mux2_1 _4390_ (.A0(net18),
    .A1(net727),
    .S(_1624_),
    .X(_2008_));
 sky130_fd_sc_hd__xnor2_1 _4391_ (.A(_2007_),
    .B(_2008_),
    .Y(\FP[28] ));
 sky130_fd_sc_hd__mux2_1 _4392_ (.A0(net687),
    .A1(\FP[28] ),
    .S(_1994_),
    .X(_2009_));
 sky130_fd_sc_hd__a22o_1 _4393_ (.A1(net140),
    .A2(_1764_),
    .B1(_1996_),
    .B2(_2009_),
    .X(_0573_));
 sky130_fd_sc_hd__inv_2 _4394_ (.A(_1448_),
    .Y(\u0.E[4] ));
 sky130_fd_sc_hd__mux2_1 _4395_ (.A0(\fifo.rd_data[23] ),
    .A1(\u0.E[4] ),
    .S(_1994_),
    .X(_2010_));
 sky130_fd_sc_hd__a22o_1 _4396_ (.A1(net139),
    .A2(_1764_),
    .B1(_1996_),
    .B2(_2010_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_4 _4397_ (.A(_0669_),
    .X(_2011_));
 sky130_fd_sc_hd__a211o_1 _4398_ (.A1(_0983_),
    .A2(_1572_),
    .B1(_1019_),
    .C1(_0984_),
    .X(_2012_));
 sky130_fd_sc_hd__and3_1 _4399_ (.A(_1007_),
    .B(_1008_),
    .C(_0959_),
    .X(_2013_));
 sky130_fd_sc_hd__mux2_1 _4400_ (.A0(_0936_),
    .A1(_1010_),
    .S(_1009_),
    .X(_2014_));
 sky130_fd_sc_hd__o221a_1 _4401_ (.A1(_1573_),
    .A2(_2013_),
    .B1(_2014_),
    .B2(_0982_),
    .C1(_1019_),
    .X(_2015_));
 sky130_fd_sc_hd__nor2_1 _4402_ (.A(_0875_),
    .B(_2015_),
    .Y(_2016_));
 sky130_fd_sc_hd__or3_1 _4403_ (.A(_0982_),
    .B(_1011_),
    .C(_1025_),
    .X(_2017_));
 sky130_fd_sc_hd__and3_1 _4404_ (.A(_1007_),
    .B(_1008_),
    .C(_0936_),
    .X(_2018_));
 sky130_fd_sc_hd__o21ai_1 _4405_ (.A1(_2018_),
    .A2(_1022_),
    .B1(_0983_),
    .Y(_2019_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(_0935_),
    .B(_1017_),
    .Y(_2020_));
 sky130_fd_sc_hd__o221a_1 _4407_ (.A1(_0982_),
    .A2(_2020_),
    .B1(_1573_),
    .B2(_2013_),
    .C1(_1019_),
    .X(_2021_));
 sky130_fd_sc_hd__a31o_1 _4408_ (.A1(_1005_),
    .A2(_2017_),
    .A3(_2019_),
    .B1(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__a22oi_2 _4409_ (.A1(_2012_),
    .A2(_2016_),
    .B1(_2022_),
    .B2(_0875_),
    .Y(_2023_));
 sky130_fd_sc_hd__mux2_1 _4410_ (.A0(net16),
    .A1(net709),
    .S(_1413_),
    .X(_2024_));
 sky130_fd_sc_hd__xor2_1 _4411_ (.A(_2023_),
    .B(_2024_),
    .X(\FP[3] ));
 sky130_fd_sc_hd__mux2_1 _4412_ (.A0(net666),
    .A1(\FP[3] ),
    .S(_1994_),
    .X(_2025_));
 sky130_fd_sc_hd__a22o_1 _4413_ (.A1(net699),
    .A2(_2011_),
    .B1(_1996_),
    .B2(_2025_),
    .X(_0571_));
 sky130_fd_sc_hd__inv_2 _4414_ (.A(_1100_),
    .Y(\u0.E[16] ));
 sky130_fd_sc_hd__mux2_1 _4415_ (.A0(net662),
    .A1(\u0.E[16] ),
    .S(_1994_),
    .X(_2026_));
 sky130_fd_sc_hd__a22o_1 _4416_ (.A1(net707),
    .A2(_2011_),
    .B1(_1996_),
    .B2(_2026_),
    .X(_0570_));
 sky130_fd_sc_hd__or2_1 _4417_ (.A(_1802_),
    .B(_1800_),
    .X(_2027_));
 sky130_fd_sc_hd__a21oi_1 _4418_ (.A1(_2027_),
    .A2(_1854_),
    .B1(_1850_),
    .Y(_2028_));
 sky130_fd_sc_hd__o21a_1 _4419_ (.A1(_1855_),
    .A2(_2028_),
    .B1(_1817_),
    .X(_2029_));
 sky130_fd_sc_hd__a311o_1 _4420_ (.A1(_1800_),
    .A2(_1852_),
    .A3(_1845_),
    .B1(_1867_),
    .C1(_1865_),
    .X(_2030_));
 sky130_fd_sc_hd__mux2_1 _4421_ (.A0(_1790_),
    .A1(_1800_),
    .S(_1777_),
    .X(_2031_));
 sky130_fd_sc_hd__or2_1 _4422_ (.A(_1850_),
    .B(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__a31o_1 _4423_ (.A1(_1829_),
    .A2(_2030_),
    .A3(_2032_),
    .B1(_1841_),
    .X(_2033_));
 sky130_fd_sc_hd__a21oi_1 _4424_ (.A1(_1847_),
    .A2(_1854_),
    .B1(_1850_),
    .Y(_2034_));
 sky130_fd_sc_hd__a21o_1 _4425_ (.A1(_1850_),
    .A2(_2031_),
    .B1(_1817_),
    .X(_2035_));
 sky130_fd_sc_hd__a21oi_1 _4426_ (.A1(_1847_),
    .A2(_1876_),
    .B1(_1865_),
    .Y(_2036_));
 sky130_fd_sc_hd__a31o_1 _4427_ (.A1(_1801_),
    .A2(_1803_),
    .A3(_1865_),
    .B1(_1829_),
    .X(_2037_));
 sky130_fd_sc_hd__o22a_1 _4428_ (.A1(_2034_),
    .A2(_2035_),
    .B1(_2036_),
    .B2(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__o22a_1 _4429_ (.A1(_2029_),
    .A2(_2033_),
    .B1(_2038_),
    .B2(_1842_),
    .X(_2039_));
 sky130_fd_sc_hd__mux2_1 _4430_ (.A0(net14),
    .A1(net700),
    .S(_1413_),
    .X(_2040_));
 sky130_fd_sc_hd__xor2_1 _4431_ (.A(_2039_),
    .B(_2040_),
    .X(\FP[11] ));
 sky130_fd_sc_hd__mux2_1 _4432_ (.A0(\fifo.rd_data[20] ),
    .A1(\FP[11] ),
    .S(_1994_),
    .X(_2041_));
 sky130_fd_sc_hd__a22o_1 _4433_ (.A1(net136),
    .A2(_2011_),
    .B1(_1996_),
    .B2(_2041_),
    .X(_0569_));
 sky130_fd_sc_hd__inv_2 _4434_ (.A(_0932_),
    .Y(\u0.E[28] ));
 sky130_fd_sc_hd__mux2_1 _4435_ (.A0(net192),
    .A1(\u0.E[28] ),
    .S(_1994_),
    .X(_2042_));
 sky130_fd_sc_hd__a22o_1 _4436_ (.A1(net134),
    .A2(_2011_),
    .B1(_1996_),
    .B2(_2042_),
    .X(_0568_));
 sky130_fd_sc_hd__nor2_1 _4437_ (.A(_1817_),
    .B(_1865_),
    .Y(_2043_));
 sky130_fd_sc_hd__and2_1 _4438_ (.A(_1845_),
    .B(_1849_),
    .X(_2044_));
 sky130_fd_sc_hd__mux2_1 _4439_ (.A0(_1828_),
    .A1(_2043_),
    .S(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__o21a_1 _4440_ (.A1(_1853_),
    .A2(_1844_),
    .B1(_1845_),
    .X(_2046_));
 sky130_fd_sc_hd__a31o_1 _4441_ (.A1(_1817_),
    .A2(_1865_),
    .A3(_2046_),
    .B1(_1841_),
    .X(_2047_));
 sky130_fd_sc_hd__or2_1 _4442_ (.A(_1870_),
    .B(_1875_),
    .X(_2048_));
 sky130_fd_sc_hd__a21oi_1 _4443_ (.A1(_1853_),
    .A2(_1866_),
    .B1(_1817_),
    .Y(_2049_));
 sky130_fd_sc_hd__mux2_1 _4444_ (.A0(_1848_),
    .A1(_1852_),
    .S(_1853_),
    .X(_2050_));
 sky130_fd_sc_hd__a22o_1 _4445_ (.A1(_1870_),
    .A2(_1856_),
    .B1(_2050_),
    .B2(_1850_),
    .X(_2051_));
 sky130_fd_sc_hd__a22o_1 _4446_ (.A1(_2048_),
    .A2(_2049_),
    .B1(_2051_),
    .B2(_1817_),
    .X(_2052_));
 sky130_fd_sc_hd__a2bb2o_1 _4447_ (.A1_N(_2045_),
    .A2_N(_2047_),
    .B1(_2052_),
    .B2(_1841_),
    .X(_2053_));
 sky130_fd_sc_hd__mux2_1 _4448_ (.A0(net11),
    .A1(net723),
    .S(_1624_),
    .X(_2054_));
 sky130_fd_sc_hd__xnor2_1 _4449_ (.A(_2053_),
    .B(_2054_),
    .Y(\FP[19] ));
 sky130_fd_sc_hd__mux2_1 _4450_ (.A0(net218),
    .A1(\FP[19] ),
    .S(_1994_),
    .X(_2055_));
 sky130_fd_sc_hd__a22o_1 _4451_ (.A1(net133),
    .A2(_2011_),
    .B1(_1996_),
    .B2(_2055_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _4452_ (.A0(net405),
    .A1(\u0.E[40] ),
    .S(_1994_),
    .X(_2056_));
 sky130_fd_sc_hd__a22o_1 _4453_ (.A1(net132),
    .A2(_2011_),
    .B1(_1996_),
    .B2(_2056_),
    .X(_0566_));
 sky130_fd_sc_hd__nor3_1 _4454_ (.A(_1333_),
    .B(_1637_),
    .C(_1640_),
    .Y(_2057_));
 sky130_fd_sc_hd__o21ai_1 _4455_ (.A1(_1641_),
    .A2(_2057_),
    .B1(_1384_),
    .Y(_2058_));
 sky130_fd_sc_hd__or2b_1 _4456_ (.A(_1392_),
    .B_N(_1387_),
    .X(_2059_));
 sky130_fd_sc_hd__a21boi_1 _4457_ (.A1(_1635_),
    .A2(_2059_),
    .B1_N(_1411_),
    .Y(_2060_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(_1346_),
    .A1(_1371_),
    .S(_1358_),
    .X(_2061_));
 sky130_fd_sc_hd__mux2_1 _4459_ (.A0(_2061_),
    .A1(_1398_),
    .S(_1645_),
    .X(_2062_));
 sky130_fd_sc_hd__nand2_1 _4460_ (.A(_1391_),
    .B(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__o21ba_1 _4461_ (.A1(_1391_),
    .A2(_2062_),
    .B1_N(_1411_),
    .X(_2064_));
 sky130_fd_sc_hd__a22o_2 _4462_ (.A1(_2058_),
    .A2(_2060_),
    .B1(_2063_),
    .B2(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__mux2_1 _4463_ (.A0(net9),
    .A1(net697),
    .S(_1624_),
    .X(_2066_));
 sky130_fd_sc_hd__xnor2_1 _4464_ (.A(_2065_),
    .B(_2066_),
    .Y(\FP[27] ));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(net381),
    .A1(\FP[27] ),
    .S(_1994_),
    .X(_2067_));
 sky130_fd_sc_hd__a22o_1 _4466_ (.A1(net686),
    .A2(_2011_),
    .B1(_1996_),
    .B2(_2067_),
    .X(_0565_));
 sky130_fd_sc_hd__buf_4 _4467_ (.A(_1301_),
    .X(_2068_));
 sky130_fd_sc_hd__mux2_1 _4468_ (.A0(net561),
    .A1(\u0.E[3] ),
    .S(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__a22o_1 _4469_ (.A1(net130),
    .A2(_2011_),
    .B1(_1996_),
    .B2(_2069_),
    .X(_0564_));
 sky130_fd_sc_hd__buf_4 _4470_ (.A(_0678_),
    .X(_2070_));
 sky130_fd_sc_hd__nand2_1 _4471_ (.A(_1706_),
    .B(_1704_),
    .Y(_2071_));
 sky130_fd_sc_hd__and3_1 _4472_ (.A(_1701_),
    .B(_1707_),
    .C(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__a21oi_1 _4473_ (.A1(_1707_),
    .A2(_2071_),
    .B1(_1701_),
    .Y(_2073_));
 sky130_fd_sc_hd__or3_1 _4474_ (.A(_2000_),
    .B(_2072_),
    .C(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__nand2_1 _4475_ (.A(_1706_),
    .B(_1740_),
    .Y(_2075_));
 sky130_fd_sc_hd__nand2_1 _4476_ (.A(_1662_),
    .B(_1708_),
    .Y(_2076_));
 sky130_fd_sc_hd__a221o_1 _4477_ (.A1(_2002_),
    .A2(_2075_),
    .B1(_2076_),
    .B2(_1738_),
    .C1(_1721_),
    .X(_2077_));
 sky130_fd_sc_hd__and2_1 _4478_ (.A(_1734_),
    .B(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__nand2_1 _4479_ (.A(_1662_),
    .B(_1740_),
    .Y(_2079_));
 sky130_fd_sc_hd__o211a_1 _4480_ (.A1(_1740_),
    .A2(_1744_),
    .B1(_2079_),
    .C1(_1701_),
    .X(_2080_));
 sky130_fd_sc_hd__nor2_1 _4481_ (.A(_1700_),
    .B(_1708_),
    .Y(_2081_));
 sky130_fd_sc_hd__a21o_1 _4482_ (.A1(_2075_),
    .A2(_2081_),
    .B1(_1722_),
    .X(_2082_));
 sky130_fd_sc_hd__nand2_1 _4483_ (.A(_1662_),
    .B(_1705_),
    .Y(_2083_));
 sky130_fd_sc_hd__o221a_1 _4484_ (.A1(_1662_),
    .A2(_1997_),
    .B1(_2081_),
    .B2(_2083_),
    .C1(_1722_),
    .X(_2084_));
 sky130_fd_sc_hd__o21ba_1 _4485_ (.A1(_2080_),
    .A2(_2082_),
    .B1_N(_2084_),
    .X(_2085_));
 sky130_fd_sc_hd__o2bb2a_1 _4486_ (.A1_N(_2074_),
    .A2_N(_2078_),
    .B1(_2085_),
    .B2(_1734_),
    .X(_2086_));
 sky130_fd_sc_hd__mux2_1 _4487_ (.A0(net7),
    .A1(net726),
    .S(_1413_),
    .X(_2087_));
 sky130_fd_sc_hd__xor2_1 _4488_ (.A(_2086_),
    .B(_2087_),
    .X(\FP[2] ));
 sky130_fd_sc_hd__mux2_1 _4489_ (.A0(net433),
    .A1(\FP[2] ),
    .S(_2068_),
    .X(_2088_));
 sky130_fd_sc_hd__a22o_1 _4490_ (.A1(net129),
    .A2(_2011_),
    .B1(_2070_),
    .B2(_2088_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _4491_ (.A0(net488),
    .A1(\u0.E[15] ),
    .S(_2068_),
    .X(_2089_));
 sky130_fd_sc_hd__a22o_1 _4492_ (.A1(net128),
    .A2(_2011_),
    .B1(_2070_),
    .B2(_2089_),
    .X(_0562_));
 sky130_fd_sc_hd__buf_4 _4493_ (.A(_0669_),
    .X(_2090_));
 sky130_fd_sc_hd__or2_1 _4494_ (.A(_1914_),
    .B(_1939_),
    .X(_2091_));
 sky130_fd_sc_hd__a22o_1 _4495_ (.A1(_1961_),
    .A2(_1967_),
    .B1(_2091_),
    .B2(_1962_),
    .X(_2092_));
 sky130_fd_sc_hd__or2_1 _4496_ (.A(_1982_),
    .B(_2092_),
    .X(_2093_));
 sky130_fd_sc_hd__a21oi_1 _4497_ (.A1(_1966_),
    .A2(_1959_),
    .B1(_1964_),
    .Y(_2094_));
 sky130_fd_sc_hd__a2bb2o_1 _4498_ (.A1_N(_1961_),
    .A2_N(_2094_),
    .B1(_1987_),
    .B2(_1969_),
    .X(_2095_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(_1982_),
    .B(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__nand2_1 _4500_ (.A(_1966_),
    .B(_1964_),
    .Y(_2097_));
 sky130_fd_sc_hd__a32oi_2 _4501_ (.A1(_1942_),
    .A2(_1961_),
    .A3(_1967_),
    .B1(_1988_),
    .B2(_2097_),
    .Y(_2098_));
 sky130_fd_sc_hd__or2_1 _4502_ (.A(_1982_),
    .B(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__o2bb2a_1 _4503_ (.A1_N(_1968_),
    .A2_N(_1969_),
    .B1(_1944_),
    .B2(_1961_),
    .X(_2100_));
 sky130_fd_sc_hd__o21ba_1 _4504_ (.A1(_1980_),
    .A2(_2100_),
    .B1_N(_1901_),
    .X(_2101_));
 sky130_fd_sc_hd__a32o_1 _4505_ (.A1(_1901_),
    .A2(_2093_),
    .A3(_2096_),
    .B1(_2099_),
    .B2(_2101_),
    .X(_2102_));
 sky130_fd_sc_hd__mux2_1 _4506_ (.A0(net5),
    .A1(net721),
    .S(_1624_),
    .X(_2103_));
 sky130_fd_sc_hd__xnor2_1 _4507_ (.A(_2102_),
    .B(_2103_),
    .Y(\FP[10] ));
 sky130_fd_sc_hd__mux2_1 _4508_ (.A0(net207),
    .A1(\FP[10] ),
    .S(_2068_),
    .X(_2104_));
 sky130_fd_sc_hd__a22o_1 _4509_ (.A1(net127),
    .A2(_2090_),
    .B1(_2070_),
    .B2(_2104_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _4510_ (.A0(\fifo.rd_data[11] ),
    .A1(\u0.E[27] ),
    .S(_2068_),
    .X(_2105_));
 sky130_fd_sc_hd__a22o_1 _4511_ (.A1(net126),
    .A2(_2090_),
    .B1(_2070_),
    .B2(_2105_),
    .X(_0560_));
 sky130_fd_sc_hd__nand2_1 _4512_ (.A(_2001_),
    .B(_1744_),
    .Y(_2106_));
 sky130_fd_sc_hd__a21o_1 _4513_ (.A1(_1707_),
    .A2(_2075_),
    .B1(_2001_),
    .X(_2107_));
 sky130_fd_sc_hd__a21oi_1 _4514_ (.A1(_2106_),
    .A2(_2107_),
    .B1(_1722_),
    .Y(_2108_));
 sky130_fd_sc_hd__o211a_1 _4515_ (.A1(_1662_),
    .A2(_1737_),
    .B1(_1705_),
    .C1(_2001_),
    .X(_2109_));
 sky130_fd_sc_hd__a211oi_1 _4516_ (.A1(_1701_),
    .A2(_1740_),
    .B1(_2109_),
    .C1(_2000_),
    .Y(_2110_));
 sky130_fd_sc_hd__o31a_1 _4517_ (.A1(_2001_),
    .A2(_1662_),
    .A3(_1735_),
    .B1(_2079_),
    .X(_2111_));
 sky130_fd_sc_hd__a21oi_1 _4518_ (.A1(_1746_),
    .A2(_2111_),
    .B1(_2000_),
    .Y(_2112_));
 sky130_fd_sc_hd__o21ai_1 _4519_ (.A1(_1706_),
    .A2(_1737_),
    .B1(_1705_),
    .Y(_2113_));
 sky130_fd_sc_hd__nor2_1 _4520_ (.A(_2001_),
    .B(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__a21o_1 _4521_ (.A1(_2001_),
    .A2(_2113_),
    .B1(_1722_),
    .X(_2115_));
 sky130_fd_sc_hd__o21ai_1 _4522_ (.A1(_2114_),
    .A2(_2115_),
    .B1(_1734_),
    .Y(_2116_));
 sky130_fd_sc_hd__o32a_2 _4523_ (.A1(_1734_),
    .A2(_2108_),
    .A3(_2110_),
    .B1(_2112_),
    .B2(_2116_),
    .X(_2117_));
 sky130_fd_sc_hd__mux2_1 _4524_ (.A0(net3),
    .A1(net711),
    .S(_1413_),
    .X(_2118_));
 sky130_fd_sc_hd__xor2_1 _4525_ (.A(_2117_),
    .B(_2118_),
    .X(\FP[18] ));
 sky130_fd_sc_hd__mux2_1 _4526_ (.A0(\fifo.rd_data[10] ),
    .A1(\FP[18] ),
    .S(_2068_),
    .X(_2119_));
 sky130_fd_sc_hd__a22o_1 _4527_ (.A1(net125),
    .A2(_2090_),
    .B1(_2070_),
    .B2(_2119_),
    .X(_0559_));
 sky130_fd_sc_hd__mux2_1 _4528_ (.A0(\fifo.rd_data[9] ),
    .A1(\u0.E[39] ),
    .S(_2068_),
    .X(_2120_));
 sky130_fd_sc_hd__a22o_1 _4529_ (.A1(net717),
    .A2(_2090_),
    .B1(_2070_),
    .B2(_2120_),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _4530_ (.A(_1980_),
    .B(_1963_),
    .Y(_2121_));
 sky130_fd_sc_hd__or2_1 _4531_ (.A(_1980_),
    .B(_1970_),
    .X(_2122_));
 sky130_fd_sc_hd__or2_1 _4532_ (.A(_1982_),
    .B(_1985_),
    .X(_2123_));
 sky130_fd_sc_hd__a21oi_1 _4533_ (.A1(_1982_),
    .A2(_1989_),
    .B1(_1901_),
    .Y(_2124_));
 sky130_fd_sc_hd__a32o_1 _4534_ (.A1(_1901_),
    .A2(_2121_),
    .A3(_2122_),
    .B1(_2123_),
    .B2(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__mux2_1 _4535_ (.A0(net64),
    .A1(net434),
    .S(_1624_),
    .X(_2126_));
 sky130_fd_sc_hd__xnor2_1 _4536_ (.A(_2125_),
    .B(_2126_),
    .Y(\FP[26] ));
 sky130_fd_sc_hd__mux2_1 _4537_ (.A0(net502),
    .A1(\FP[26] ),
    .S(_2068_),
    .X(_2127_));
 sky130_fd_sc_hd__a22o_1 _4538_ (.A1(net186),
    .A2(_2090_),
    .B1(_2070_),
    .B2(_2127_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _4539_ (.A0(\fifo.rd_data[7] ),
    .A1(\u0.E[2] ),
    .S(_2068_),
    .X(_2128_));
 sky130_fd_sc_hd__a22o_1 _4540_ (.A1(net185),
    .A2(_2090_),
    .B1(_2070_),
    .B2(_2128_),
    .X(_0556_));
 sky130_fd_sc_hd__or2_1 _4541_ (.A(_1980_),
    .B(_2098_),
    .X(_2129_));
 sky130_fd_sc_hd__a21oi_1 _4542_ (.A1(_1980_),
    .A2(_2100_),
    .B1(_1901_),
    .Y(_2130_));
 sky130_fd_sc_hd__mux2_1 _4543_ (.A0(_2095_),
    .A1(_2092_),
    .S(_1982_),
    .X(_2131_));
 sky130_fd_sc_hd__a22o_1 _4544_ (.A1(_2129_),
    .A2(_2130_),
    .B1(_2131_),
    .B2(_1901_),
    .X(_2132_));
 sky130_fd_sc_hd__mux2_1 _4545_ (.A0(net62),
    .A1(net714),
    .S(_1624_),
    .X(_2133_));
 sky130_fd_sc_hd__xnor2_1 _4546_ (.A(_2132_),
    .B(_2133_),
    .Y(\FP[1] ));
 sky130_fd_sc_hd__mux2_1 _4547_ (.A0(\fifo.rd_data[6] ),
    .A1(\FP[1] ),
    .S(_2068_),
    .X(_2134_));
 sky130_fd_sc_hd__a22o_1 _4548_ (.A1(net184),
    .A2(_2090_),
    .B1(_2070_),
    .B2(_2134_),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _4549_ (.A0(net542),
    .A1(\u0.E[12] ),
    .S(_1302_),
    .X(_2135_));
 sky130_fd_sc_hd__a22o_1 _4550_ (.A1(net704),
    .A2(_2090_),
    .B1(_2070_),
    .B2(_2135_),
    .X(_0554_));
 sky130_fd_sc_hd__a21oi_1 _4551_ (.A1(_1486_),
    .A2(_1487_),
    .B1(_1537_),
    .Y(_2136_));
 sky130_fd_sc_hd__o21bai_1 _4552_ (.A1(_1434_),
    .A2(_1451_),
    .B1_N(_1535_),
    .Y(_2137_));
 sky130_fd_sc_hd__mux2_1 _4553_ (.A0(_2136_),
    .A1(_2137_),
    .S(_1483_),
    .X(_2138_));
 sky130_fd_sc_hd__or2_1 _4554_ (.A(_1535_),
    .B(_1537_),
    .X(_2139_));
 sky130_fd_sc_hd__a211oi_1 _4555_ (.A1(_1486_),
    .A2(_1487_),
    .B1(_1537_),
    .C1(_1480_),
    .Y(_2140_));
 sky130_fd_sc_hd__a21o_1 _4556_ (.A1(_1480_),
    .A2(_2139_),
    .B1(_2140_),
    .X(_2141_));
 sky130_fd_sc_hd__a21o_1 _4557_ (.A1(_1434_),
    .A2(_1486_),
    .B1(_1480_),
    .X(_2142_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_1452_),
    .B(_1487_),
    .Y(_2143_));
 sky130_fd_sc_hd__xnor2_1 _4559_ (.A(_2142_),
    .B(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__a21o_1 _4560_ (.A1(_1486_),
    .A2(_1487_),
    .B1(_1434_),
    .X(_2145_));
 sky130_fd_sc_hd__and2b_1 _4561_ (.A_N(_1484_),
    .B(_1538_),
    .X(_2146_));
 sky130_fd_sc_hd__a31oi_1 _4562_ (.A1(_1483_),
    .A2(_1509_),
    .A3(_2145_),
    .B1(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__mux4_1 _4563_ (.A0(_2138_),
    .A1(_2141_),
    .A2(_2144_),
    .A3(_2147_),
    .S0(_1516_),
    .S1(_1534_),
    .X(_2148_));
 sky130_fd_sc_hd__mux2_1 _4564_ (.A0(net46),
    .A1(net715),
    .S(_0905_),
    .X(_2149_));
 sky130_fd_sc_hd__xnor2_1 _4565_ (.A(_2148_),
    .B(_2149_),
    .Y(\FP[9] ));
 sky130_fd_sc_hd__mux2_1 _4566_ (.A0(net734),
    .A1(\FP[9] ),
    .S(_1302_),
    .X(_2150_));
 sky130_fd_sc_hd__a22o_1 _4567_ (.A1(net168),
    .A2(_2090_),
    .B1(_1305_),
    .B2(_2150_),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _4568_ (.A0(net604),
    .A1(\u0.E[24] ),
    .S(_1302_),
    .X(_2151_));
 sky130_fd_sc_hd__a22o_1 _4569_ (.A1(net157),
    .A2(_2090_),
    .B1(_1305_),
    .B2(_2151_),
    .X(_0552_));
 sky130_fd_sc_hd__a211oi_1 _4570_ (.A1(_1480_),
    .A2(_2137_),
    .B1(_2140_),
    .C1(_1516_),
    .Y(_2152_));
 sky130_fd_sc_hd__a21o_1 _4571_ (.A1(_1509_),
    .A2(_1512_),
    .B1(_1480_),
    .X(_2153_));
 sky130_fd_sc_hd__o31ai_1 _4572_ (.A1(_1434_),
    .A2(_1486_),
    .A3(_1487_),
    .B1(_1538_),
    .Y(_2154_));
 sky130_fd_sc_hd__a31o_1 _4573_ (.A1(_1516_),
    .A2(_2153_),
    .A3(_2154_),
    .B1(_1529_),
    .X(_2155_));
 sky130_fd_sc_hd__a21oi_1 _4574_ (.A1(_1452_),
    .A2(_1469_),
    .B1(_1483_),
    .Y(_2156_));
 sky130_fd_sc_hd__o31ai_1 _4575_ (.A1(_1480_),
    .A2(_1535_),
    .A3(_1536_),
    .B1(_1516_),
    .Y(_2157_));
 sky130_fd_sc_hd__o32a_1 _4576_ (.A1(_1483_),
    .A2(_1484_),
    .A3(_1488_),
    .B1(_2142_),
    .B2(_1537_),
    .X(_2158_));
 sky130_fd_sc_hd__o22a_1 _4577_ (.A1(_2156_),
    .A2(_2157_),
    .B1(_2158_),
    .B2(_1516_),
    .X(_2159_));
 sky130_fd_sc_hd__o22a_1 _4578_ (.A1(_2152_),
    .A2(_2155_),
    .B1(_2159_),
    .B2(_1534_),
    .X(_2160_));
 sky130_fd_sc_hd__mux2_1 _4579_ (.A0(net24),
    .A1(net191),
    .S(_1413_),
    .X(_2161_));
 sky130_fd_sc_hd__xor2_1 _4580_ (.A(_2160_),
    .B(_2161_),
    .X(\FP[17] ));
 sky130_fd_sc_hd__mux2_1 _4581_ (.A0(\fifo.rd_data[2] ),
    .A1(\FP[17] ),
    .S(_1302_),
    .X(_2162_));
 sky130_fd_sc_hd__a22o_1 _4582_ (.A1(net146),
    .A2(_0670_),
    .B1(_1305_),
    .B2(_2162_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _4583_ (.A0(net420),
    .A1(\u0.E[36] ),
    .S(_1302_),
    .X(_2163_));
 sky130_fd_sc_hd__a22o_1 _4584_ (.A1(net135),
    .A2(_0670_),
    .B1(_1305_),
    .B2(_2163_),
    .X(_0550_));
 sky130_fd_sc_hd__nor2_1 _4585_ (.A(_1010_),
    .B(_1018_),
    .Y(_2164_));
 sky130_fd_sc_hd__o311a_1 _4586_ (.A1(_0983_),
    .A2(_1025_),
    .A3(_2164_),
    .B1(_1026_),
    .C1(_0875_),
    .X(_2165_));
 sky130_fd_sc_hd__o21a_1 _4587_ (.A1(_0936_),
    .A2(_1010_),
    .B1(_0935_),
    .X(_2166_));
 sky130_fd_sc_hd__o221a_1 _4588_ (.A1(_2020_),
    .A2(_1573_),
    .B1(_2166_),
    .B2(_0987_),
    .C1(_1570_),
    .X(_2167_));
 sky130_fd_sc_hd__nor2_1 _4589_ (.A(_0983_),
    .B(_0960_),
    .Y(_2168_));
 sky130_fd_sc_hd__o211a_1 _4590_ (.A1(_1009_),
    .A2(_0936_),
    .B1(_1577_),
    .C1(_0982_),
    .X(_2169_));
 sky130_fd_sc_hd__o21a_1 _4591_ (.A1(_2168_),
    .A2(_2169_),
    .B1(_0875_),
    .X(_2170_));
 sky130_fd_sc_hd__a22o_1 _4592_ (.A1(_0985_),
    .A2(_1571_),
    .B1(_1575_),
    .B2(_0987_),
    .X(_2171_));
 sky130_fd_sc_hd__a21o_1 _4593_ (.A1(_1570_),
    .A2(_2171_),
    .B1(_1019_),
    .X(_2172_));
 sky130_fd_sc_hd__o32a_2 _4594_ (.A1(_1005_),
    .A2(_2165_),
    .A3(_2167_),
    .B1(_2170_),
    .B2(_2172_),
    .X(_2173_));
 sky130_fd_sc_hd__mux2_1 _4595_ (.A0(net2),
    .A1(\L[25] ),
    .S(_0905_),
    .X(_2174_));
 sky130_fd_sc_hd__xnor2_2 _4596_ (.A(_2173_),
    .B(_2174_),
    .Y(\FP[25] ));
 sky130_fd_sc_hd__mux2_1 _4597_ (.A0(net222),
    .A1(\FP[25] ),
    .S(_1302_),
    .X(_2175_));
 sky130_fd_sc_hd__a22o_1 _4598_ (.A1(net124),
    .A2(_0670_),
    .B1(_1305_),
    .B2(_2175_),
    .X(_0549_));
 sky130_fd_sc_hd__and3b_4 _4599_ (.A_N(\fifo.fifo_empty ),
    .B(_0767_),
    .C(_0793_),
    .X(_2176_));
 sky130_fd_sc_hd__clkbuf_8 _4600_ (.A(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__nand2_1 _4601_ (.A(_0785_),
    .B(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__nor2_1 _4602_ (.A(_0783_),
    .B(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__xnor2_1 _4603_ (.A(_0781_),
    .B(_2179_),
    .Y(_0380_));
 sky130_fd_sc_hd__xnor2_1 _4604_ (.A(_0789_),
    .B(_2178_),
    .Y(_0379_));
 sky130_fd_sc_hd__buf_4 _4605_ (.A(_2176_),
    .X(_2180_));
 sky130_fd_sc_hd__xor2_1 _4606_ (.A(_0785_),
    .B(_2180_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_1 _4607_ (.A(_1606_),
    .B(_1607_),
    .Y(\FP[22] ));
 sky130_fd_sc_hd__and2_1 _4608_ (.A(_1315_),
    .B(_1316_),
    .X(_2181_));
 sky130_fd_sc_hd__clkbuf_1 _4609_ (.A(_2181_),
    .X(\FP[7] ));
 sky130_fd_sc_hd__and3_1 _4610_ (.A(\fifo.wr_ptr[2] ),
    .B(_0788_),
    .C(_0770_),
    .X(_2182_));
 sky130_fd_sc_hd__clkbuf_8 _4611_ (.A(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__buf_4 _4612_ (.A(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__mux2_1 _4613_ (.A0(net453),
    .A1(_1347_),
    .S(_2184_),
    .X(_2185_));
 sky130_fd_sc_hd__clkbuf_1 _4614_ (.A(_2185_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _4615_ (.A0(net547),
    .A1(_0943_),
    .S(_2184_),
    .X(_2186_));
 sky130_fd_sc_hd__clkbuf_1 _4616_ (.A(_2186_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _4617_ (.A0(net314),
    .A1(_0845_),
    .S(_2184_),
    .X(_2187_));
 sky130_fd_sc_hd__clkbuf_1 _4618_ (.A(_2187_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _4619_ (.A0(net357),
    .A1(_0705_),
    .S(_2184_),
    .X(_2188_));
 sky130_fd_sc_hd__clkbuf_1 _4620_ (.A(_2188_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _4621_ (.A0(net307),
    .A1(_0703_),
    .S(_2184_),
    .X(_2189_));
 sky130_fd_sc_hd__clkbuf_1 _4622_ (.A(_2189_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _4623_ (.A0(net351),
    .A1(_0702_),
    .S(_2184_),
    .X(_2190_));
 sky130_fd_sc_hd__clkbuf_1 _4624_ (.A(_2190_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _4625_ (.A0(net204),
    .A1(_1048_),
    .S(_2184_),
    .X(_2191_));
 sky130_fd_sc_hd__clkbuf_1 _4626_ (.A(_2191_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _4627_ (.A0(net648),
    .A1(_0847_),
    .S(_2184_),
    .X(_2192_));
 sky130_fd_sc_hd__clkbuf_1 _4628_ (.A(_2192_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _4629_ (.A0(net224),
    .A1(_0713_),
    .S(_2184_),
    .X(_2193_));
 sky130_fd_sc_hd__clkbuf_1 _4630_ (.A(_2193_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _4631_ (.A0(net450),
    .A1(_0714_),
    .S(_2184_),
    .X(_2194_));
 sky130_fd_sc_hd__clkbuf_1 _4632_ (.A(_2194_),
    .X(_0632_));
 sky130_fd_sc_hd__buf_4 _4633_ (.A(_2183_),
    .X(_2195_));
 sky130_fd_sc_hd__mux2_1 _4634_ (.A0(net354),
    .A1(_1518_),
    .S(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__clkbuf_1 _4635_ (.A(_2196_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _4636_ (.A0(net484),
    .A1(_0715_),
    .S(_2195_),
    .X(_2197_));
 sky130_fd_sc_hd__clkbuf_1 _4637_ (.A(_2197_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _4638_ (.A0(net629),
    .A1(_0708_),
    .S(_2195_),
    .X(_2198_));
 sky130_fd_sc_hd__clkbuf_1 _4639_ (.A(_2198_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _4640_ (.A0(net652),
    .A1(_0711_),
    .S(_2195_),
    .X(_2199_));
 sky130_fd_sc_hd__clkbuf_1 _4641_ (.A(_2199_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _4642_ (.A0(net520),
    .A1(_0710_),
    .S(_2195_),
    .X(_2200_));
 sky130_fd_sc_hd__clkbuf_1 _4643_ (.A(_2200_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _4644_ (.A0(net344),
    .A1(_0709_),
    .S(_2195_),
    .X(_2201_));
 sky130_fd_sc_hd__clkbuf_1 _4645_ (.A(_2201_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _4646_ (.A0(net442),
    .A1(_0880_),
    .S(_2195_),
    .X(_2202_));
 sky130_fd_sc_hd__clkbuf_1 _4647_ (.A(_2202_),
    .X(_0639_));
 sky130_fd_sc_hd__mux2_1 _4648_ (.A0(net286),
    .A1(_0718_),
    .S(_2195_),
    .X(_2203_));
 sky130_fd_sc_hd__clkbuf_1 _4649_ (.A(_2203_),
    .X(_0640_));
 sky130_fd_sc_hd__mux2_1 _4650_ (.A0(net512),
    .A1(_1493_),
    .S(_2195_),
    .X(_2204_));
 sky130_fd_sc_hd__clkbuf_1 _4651_ (.A(_2204_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_1 _4652_ (.A0(net379),
    .A1(_0719_),
    .S(_2195_),
    .X(_2205_));
 sky130_fd_sc_hd__clkbuf_1 _4653_ (.A(_2205_),
    .X(_0642_));
 sky130_fd_sc_hd__buf_4 _4654_ (.A(_2183_),
    .X(_2206_));
 sky130_fd_sc_hd__mux2_1 _4655_ (.A0(net611),
    .A1(_0721_),
    .S(_2206_),
    .X(_2207_));
 sky130_fd_sc_hd__clkbuf_1 _4656_ (.A(_2207_),
    .X(_0643_));
 sky130_fd_sc_hd__mux2_1 _4657_ (.A0(net197),
    .A1(_0724_),
    .S(_2206_),
    .X(_2208_));
 sky130_fd_sc_hd__clkbuf_1 _4658_ (.A(_2208_),
    .X(_0644_));
 sky130_fd_sc_hd__mux2_1 _4659_ (.A0(net401),
    .A1(_0723_),
    .S(_2206_),
    .X(_2209_));
 sky130_fd_sc_hd__clkbuf_1 _4660_ (.A(_2209_),
    .X(_0645_));
 sky130_fd_sc_hd__mux2_1 _4661_ (.A0(net356),
    .A1(_0722_),
    .S(_2206_),
    .X(_2210_));
 sky130_fd_sc_hd__clkbuf_1 _4662_ (.A(_2210_),
    .X(_0646_));
 sky130_fd_sc_hd__mux2_1 _4663_ (.A0(net303),
    .A1(_0750_),
    .S(_2206_),
    .X(_2211_));
 sky130_fd_sc_hd__clkbuf_1 _4664_ (.A(_2211_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2_1 _4665_ (.A0(net501),
    .A1(_0752_),
    .S(_2206_),
    .X(_2212_));
 sky130_fd_sc_hd__clkbuf_1 _4666_ (.A(_2212_),
    .X(_0648_));
 sky130_fd_sc_hd__mux2_1 _4667_ (.A0(net429),
    .A1(_0751_),
    .S(_2206_),
    .X(_2213_));
 sky130_fd_sc_hd__clkbuf_1 _4668_ (.A(_2213_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _4669_ (.A0(net508),
    .A1(_1731_),
    .S(_2206_),
    .X(_2214_));
 sky130_fd_sc_hd__clkbuf_1 _4670_ (.A(_2214_),
    .X(_0650_));
 sky130_fd_sc_hd__mux2_1 _4671_ (.A0(net315),
    .A1(_0746_),
    .S(_2206_),
    .X(_2215_));
 sky130_fd_sc_hd__clkbuf_1 _4672_ (.A(_2215_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _4673_ (.A0(net569),
    .A1(_0748_),
    .S(_2206_),
    .X(_2216_));
 sky130_fd_sc_hd__clkbuf_1 _4674_ (.A(_2216_),
    .X(_0652_));
 sky130_fd_sc_hd__buf_4 _4675_ (.A(_2183_),
    .X(_2217_));
 sky130_fd_sc_hd__mux2_1 _4676_ (.A0(net447),
    .A1(_0857_),
    .S(_2217_),
    .X(_2218_));
 sky130_fd_sc_hd__clkbuf_1 _4677_ (.A(_2218_),
    .X(_0653_));
 sky130_fd_sc_hd__mux2_1 _4678_ (.A0(net288),
    .A1(_0747_),
    .S(_2217_),
    .X(_2219_));
 sky130_fd_sc_hd__clkbuf_1 _4679_ (.A(_2219_),
    .X(_0654_));
 sky130_fd_sc_hd__mux2_1 _4680_ (.A0(net306),
    .A1(_0755_),
    .S(_2217_),
    .X(_2220_));
 sky130_fd_sc_hd__clkbuf_1 _4681_ (.A(_2220_),
    .X(_0655_));
 sky130_fd_sc_hd__mux2_1 _4682_ (.A0(net349),
    .A1(_0756_),
    .S(_2217_),
    .X(_2221_));
 sky130_fd_sc_hd__clkbuf_1 _4683_ (.A(_2221_),
    .X(_0656_));
 sky130_fd_sc_hd__mux2_1 _4684_ (.A0(net563),
    .A1(_0757_),
    .S(_2217_),
    .X(_2222_));
 sky130_fd_sc_hd__clkbuf_1 _4685_ (.A(_2222_),
    .X(_0657_));
 sky130_fd_sc_hd__mux2_1 _4686_ (.A0(net201),
    .A1(_0758_),
    .S(_2217_),
    .X(_2223_));
 sky130_fd_sc_hd__clkbuf_1 _4687_ (.A(_2223_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _4688_ (.A0(net266),
    .A1(_0760_),
    .S(_2217_),
    .X(_2224_));
 sky130_fd_sc_hd__clkbuf_1 _4689_ (.A(_2224_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _4690_ (.A0(net235),
    .A1(_0763_),
    .S(_2217_),
    .X(_2225_));
 sky130_fd_sc_hd__clkbuf_1 _4691_ (.A(_2225_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _4692_ (.A0(net477),
    .A1(_0762_),
    .S(_2217_),
    .X(_2226_));
 sky130_fd_sc_hd__clkbuf_1 _4693_ (.A(_2226_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _4694_ (.A0(net382),
    .A1(_0761_),
    .S(_2217_),
    .X(_2227_));
 sky130_fd_sc_hd__clkbuf_1 _4695_ (.A(_2227_),
    .X(_0081_));
 sky130_fd_sc_hd__buf_4 _4696_ (.A(_2182_),
    .X(_2228_));
 sky130_fd_sc_hd__mux2_1 _4697_ (.A0(net437),
    .A1(_1038_),
    .S(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__clkbuf_1 _4698_ (.A(_2229_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _4699_ (.A0(net206),
    .A1(_0734_),
    .S(_2228_),
    .X(_2230_));
 sky130_fd_sc_hd__clkbuf_1 _4700_ (.A(_2230_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _4701_ (.A0(net328),
    .A1(_0733_),
    .S(_2228_),
    .X(_2231_));
 sky130_fd_sc_hd__clkbuf_1 _4702_ (.A(_2231_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4703_ (.A0(net332),
    .A1(_0732_),
    .S(_2228_),
    .X(_2232_));
 sky130_fd_sc_hd__clkbuf_1 _4704_ (.A(_2232_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _4705_ (.A0(net574),
    .A1(_0729_),
    .S(_2228_),
    .X(_2233_));
 sky130_fd_sc_hd__clkbuf_1 _4706_ (.A(_2233_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _4707_ (.A0(net494),
    .A1(_0730_),
    .S(_2228_),
    .X(_2234_));
 sky130_fd_sc_hd__clkbuf_1 _4708_ (.A(_2234_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _4709_ (.A0(net227),
    .A1(_1426_),
    .S(_2228_),
    .X(_2235_));
 sky130_fd_sc_hd__clkbuf_1 _4710_ (.A(_2235_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _4711_ (.A0(net595),
    .A1(_0727_),
    .S(_2228_),
    .X(_2236_));
 sky130_fd_sc_hd__clkbuf_1 _4712_ (.A(_2236_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _4713_ (.A0(net284),
    .A1(_0738_),
    .S(_2228_),
    .X(_2237_));
 sky130_fd_sc_hd__clkbuf_1 _4714_ (.A(_2237_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _4715_ (.A0(net605),
    .A1(_0737_),
    .S(_2228_),
    .X(_2238_));
 sky130_fd_sc_hd__clkbuf_1 _4716_ (.A(_2238_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _4717_ (.A0(net377),
    .A1(_1227_),
    .S(_2183_),
    .X(_2239_));
 sky130_fd_sc_hd__clkbuf_1 _4718_ (.A(_2239_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _4719_ (.A0(net252),
    .A1(_0739_),
    .S(_2183_),
    .X(_2240_));
 sky130_fd_sc_hd__clkbuf_1 _4720_ (.A(_2240_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4721_ (.A0(net497),
    .A1(_0743_),
    .S(_2183_),
    .X(_2241_));
 sky130_fd_sc_hd__clkbuf_1 _4722_ (.A(_2241_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4723_ (.A0(net241),
    .A1(_0741_),
    .S(_2183_),
    .X(_2242_));
 sky130_fd_sc_hd__clkbuf_1 _4724_ (.A(_2242_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4725_ (.A0(net425),
    .A1(_0742_),
    .S(_2183_),
    .X(_2243_));
 sky130_fd_sc_hd__clkbuf_1 _4726_ (.A(_2243_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _4727_ (.A0(net360),
    .A1(_1954_),
    .S(_2183_),
    .X(_2244_));
 sky130_fd_sc_hd__clkbuf_1 _4728_ (.A(_2244_),
    .X(_0097_));
 sky130_fd_sc_hd__mux4_1 _4729_ (.A0(\fifo.fifo[4][0] ),
    .A1(\fifo.fifo[5][0] ),
    .A2(\fifo.fifo[6][0] ),
    .A3(\fifo.fifo[7][0] ),
    .S0(_0785_),
    .S1(_0789_),
    .X(_2245_));
 sky130_fd_sc_hd__buf_4 _4730_ (.A(\fifo.rd_ptr[0] ),
    .X(_2246_));
 sky130_fd_sc_hd__clkbuf_8 _4731_ (.A(_0782_),
    .X(_2247_));
 sky130_fd_sc_hd__mux4_1 _4732_ (.A0(\fifo.fifo[0][0] ),
    .A1(\fifo.fifo[1][0] ),
    .A2(\fifo.fifo[2][0] ),
    .A3(\fifo.fifo[3][0] ),
    .S0(_2246_),
    .S1(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__mux2_1 _4733_ (.A0(_2245_),
    .A1(_2248_),
    .S(_0781_),
    .X(_2249_));
 sky130_fd_sc_hd__mux2_1 _4734_ (.A0(net222),
    .A1(_2249_),
    .S(_2180_),
    .X(_2250_));
 sky130_fd_sc_hd__clkbuf_1 _4735_ (.A(_2250_),
    .X(_0098_));
 sky130_fd_sc_hd__mux4_1 _4736_ (.A0(\fifo.fifo[4][1] ),
    .A1(\fifo.fifo[5][1] ),
    .A2(\fifo.fifo[6][1] ),
    .A3(\fifo.fifo[7][1] ),
    .S0(_0785_),
    .S1(_0789_),
    .X(_2251_));
 sky130_fd_sc_hd__mux4_1 _4737_ (.A0(\fifo.fifo[0][1] ),
    .A1(\fifo.fifo[1][1] ),
    .A2(\fifo.fifo[2][1] ),
    .A3(\fifo.fifo[3][1] ),
    .S0(_2246_),
    .S1(_2247_),
    .X(_2252_));
 sky130_fd_sc_hd__mux2_1 _4738_ (.A0(_2251_),
    .A1(_2252_),
    .S(_0781_),
    .X(_2253_));
 sky130_fd_sc_hd__mux2_1 _4739_ (.A0(net420),
    .A1(_2253_),
    .S(_2180_),
    .X(_2254_));
 sky130_fd_sc_hd__clkbuf_1 _4740_ (.A(_2254_),
    .X(_0099_));
 sky130_fd_sc_hd__mux4_1 _4741_ (.A0(\fifo.fifo[4][2] ),
    .A1(\fifo.fifo[5][2] ),
    .A2(\fifo.fifo[6][2] ),
    .A3(\fifo.fifo[7][2] ),
    .S0(_0785_),
    .S1(_0789_),
    .X(_2255_));
 sky130_fd_sc_hd__buf_4 _4742_ (.A(\fifo.rd_ptr[1] ),
    .X(_2256_));
 sky130_fd_sc_hd__mux4_1 _4743_ (.A0(\fifo.fifo[0][2] ),
    .A1(\fifo.fifo[1][2] ),
    .A2(\fifo.fifo[2][2] ),
    .A3(\fifo.fifo[3][2] ),
    .S0(_2246_),
    .S1(_2256_),
    .X(_2257_));
 sky130_fd_sc_hd__mux2_1 _4744_ (.A0(_2255_),
    .A1(_2257_),
    .S(_0781_),
    .X(_2258_));
 sky130_fd_sc_hd__mux2_1 _4745_ (.A0(net682),
    .A1(_2258_),
    .S(_2180_),
    .X(_2259_));
 sky130_fd_sc_hd__clkbuf_1 _4746_ (.A(_2259_),
    .X(_0100_));
 sky130_fd_sc_hd__mux4_1 _4747_ (.A0(\fifo.fifo[4][3] ),
    .A1(\fifo.fifo[5][3] ),
    .A2(\fifo.fifo[6][3] ),
    .A3(\fifo.fifo[7][3] ),
    .S0(_0785_),
    .S1(_0789_),
    .X(_2260_));
 sky130_fd_sc_hd__mux4_1 _4748_ (.A0(\fifo.fifo[0][3] ),
    .A1(\fifo.fifo[1][3] ),
    .A2(\fifo.fifo[2][3] ),
    .A3(\fifo.fifo[3][3] ),
    .S0(_2246_),
    .S1(_2256_),
    .X(_2261_));
 sky130_fd_sc_hd__mux2_1 _4749_ (.A0(_2260_),
    .A1(_2261_),
    .S(_0781_),
    .X(_2262_));
 sky130_fd_sc_hd__mux2_1 _4750_ (.A0(net604),
    .A1(_2262_),
    .S(_2180_),
    .X(_2263_));
 sky130_fd_sc_hd__clkbuf_1 _4751_ (.A(_2263_),
    .X(_0101_));
 sky130_fd_sc_hd__mux4_1 _4752_ (.A0(\fifo.fifo[4][4] ),
    .A1(\fifo.fifo[5][4] ),
    .A2(\fifo.fifo[6][4] ),
    .A3(\fifo.fifo[7][4] ),
    .S0(_0785_),
    .S1(_0789_),
    .X(_2264_));
 sky130_fd_sc_hd__mux4_1 _4753_ (.A0(\fifo.fifo[0][4] ),
    .A1(\fifo.fifo[1][4] ),
    .A2(\fifo.fifo[2][4] ),
    .A3(\fifo.fifo[3][4] ),
    .S0(_2246_),
    .S1(_2256_),
    .X(_2265_));
 sky130_fd_sc_hd__mux2_1 _4754_ (.A0(_2264_),
    .A1(_2265_),
    .S(_0781_),
    .X(_2266_));
 sky130_fd_sc_hd__mux2_1 _4755_ (.A0(net684),
    .A1(_2266_),
    .S(_2180_),
    .X(_2267_));
 sky130_fd_sc_hd__clkbuf_1 _4756_ (.A(_2267_),
    .X(_0102_));
 sky130_fd_sc_hd__mux4_1 _4757_ (.A0(\fifo.fifo[4][5] ),
    .A1(\fifo.fifo[5][5] ),
    .A2(\fifo.fifo[6][5] ),
    .A3(\fifo.fifo[7][5] ),
    .S0(_0785_),
    .S1(_0789_),
    .X(_2268_));
 sky130_fd_sc_hd__mux4_1 _4758_ (.A0(\fifo.fifo[0][5] ),
    .A1(\fifo.fifo[1][5] ),
    .A2(\fifo.fifo[2][5] ),
    .A3(\fifo.fifo[3][5] ),
    .S0(_2246_),
    .S1(_2256_),
    .X(_2269_));
 sky130_fd_sc_hd__mux2_1 _4759_ (.A0(_2268_),
    .A1(_2269_),
    .S(_0781_),
    .X(_2270_));
 sky130_fd_sc_hd__mux2_1 _4760_ (.A0(net542),
    .A1(_2270_),
    .S(_2180_),
    .X(_2271_));
 sky130_fd_sc_hd__clkbuf_1 _4761_ (.A(_2271_),
    .X(_0103_));
 sky130_fd_sc_hd__buf_4 _4762_ (.A(_0784_),
    .X(_2272_));
 sky130_fd_sc_hd__mux4_1 _4763_ (.A0(\fifo.fifo[4][6] ),
    .A1(\fifo.fifo[5][6] ),
    .A2(\fifo.fifo[6][6] ),
    .A3(\fifo.fifo[7][6] ),
    .S0(_2272_),
    .S1(_0789_),
    .X(_2273_));
 sky130_fd_sc_hd__mux4_1 _4764_ (.A0(\fifo.fifo[0][6] ),
    .A1(\fifo.fifo[1][6] ),
    .A2(\fifo.fifo[2][6] ),
    .A3(\fifo.fifo[3][6] ),
    .S0(_2246_),
    .S1(_2256_),
    .X(_2274_));
 sky130_fd_sc_hd__mux2_1 _4765_ (.A0(_2273_),
    .A1(_2274_),
    .S(_0781_),
    .X(_2275_));
 sky130_fd_sc_hd__mux2_1 _4766_ (.A0(net693),
    .A1(_2275_),
    .S(_2180_),
    .X(_2276_));
 sky130_fd_sc_hd__clkbuf_1 _4767_ (.A(_2276_),
    .X(_0104_));
 sky130_fd_sc_hd__mux4_1 _4768_ (.A0(\fifo.fifo[4][7] ),
    .A1(\fifo.fifo[5][7] ),
    .A2(\fifo.fifo[6][7] ),
    .A3(\fifo.fifo[7][7] ),
    .S0(_2272_),
    .S1(_0789_),
    .X(_2277_));
 sky130_fd_sc_hd__mux4_1 _4769_ (.A0(\fifo.fifo[0][7] ),
    .A1(\fifo.fifo[1][7] ),
    .A2(\fifo.fifo[2][7] ),
    .A3(\fifo.fifo[3][7] ),
    .S0(_2246_),
    .S1(_2256_),
    .X(_2278_));
 sky130_fd_sc_hd__mux2_1 _4770_ (.A0(_2277_),
    .A1(_2278_),
    .S(_0781_),
    .X(_2279_));
 sky130_fd_sc_hd__mux2_1 _4771_ (.A0(net661),
    .A1(_2279_),
    .S(_2180_),
    .X(_2280_));
 sky130_fd_sc_hd__clkbuf_1 _4772_ (.A(_2280_),
    .X(_0105_));
 sky130_fd_sc_hd__buf_4 _4773_ (.A(_0782_),
    .X(_2281_));
 sky130_fd_sc_hd__mux4_1 _4774_ (.A0(\fifo.fifo[4][8] ),
    .A1(\fifo.fifo[5][8] ),
    .A2(\fifo.fifo[6][8] ),
    .A3(\fifo.fifo[7][8] ),
    .S0(_2272_),
    .S1(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__mux4_1 _4775_ (.A0(\fifo.fifo[0][8] ),
    .A1(\fifo.fifo[1][8] ),
    .A2(\fifo.fifo[2][8] ),
    .A3(\fifo.fifo[3][8] ),
    .S0(_2246_),
    .S1(_2256_),
    .X(_2283_));
 sky130_fd_sc_hd__buf_4 _4776_ (.A(_0780_),
    .X(_2284_));
 sky130_fd_sc_hd__buf_4 _4777_ (.A(_2284_),
    .X(_2285_));
 sky130_fd_sc_hd__mux2_1 _4778_ (.A0(_2282_),
    .A1(_2283_),
    .S(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__mux2_1 _4779_ (.A0(net502),
    .A1(_2286_),
    .S(_2180_),
    .X(_2287_));
 sky130_fd_sc_hd__clkbuf_1 _4780_ (.A(_2287_),
    .X(_0106_));
 sky130_fd_sc_hd__mux4_1 _4781_ (.A0(\fifo.fifo[4][9] ),
    .A1(\fifo.fifo[5][9] ),
    .A2(\fifo.fifo[6][9] ),
    .A3(\fifo.fifo[7][9] ),
    .S0(_2272_),
    .S1(_2281_),
    .X(_2288_));
 sky130_fd_sc_hd__mux4_1 _4782_ (.A0(\fifo.fifo[0][9] ),
    .A1(\fifo.fifo[1][9] ),
    .A2(\fifo.fifo[2][9] ),
    .A3(\fifo.fifo[3][9] ),
    .S0(_2246_),
    .S1(_2256_),
    .X(_2289_));
 sky130_fd_sc_hd__mux2_1 _4783_ (.A0(_2288_),
    .A1(_2289_),
    .S(_2285_),
    .X(_2290_));
 sky130_fd_sc_hd__clkbuf_4 _4784_ (.A(_2177_),
    .X(_2291_));
 sky130_fd_sc_hd__mux2_1 _4785_ (.A0(net675),
    .A1(_2290_),
    .S(_2291_),
    .X(_2292_));
 sky130_fd_sc_hd__clkbuf_1 _4786_ (.A(_2292_),
    .X(_0107_));
 sky130_fd_sc_hd__mux4_1 _4787_ (.A0(\fifo.fifo[4][10] ),
    .A1(\fifo.fifo[5][10] ),
    .A2(\fifo.fifo[6][10] ),
    .A3(\fifo.fifo[7][10] ),
    .S0(_2272_),
    .S1(_2281_),
    .X(_2293_));
 sky130_fd_sc_hd__buf_4 _4788_ (.A(\fifo.rd_ptr[0] ),
    .X(_2294_));
 sky130_fd_sc_hd__mux4_1 _4789_ (.A0(\fifo.fifo[0][10] ),
    .A1(\fifo.fifo[1][10] ),
    .A2(\fifo.fifo[2][10] ),
    .A3(\fifo.fifo[3][10] ),
    .S0(_2294_),
    .S1(_2256_),
    .X(_2295_));
 sky130_fd_sc_hd__mux2_1 _4790_ (.A0(_2293_),
    .A1(_2295_),
    .S(_2285_),
    .X(_2296_));
 sky130_fd_sc_hd__mux2_1 _4791_ (.A0(net696),
    .A1(_2296_),
    .S(_2291_),
    .X(_2297_));
 sky130_fd_sc_hd__clkbuf_1 _4792_ (.A(_2297_),
    .X(_0108_));
 sky130_fd_sc_hd__mux4_1 _4793_ (.A0(\fifo.fifo[4][11] ),
    .A1(\fifo.fifo[5][11] ),
    .A2(\fifo.fifo[6][11] ),
    .A3(\fifo.fifo[7][11] ),
    .S0(_2272_),
    .S1(_2281_),
    .X(_2298_));
 sky130_fd_sc_hd__mux4_1 _4794_ (.A0(\fifo.fifo[0][11] ),
    .A1(\fifo.fifo[1][11] ),
    .A2(\fifo.fifo[2][11] ),
    .A3(\fifo.fifo[3][11] ),
    .S0(_2294_),
    .S1(_2256_),
    .X(_2299_));
 sky130_fd_sc_hd__mux2_1 _4795_ (.A0(_2298_),
    .A1(_2299_),
    .S(_2285_),
    .X(_2300_));
 sky130_fd_sc_hd__mux2_1 _4796_ (.A0(net681),
    .A1(_2300_),
    .S(_2291_),
    .X(_2301_));
 sky130_fd_sc_hd__clkbuf_1 _4797_ (.A(_2301_),
    .X(_0109_));
 sky130_fd_sc_hd__mux4_1 _4798_ (.A0(\fifo.fifo[4][12] ),
    .A1(\fifo.fifo[5][12] ),
    .A2(\fifo.fifo[6][12] ),
    .A3(\fifo.fifo[7][12] ),
    .S0(_2272_),
    .S1(_2281_),
    .X(_2302_));
 sky130_fd_sc_hd__clkbuf_4 _4799_ (.A(\fifo.rd_ptr[1] ),
    .X(_2303_));
 sky130_fd_sc_hd__mux4_1 _4800_ (.A0(\fifo.fifo[0][12] ),
    .A1(\fifo.fifo[1][12] ),
    .A2(\fifo.fifo[2][12] ),
    .A3(\fifo.fifo[3][12] ),
    .S0(_2294_),
    .S1(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__mux2_1 _4801_ (.A0(_2302_),
    .A1(_2304_),
    .S(_2285_),
    .X(_2305_));
 sky130_fd_sc_hd__mux2_1 _4802_ (.A0(net207),
    .A1(_2305_),
    .S(_2291_),
    .X(_2306_));
 sky130_fd_sc_hd__clkbuf_1 _4803_ (.A(_2306_),
    .X(_0110_));
 sky130_fd_sc_hd__mux4_1 _4804_ (.A0(\fifo.fifo[4][13] ),
    .A1(\fifo.fifo[5][13] ),
    .A2(\fifo.fifo[6][13] ),
    .A3(\fifo.fifo[7][13] ),
    .S0(_2272_),
    .S1(_2281_),
    .X(_2307_));
 sky130_fd_sc_hd__mux4_1 _4805_ (.A0(\fifo.fifo[0][13] ),
    .A1(\fifo.fifo[1][13] ),
    .A2(\fifo.fifo[2][13] ),
    .A3(\fifo.fifo[3][13] ),
    .S0(_2294_),
    .S1(_2303_),
    .X(_2308_));
 sky130_fd_sc_hd__mux2_1 _4806_ (.A0(_2307_),
    .A1(_2308_),
    .S(_2285_),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_1 _4807_ (.A0(net488),
    .A1(_2309_),
    .S(_2291_),
    .X(_2310_));
 sky130_fd_sc_hd__clkbuf_1 _4808_ (.A(_2310_),
    .X(_0111_));
 sky130_fd_sc_hd__mux4_1 _4809_ (.A0(\fifo.fifo[4][14] ),
    .A1(\fifo.fifo[5][14] ),
    .A2(\fifo.fifo[6][14] ),
    .A3(\fifo.fifo[7][14] ),
    .S0(_2272_),
    .S1(_2281_),
    .X(_2311_));
 sky130_fd_sc_hd__mux4_1 _4810_ (.A0(\fifo.fifo[0][14] ),
    .A1(\fifo.fifo[1][14] ),
    .A2(\fifo.fifo[2][14] ),
    .A3(\fifo.fifo[3][14] ),
    .S0(_2294_),
    .S1(_2303_),
    .X(_2312_));
 sky130_fd_sc_hd__mux2_1 _4811_ (.A0(_2311_),
    .A1(_2312_),
    .S(_2285_),
    .X(_2313_));
 sky130_fd_sc_hd__mux2_1 _4812_ (.A0(net433),
    .A1(_2313_),
    .S(_2291_),
    .X(_2314_));
 sky130_fd_sc_hd__clkbuf_1 _4813_ (.A(_2314_),
    .X(_0112_));
 sky130_fd_sc_hd__mux4_1 _4814_ (.A0(\fifo.fifo[4][15] ),
    .A1(\fifo.fifo[5][15] ),
    .A2(\fifo.fifo[6][15] ),
    .A3(\fifo.fifo[7][15] ),
    .S0(_2272_),
    .S1(_2281_),
    .X(_2315_));
 sky130_fd_sc_hd__mux4_1 _4815_ (.A0(\fifo.fifo[0][15] ),
    .A1(\fifo.fifo[1][15] ),
    .A2(\fifo.fifo[2][15] ),
    .A3(\fifo.fifo[3][15] ),
    .S0(_2294_),
    .S1(_2303_),
    .X(_2316_));
 sky130_fd_sc_hd__mux2_1 _4816_ (.A0(_2315_),
    .A1(_2316_),
    .S(_2285_),
    .X(_2317_));
 sky130_fd_sc_hd__mux2_1 _4817_ (.A0(net561),
    .A1(_2317_),
    .S(_2291_),
    .X(_2318_));
 sky130_fd_sc_hd__clkbuf_1 _4818_ (.A(_2318_),
    .X(_0113_));
 sky130_fd_sc_hd__buf_4 _4819_ (.A(_0784_),
    .X(_2319_));
 sky130_fd_sc_hd__mux4_1 _4820_ (.A0(\fifo.fifo[4][16] ),
    .A1(\fifo.fifo[5][16] ),
    .A2(\fifo.fifo[6][16] ),
    .A3(\fifo.fifo[7][16] ),
    .S0(_2319_),
    .S1(_2281_),
    .X(_2320_));
 sky130_fd_sc_hd__mux4_1 _4821_ (.A0(\fifo.fifo[0][16] ),
    .A1(\fifo.fifo[1][16] ),
    .A2(\fifo.fifo[2][16] ),
    .A3(\fifo.fifo[3][16] ),
    .S0(_2294_),
    .S1(_2303_),
    .X(_2321_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(_2320_),
    .A1(_2321_),
    .S(_2285_),
    .X(_2322_));
 sky130_fd_sc_hd__mux2_1 _4823_ (.A0(net381),
    .A1(_2322_),
    .S(_2291_),
    .X(_2323_));
 sky130_fd_sc_hd__clkbuf_1 _4824_ (.A(_2323_),
    .X(_0114_));
 sky130_fd_sc_hd__mux4_1 _4825_ (.A0(\fifo.fifo[4][17] ),
    .A1(\fifo.fifo[5][17] ),
    .A2(\fifo.fifo[6][17] ),
    .A3(\fifo.fifo[7][17] ),
    .S0(_2319_),
    .S1(_2281_),
    .X(_2324_));
 sky130_fd_sc_hd__mux4_1 _4826_ (.A0(\fifo.fifo[0][17] ),
    .A1(\fifo.fifo[1][17] ),
    .A2(\fifo.fifo[2][17] ),
    .A3(\fifo.fifo[3][17] ),
    .S0(_2294_),
    .S1(_2303_),
    .X(_2325_));
 sky130_fd_sc_hd__mux2_1 _4827_ (.A0(_2324_),
    .A1(_2325_),
    .S(_2285_),
    .X(_2326_));
 sky130_fd_sc_hd__mux2_1 _4828_ (.A0(net405),
    .A1(_2326_),
    .S(_2291_),
    .X(_2327_));
 sky130_fd_sc_hd__clkbuf_1 _4829_ (.A(_2327_),
    .X(_0115_));
 sky130_fd_sc_hd__buf_4 _4830_ (.A(_0782_),
    .X(_2328_));
 sky130_fd_sc_hd__mux4_1 _4831_ (.A0(\fifo.fifo[4][18] ),
    .A1(\fifo.fifo[5][18] ),
    .A2(\fifo.fifo[6][18] ),
    .A3(\fifo.fifo[7][18] ),
    .S0(_2319_),
    .S1(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__mux4_1 _4832_ (.A0(\fifo.fifo[0][18] ),
    .A1(\fifo.fifo[1][18] ),
    .A2(\fifo.fifo[2][18] ),
    .A3(\fifo.fifo[3][18] ),
    .S0(_2294_),
    .S1(_2303_),
    .X(_2330_));
 sky130_fd_sc_hd__buf_4 _4833_ (.A(_2284_),
    .X(_2331_));
 sky130_fd_sc_hd__mux2_1 _4834_ (.A0(_2329_),
    .A1(_2330_),
    .S(_2331_),
    .X(_2332_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(net218),
    .A1(_2332_),
    .S(_2291_),
    .X(_2333_));
 sky130_fd_sc_hd__clkbuf_1 _4836_ (.A(_2333_),
    .X(_0116_));
 sky130_fd_sc_hd__mux4_1 _4837_ (.A0(\fifo.fifo[4][19] ),
    .A1(\fifo.fifo[5][19] ),
    .A2(\fifo.fifo[6][19] ),
    .A3(\fifo.fifo[7][19] ),
    .S0(_2319_),
    .S1(_2328_),
    .X(_2334_));
 sky130_fd_sc_hd__mux4_1 _4838_ (.A0(\fifo.fifo[0][19] ),
    .A1(\fifo.fifo[1][19] ),
    .A2(\fifo.fifo[2][19] ),
    .A3(\fifo.fifo[3][19] ),
    .S0(_2294_),
    .S1(_2303_),
    .X(_2335_));
 sky130_fd_sc_hd__mux2_1 _4839_ (.A0(_2334_),
    .A1(_2335_),
    .S(_2331_),
    .X(_2336_));
 sky130_fd_sc_hd__clkbuf_4 _4840_ (.A(_2177_),
    .X(_2337_));
 sky130_fd_sc_hd__mux2_1 _4841_ (.A0(net192),
    .A1(_2336_),
    .S(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__clkbuf_1 _4842_ (.A(_2338_),
    .X(_0117_));
 sky130_fd_sc_hd__mux4_1 _4843_ (.A0(\fifo.fifo[4][20] ),
    .A1(\fifo.fifo[5][20] ),
    .A2(\fifo.fifo[6][20] ),
    .A3(\fifo.fifo[7][20] ),
    .S0(_2319_),
    .S1(_2328_),
    .X(_2339_));
 sky130_fd_sc_hd__buf_4 _4844_ (.A(\fifo.rd_ptr[0] ),
    .X(_2340_));
 sky130_fd_sc_hd__mux4_1 _4845_ (.A0(\fifo.fifo[0][20] ),
    .A1(\fifo.fifo[1][20] ),
    .A2(\fifo.fifo[2][20] ),
    .A3(\fifo.fifo[3][20] ),
    .S0(_2340_),
    .S1(_2303_),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _4846_ (.A0(_2339_),
    .A1(_2341_),
    .S(_2331_),
    .X(_2342_));
 sky130_fd_sc_hd__mux2_1 _4847_ (.A0(net698),
    .A1(_2342_),
    .S(_2337_),
    .X(_2343_));
 sky130_fd_sc_hd__clkbuf_1 _4848_ (.A(_2343_),
    .X(_0118_));
 sky130_fd_sc_hd__mux4_1 _4849_ (.A0(\fifo.fifo[4][21] ),
    .A1(\fifo.fifo[5][21] ),
    .A2(\fifo.fifo[6][21] ),
    .A3(\fifo.fifo[7][21] ),
    .S0(_2319_),
    .S1(_2328_),
    .X(_2344_));
 sky130_fd_sc_hd__mux4_1 _4850_ (.A0(\fifo.fifo[0][21] ),
    .A1(\fifo.fifo[1][21] ),
    .A2(\fifo.fifo[2][21] ),
    .A3(\fifo.fifo[3][21] ),
    .S0(_2340_),
    .S1(_2303_),
    .X(_2345_));
 sky130_fd_sc_hd__mux2_1 _4851_ (.A0(_2344_),
    .A1(_2345_),
    .S(_2331_),
    .X(_2346_));
 sky130_fd_sc_hd__mux2_1 _4852_ (.A0(net662),
    .A1(_2346_),
    .S(_2337_),
    .X(_2347_));
 sky130_fd_sc_hd__clkbuf_1 _4853_ (.A(_2347_),
    .X(_0119_));
 sky130_fd_sc_hd__mux4_1 _4854_ (.A0(\fifo.fifo[4][22] ),
    .A1(\fifo.fifo[5][22] ),
    .A2(\fifo.fifo[6][22] ),
    .A3(\fifo.fifo[7][22] ),
    .S0(_2319_),
    .S1(_2328_),
    .X(_2348_));
 sky130_fd_sc_hd__clkbuf_4 _4855_ (.A(\fifo.rd_ptr[1] ),
    .X(_2349_));
 sky130_fd_sc_hd__mux4_1 _4856_ (.A0(\fifo.fifo[0][22] ),
    .A1(\fifo.fifo[1][22] ),
    .A2(\fifo.fifo[2][22] ),
    .A3(\fifo.fifo[3][22] ),
    .S0(_2340_),
    .S1(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__mux2_1 _4857_ (.A0(_2348_),
    .A1(_2350_),
    .S(_2331_),
    .X(_2351_));
 sky130_fd_sc_hd__mux2_1 _4858_ (.A0(net666),
    .A1(_2351_),
    .S(_2337_),
    .X(_2352_));
 sky130_fd_sc_hd__clkbuf_1 _4859_ (.A(_2352_),
    .X(_0120_));
 sky130_fd_sc_hd__mux4_1 _4860_ (.A0(\fifo.fifo[4][23] ),
    .A1(\fifo.fifo[5][23] ),
    .A2(\fifo.fifo[6][23] ),
    .A3(\fifo.fifo[7][23] ),
    .S0(_2319_),
    .S1(_2328_),
    .X(_2353_));
 sky130_fd_sc_hd__mux4_1 _4861_ (.A0(\fifo.fifo[0][23] ),
    .A1(\fifo.fifo[1][23] ),
    .A2(\fifo.fifo[2][23] ),
    .A3(\fifo.fifo[3][23] ),
    .S0(_2340_),
    .S1(_2349_),
    .X(_2354_));
 sky130_fd_sc_hd__mux2_1 _4862_ (.A0(_2353_),
    .A1(_2354_),
    .S(_2331_),
    .X(_2355_));
 sky130_fd_sc_hd__mux2_1 _4863_ (.A0(net722),
    .A1(_2355_),
    .S(_2337_),
    .X(_2356_));
 sky130_fd_sc_hd__clkbuf_1 _4864_ (.A(_2356_),
    .X(_0121_));
 sky130_fd_sc_hd__mux4_1 _4865_ (.A0(\fifo.fifo[4][24] ),
    .A1(\fifo.fifo[5][24] ),
    .A2(\fifo.fifo[6][24] ),
    .A3(\fifo.fifo[7][24] ),
    .S0(_2319_),
    .S1(_2328_),
    .X(_2357_));
 sky130_fd_sc_hd__mux4_1 _4866_ (.A0(\fifo.fifo[0][24] ),
    .A1(\fifo.fifo[1][24] ),
    .A2(\fifo.fifo[2][24] ),
    .A3(\fifo.fifo[3][24] ),
    .S0(_2340_),
    .S1(_2349_),
    .X(_2358_));
 sky130_fd_sc_hd__mux2_1 _4867_ (.A0(_2357_),
    .A1(_2358_),
    .S(_2331_),
    .X(_2359_));
 sky130_fd_sc_hd__mux2_1 _4868_ (.A0(net732),
    .A1(_2359_),
    .S(_2337_),
    .X(_2360_));
 sky130_fd_sc_hd__clkbuf_1 _4869_ (.A(_2360_),
    .X(_0122_));
 sky130_fd_sc_hd__mux4_1 _4870_ (.A0(\fifo.fifo[4][25] ),
    .A1(\fifo.fifo[5][25] ),
    .A2(\fifo.fifo[6][25] ),
    .A3(\fifo.fifo[7][25] ),
    .S0(_2319_),
    .S1(_2328_),
    .X(_2361_));
 sky130_fd_sc_hd__mux4_1 _4871_ (.A0(\fifo.fifo[0][25] ),
    .A1(\fifo.fifo[1][25] ),
    .A2(\fifo.fifo[2][25] ),
    .A3(\fifo.fifo[3][25] ),
    .S0(_2340_),
    .S1(_2349_),
    .X(_2362_));
 sky130_fd_sc_hd__mux2_1 _4872_ (.A0(_2361_),
    .A1(_2362_),
    .S(_2331_),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_1 _4873_ (.A0(net712),
    .A1(_2363_),
    .S(_2337_),
    .X(_2364_));
 sky130_fd_sc_hd__clkbuf_1 _4874_ (.A(_2364_),
    .X(_0123_));
 sky130_fd_sc_hd__buf_4 _4875_ (.A(_0784_),
    .X(_2365_));
 sky130_fd_sc_hd__mux4_1 _4876_ (.A0(\fifo.fifo[4][26] ),
    .A1(\fifo.fifo[5][26] ),
    .A2(\fifo.fifo[6][26] ),
    .A3(\fifo.fifo[7][26] ),
    .S0(_2365_),
    .S1(_2328_),
    .X(_2366_));
 sky130_fd_sc_hd__mux4_1 _4877_ (.A0(\fifo.fifo[0][26] ),
    .A1(\fifo.fifo[1][26] ),
    .A2(\fifo.fifo[2][26] ),
    .A3(\fifo.fifo[3][26] ),
    .S0(_2340_),
    .S1(_2349_),
    .X(_2367_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(_2366_),
    .A1(_2367_),
    .S(_2331_),
    .X(_2368_));
 sky130_fd_sc_hd__mux2_1 _4879_ (.A0(net194),
    .A1(_2368_),
    .S(_2337_),
    .X(_2369_));
 sky130_fd_sc_hd__clkbuf_1 _4880_ (.A(_2369_),
    .X(_0124_));
 sky130_fd_sc_hd__mux4_1 _4881_ (.A0(\fifo.fifo[4][27] ),
    .A1(\fifo.fifo[5][27] ),
    .A2(\fifo.fifo[6][27] ),
    .A3(\fifo.fifo[7][27] ),
    .S0(_2365_),
    .S1(_2328_),
    .X(_2370_));
 sky130_fd_sc_hd__mux4_1 _4882_ (.A0(\fifo.fifo[0][27] ),
    .A1(\fifo.fifo[1][27] ),
    .A2(\fifo.fifo[2][27] ),
    .A3(\fifo.fifo[3][27] ),
    .S0(_2340_),
    .S1(_2349_),
    .X(_2371_));
 sky130_fd_sc_hd__mux2_1 _4883_ (.A0(_2370_),
    .A1(_2371_),
    .S(_2331_),
    .X(_2372_));
 sky130_fd_sc_hd__mux2_1 _4884_ (.A0(net279),
    .A1(_2372_),
    .S(_2337_),
    .X(_2373_));
 sky130_fd_sc_hd__clkbuf_1 _4885_ (.A(_2373_),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_4 _4886_ (.A(_0782_),
    .X(_2374_));
 sky130_fd_sc_hd__mux4_1 _4887_ (.A0(\fifo.fifo[4][28] ),
    .A1(\fifo.fifo[5][28] ),
    .A2(\fifo.fifo[6][28] ),
    .A3(\fifo.fifo[7][28] ),
    .S0(_2365_),
    .S1(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__mux4_1 _4888_ (.A0(\fifo.fifo[0][28] ),
    .A1(\fifo.fifo[1][28] ),
    .A2(\fifo.fifo[2][28] ),
    .A3(\fifo.fifo[3][28] ),
    .S0(_2340_),
    .S1(_2349_),
    .X(_2376_));
 sky130_fd_sc_hd__buf_4 _4889_ (.A(_0780_),
    .X(_2377_));
 sky130_fd_sc_hd__mux2_1 _4890_ (.A0(_2375_),
    .A1(_2376_),
    .S(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__mux2_1 _4891_ (.A0(net672),
    .A1(_2378_),
    .S(_2337_),
    .X(_2379_));
 sky130_fd_sc_hd__clkbuf_1 _4892_ (.A(_2379_),
    .X(_0126_));
 sky130_fd_sc_hd__mux4_1 _4893_ (.A0(\fifo.fifo[4][29] ),
    .A1(\fifo.fifo[5][29] ),
    .A2(\fifo.fifo[6][29] ),
    .A3(\fifo.fifo[7][29] ),
    .S0(_2365_),
    .S1(_2374_),
    .X(_2380_));
 sky130_fd_sc_hd__mux4_1 _4894_ (.A0(\fifo.fifo[0][29] ),
    .A1(\fifo.fifo[1][29] ),
    .A2(\fifo.fifo[2][29] ),
    .A3(\fifo.fifo[3][29] ),
    .S0(_2340_),
    .S1(_2349_),
    .X(_2381_));
 sky130_fd_sc_hd__mux2_1 _4895_ (.A0(_2380_),
    .A1(_2381_),
    .S(_2377_),
    .X(_2382_));
 sky130_fd_sc_hd__buf_4 _4896_ (.A(_2176_),
    .X(_2383_));
 sky130_fd_sc_hd__mux2_1 _4897_ (.A0(\fifo.rd_data[29] ),
    .A1(_2382_),
    .S(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__clkbuf_1 _4898_ (.A(_2384_),
    .X(_0127_));
 sky130_fd_sc_hd__mux4_1 _4899_ (.A0(\fifo.fifo[4][30] ),
    .A1(\fifo.fifo[5][30] ),
    .A2(\fifo.fifo[6][30] ),
    .A3(\fifo.fifo[7][30] ),
    .S0(_2365_),
    .S1(_2374_),
    .X(_2385_));
 sky130_fd_sc_hd__buf_4 _4900_ (.A(\fifo.rd_ptr[0] ),
    .X(_2386_));
 sky130_fd_sc_hd__mux4_1 _4901_ (.A0(\fifo.fifo[0][30] ),
    .A1(\fifo.fifo[1][30] ),
    .A2(\fifo.fifo[2][30] ),
    .A3(\fifo.fifo[3][30] ),
    .S0(_2386_),
    .S1(_2349_),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _4902_ (.A0(_2385_),
    .A1(_2387_),
    .S(_2377_),
    .X(_2388_));
 sky130_fd_sc_hd__mux2_1 _4903_ (.A0(net669),
    .A1(_2388_),
    .S(_2383_),
    .X(_2389_));
 sky130_fd_sc_hd__clkbuf_1 _4904_ (.A(_2389_),
    .X(_0128_));
 sky130_fd_sc_hd__mux4_1 _4905_ (.A0(\fifo.fifo[4][31] ),
    .A1(\fifo.fifo[5][31] ),
    .A2(\fifo.fifo[6][31] ),
    .A3(\fifo.fifo[7][31] ),
    .S0(_2365_),
    .S1(_2374_),
    .X(_2390_));
 sky130_fd_sc_hd__mux4_1 _4906_ (.A0(\fifo.fifo[0][31] ),
    .A1(\fifo.fifo[1][31] ),
    .A2(\fifo.fifo[2][31] ),
    .A3(\fifo.fifo[3][31] ),
    .S0(_2386_),
    .S1(_2349_),
    .X(_2391_));
 sky130_fd_sc_hd__mux2_1 _4907_ (.A0(_2390_),
    .A1(_2391_),
    .S(_2377_),
    .X(_2392_));
 sky130_fd_sc_hd__mux2_1 _4908_ (.A0(net683),
    .A1(_2392_),
    .S(_2383_),
    .X(_2393_));
 sky130_fd_sc_hd__clkbuf_1 _4909_ (.A(_2393_),
    .X(_0129_));
 sky130_fd_sc_hd__mux4_1 _4910_ (.A0(\fifo.fifo[4][32] ),
    .A1(\fifo.fifo[5][32] ),
    .A2(\fifo.fifo[6][32] ),
    .A3(\fifo.fifo[7][32] ),
    .S0(_2365_),
    .S1(_2374_),
    .X(_2394_));
 sky130_fd_sc_hd__buf_4 _4911_ (.A(\fifo.rd_ptr[1] ),
    .X(_2395_));
 sky130_fd_sc_hd__mux4_1 _4912_ (.A0(\fifo.fifo[0][32] ),
    .A1(\fifo.fifo[1][32] ),
    .A2(\fifo.fifo[2][32] ),
    .A3(\fifo.fifo[3][32] ),
    .S0(_2386_),
    .S1(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__mux2_1 _4913_ (.A0(_2394_),
    .A1(_2396_),
    .S(_2377_),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _4914_ (.A0(\fifo.rd_data[32] ),
    .A1(_2397_),
    .S(_2383_),
    .X(_2398_));
 sky130_fd_sc_hd__clkbuf_1 _4915_ (.A(_2398_),
    .X(_0130_));
 sky130_fd_sc_hd__mux4_1 _4916_ (.A0(\fifo.fifo[4][33] ),
    .A1(\fifo.fifo[5][33] ),
    .A2(\fifo.fifo[6][33] ),
    .A3(\fifo.fifo[7][33] ),
    .S0(_2365_),
    .S1(_2374_),
    .X(_2399_));
 sky130_fd_sc_hd__mux4_1 _4917_ (.A0(\fifo.fifo[0][33] ),
    .A1(\fifo.fifo[1][33] ),
    .A2(\fifo.fifo[2][33] ),
    .A3(\fifo.fifo[3][33] ),
    .S0(_2386_),
    .S1(_2395_),
    .X(_2400_));
 sky130_fd_sc_hd__mux2_1 _4918_ (.A0(_2399_),
    .A1(_2400_),
    .S(_2377_),
    .X(_2401_));
 sky130_fd_sc_hd__mux2_1 _4919_ (.A0(net394),
    .A1(_2401_),
    .S(_2383_),
    .X(_2402_));
 sky130_fd_sc_hd__clkbuf_1 _4920_ (.A(_2402_),
    .X(_0131_));
 sky130_fd_sc_hd__mux4_1 _4921_ (.A0(\fifo.fifo[4][34] ),
    .A1(\fifo.fifo[5][34] ),
    .A2(\fifo.fifo[6][34] ),
    .A3(\fifo.fifo[7][34] ),
    .S0(_2365_),
    .S1(_2374_),
    .X(_2403_));
 sky130_fd_sc_hd__mux4_1 _4922_ (.A0(\fifo.fifo[0][34] ),
    .A1(\fifo.fifo[1][34] ),
    .A2(\fifo.fifo[2][34] ),
    .A3(\fifo.fifo[3][34] ),
    .S0(_2386_),
    .S1(_2395_),
    .X(_2404_));
 sky130_fd_sc_hd__mux2_1 _4923_ (.A0(_2403_),
    .A1(_2404_),
    .S(_2377_),
    .X(_2405_));
 sky130_fd_sc_hd__mux2_1 _4924_ (.A0(net202),
    .A1(_2405_),
    .S(_2383_),
    .X(_2406_));
 sky130_fd_sc_hd__clkbuf_1 _4925_ (.A(_2406_),
    .X(_0132_));
 sky130_fd_sc_hd__mux4_1 _4926_ (.A0(\fifo.fifo[4][35] ),
    .A1(\fifo.fifo[5][35] ),
    .A2(\fifo.fifo[6][35] ),
    .A3(\fifo.fifo[7][35] ),
    .S0(_2365_),
    .S1(_2374_),
    .X(_2407_));
 sky130_fd_sc_hd__mux4_1 _4927_ (.A0(\fifo.fifo[0][35] ),
    .A1(\fifo.fifo[1][35] ),
    .A2(\fifo.fifo[2][35] ),
    .A3(\fifo.fifo[3][35] ),
    .S0(_2386_),
    .S1(_2395_),
    .X(_2408_));
 sky130_fd_sc_hd__mux2_1 _4928_ (.A0(_2407_),
    .A1(_2408_),
    .S(_2377_),
    .X(_2409_));
 sky130_fd_sc_hd__mux2_1 _4929_ (.A0(net511),
    .A1(_2409_),
    .S(_2383_),
    .X(_2410_));
 sky130_fd_sc_hd__clkbuf_1 _4930_ (.A(_2410_),
    .X(_0133_));
 sky130_fd_sc_hd__buf_4 _4931_ (.A(\fifo.rd_ptr[0] ),
    .X(_2411_));
 sky130_fd_sc_hd__mux4_1 _4932_ (.A0(\fifo.fifo[4][36] ),
    .A1(\fifo.fifo[5][36] ),
    .A2(\fifo.fifo[6][36] ),
    .A3(\fifo.fifo[7][36] ),
    .S0(_2411_),
    .S1(_2374_),
    .X(_2412_));
 sky130_fd_sc_hd__mux4_1 _4933_ (.A0(\fifo.fifo[0][36] ),
    .A1(\fifo.fifo[1][36] ),
    .A2(\fifo.fifo[2][36] ),
    .A3(\fifo.fifo[3][36] ),
    .S0(_2386_),
    .S1(_2395_),
    .X(_2413_));
 sky130_fd_sc_hd__mux2_1 _4934_ (.A0(_2412_),
    .A1(_2413_),
    .S(_2377_),
    .X(_2414_));
 sky130_fd_sc_hd__mux2_1 _4935_ (.A0(net724),
    .A1(_2414_),
    .S(_2383_),
    .X(_2415_));
 sky130_fd_sc_hd__clkbuf_1 _4936_ (.A(_2415_),
    .X(_0134_));
 sky130_fd_sc_hd__mux4_1 _4937_ (.A0(\fifo.fifo[4][37] ),
    .A1(\fifo.fifo[5][37] ),
    .A2(\fifo.fifo[6][37] ),
    .A3(\fifo.fifo[7][37] ),
    .S0(_2411_),
    .S1(_2374_),
    .X(_2416_));
 sky130_fd_sc_hd__mux4_1 _4938_ (.A0(\fifo.fifo[0][37] ),
    .A1(\fifo.fifo[1][37] ),
    .A2(\fifo.fifo[2][37] ),
    .A3(\fifo.fifo[3][37] ),
    .S0(_2386_),
    .S1(_2395_),
    .X(_2417_));
 sky130_fd_sc_hd__mux2_1 _4939_ (.A0(_2416_),
    .A1(_2417_),
    .S(_2377_),
    .X(_2418_));
 sky130_fd_sc_hd__mux2_1 _4940_ (.A0(net706),
    .A1(_2418_),
    .S(_2383_),
    .X(_2419_));
 sky130_fd_sc_hd__clkbuf_1 _4941_ (.A(_2419_),
    .X(_0135_));
 sky130_fd_sc_hd__buf_4 _4942_ (.A(_0782_),
    .X(_2420_));
 sky130_fd_sc_hd__mux4_1 _4943_ (.A0(\fifo.fifo[4][38] ),
    .A1(\fifo.fifo[5][38] ),
    .A2(\fifo.fifo[6][38] ),
    .A3(\fifo.fifo[7][38] ),
    .S0(_2411_),
    .S1(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__mux4_1 _4944_ (.A0(\fifo.fifo[0][38] ),
    .A1(\fifo.fifo[1][38] ),
    .A2(\fifo.fifo[2][38] ),
    .A3(\fifo.fifo[3][38] ),
    .S0(_2386_),
    .S1(_2395_),
    .X(_2422_));
 sky130_fd_sc_hd__buf_4 _4945_ (.A(_0780_),
    .X(_2423_));
 sky130_fd_sc_hd__mux2_1 _4946_ (.A0(_2421_),
    .A1(_2422_),
    .S(_2423_),
    .X(_2424_));
 sky130_fd_sc_hd__mux2_1 _4947_ (.A0(\fifo.rd_data[38] ),
    .A1(_2424_),
    .S(_2383_),
    .X(_2425_));
 sky130_fd_sc_hd__clkbuf_1 _4948_ (.A(_2425_),
    .X(_0136_));
 sky130_fd_sc_hd__mux4_1 _4949_ (.A0(\fifo.fifo[4][39] ),
    .A1(\fifo.fifo[5][39] ),
    .A2(\fifo.fifo[6][39] ),
    .A3(\fifo.fifo[7][39] ),
    .S0(_2411_),
    .S1(_2420_),
    .X(_2426_));
 sky130_fd_sc_hd__mux4_1 _4950_ (.A0(\fifo.fifo[0][39] ),
    .A1(\fifo.fifo[1][39] ),
    .A2(\fifo.fifo[2][39] ),
    .A3(\fifo.fifo[3][39] ),
    .S0(_2386_),
    .S1(_2395_),
    .X(_2427_));
 sky130_fd_sc_hd__mux2_2 _4951_ (.A0(_2426_),
    .A1(_2427_),
    .S(_2423_),
    .X(_2428_));
 sky130_fd_sc_hd__clkbuf_4 _4952_ (.A(_2176_),
    .X(_2429_));
 sky130_fd_sc_hd__mux2_1 _4953_ (.A0(net733),
    .A1(_2428_),
    .S(_2429_),
    .X(_2430_));
 sky130_fd_sc_hd__clkbuf_1 _4954_ (.A(_2430_),
    .X(_0137_));
 sky130_fd_sc_hd__mux4_1 _4955_ (.A0(\fifo.fifo[4][40] ),
    .A1(\fifo.fifo[5][40] ),
    .A2(\fifo.fifo[6][40] ),
    .A3(\fifo.fifo[7][40] ),
    .S0(_2411_),
    .S1(_2420_),
    .X(_2431_));
 sky130_fd_sc_hd__buf_4 _4956_ (.A(\fifo.rd_ptr[0] ),
    .X(_2432_));
 sky130_fd_sc_hd__mux4_1 _4957_ (.A0(\fifo.fifo[0][40] ),
    .A1(\fifo.fifo[1][40] ),
    .A2(\fifo.fifo[2][40] ),
    .A3(\fifo.fifo[3][40] ),
    .S0(_2432_),
    .S1(_2395_),
    .X(_2433_));
 sky130_fd_sc_hd__mux2_1 _4958_ (.A0(_2431_),
    .A1(_2433_),
    .S(_2423_),
    .X(_2434_));
 sky130_fd_sc_hd__mux2_1 _4959_ (.A0(\fifo.rd_data[40] ),
    .A1(_2434_),
    .S(_2429_),
    .X(_2435_));
 sky130_fd_sc_hd__clkbuf_1 _4960_ (.A(_2435_),
    .X(_0138_));
 sky130_fd_sc_hd__mux4_1 _4961_ (.A0(\fifo.fifo[4][41] ),
    .A1(\fifo.fifo[5][41] ),
    .A2(\fifo.fifo[6][41] ),
    .A3(\fifo.fifo[7][41] ),
    .S0(_2411_),
    .S1(_2420_),
    .X(_2436_));
 sky130_fd_sc_hd__mux4_1 _4962_ (.A0(\fifo.fifo[0][41] ),
    .A1(\fifo.fifo[1][41] ),
    .A2(\fifo.fifo[2][41] ),
    .A3(\fifo.fifo[3][41] ),
    .S0(_2432_),
    .S1(_2395_),
    .X(_2437_));
 sky130_fd_sc_hd__mux2_1 _4963_ (.A0(_2436_),
    .A1(_2437_),
    .S(_2423_),
    .X(_2438_));
 sky130_fd_sc_hd__mux2_1 _4964_ (.A0(net701),
    .A1(_2438_),
    .S(_2429_),
    .X(_2439_));
 sky130_fd_sc_hd__clkbuf_1 _4965_ (.A(_2439_),
    .X(_0139_));
 sky130_fd_sc_hd__mux4_1 _4966_ (.A0(\fifo.fifo[4][42] ),
    .A1(\fifo.fifo[5][42] ),
    .A2(\fifo.fifo[6][42] ),
    .A3(\fifo.fifo[7][42] ),
    .S0(_2411_),
    .S1(_2420_),
    .X(_2440_));
 sky130_fd_sc_hd__clkbuf_4 _4967_ (.A(\fifo.rd_ptr[1] ),
    .X(_2441_));
 sky130_fd_sc_hd__mux4_1 _4968_ (.A0(\fifo.fifo[0][42] ),
    .A1(\fifo.fifo[1][42] ),
    .A2(\fifo.fifo[2][42] ),
    .A3(\fifo.fifo[3][42] ),
    .S0(_2432_),
    .S1(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__mux2_1 _4969_ (.A0(_2440_),
    .A1(_2442_),
    .S(_2423_),
    .X(_2443_));
 sky130_fd_sc_hd__mux2_1 _4970_ (.A0(net499),
    .A1(_2443_),
    .S(_2429_),
    .X(_2444_));
 sky130_fd_sc_hd__clkbuf_1 _4971_ (.A(_2444_),
    .X(_0140_));
 sky130_fd_sc_hd__mux4_1 _4972_ (.A0(\fifo.fifo[4][43] ),
    .A1(\fifo.fifo[5][43] ),
    .A2(\fifo.fifo[6][43] ),
    .A3(\fifo.fifo[7][43] ),
    .S0(_2411_),
    .S1(_2420_),
    .X(_2445_));
 sky130_fd_sc_hd__mux4_1 _4973_ (.A0(\fifo.fifo[0][43] ),
    .A1(\fifo.fifo[1][43] ),
    .A2(\fifo.fifo[2][43] ),
    .A3(\fifo.fifo[3][43] ),
    .S0(_2432_),
    .S1(_2441_),
    .X(_2446_));
 sky130_fd_sc_hd__mux2_1 _4974_ (.A0(_2445_),
    .A1(_2446_),
    .S(_2423_),
    .X(_2447_));
 sky130_fd_sc_hd__mux2_1 _4975_ (.A0(net436),
    .A1(_2447_),
    .S(_2429_),
    .X(_2448_));
 sky130_fd_sc_hd__clkbuf_1 _4976_ (.A(_2448_),
    .X(_0141_));
 sky130_fd_sc_hd__mux4_1 _4977_ (.A0(\fifo.fifo[4][44] ),
    .A1(\fifo.fifo[5][44] ),
    .A2(\fifo.fifo[6][44] ),
    .A3(\fifo.fifo[7][44] ),
    .S0(_2411_),
    .S1(_2420_),
    .X(_2449_));
 sky130_fd_sc_hd__mux4_1 _4978_ (.A0(\fifo.fifo[0][44] ),
    .A1(\fifo.fifo[1][44] ),
    .A2(\fifo.fifo[2][44] ),
    .A3(\fifo.fifo[3][44] ),
    .S0(_2432_),
    .S1(_2441_),
    .X(_2450_));
 sky130_fd_sc_hd__mux2_1 _4979_ (.A0(_2449_),
    .A1(_2450_),
    .S(_2423_),
    .X(_2451_));
 sky130_fd_sc_hd__mux2_1 _4980_ (.A0(net232),
    .A1(_2451_),
    .S(_2429_),
    .X(_2452_));
 sky130_fd_sc_hd__clkbuf_1 _4981_ (.A(_2452_),
    .X(_0142_));
 sky130_fd_sc_hd__mux4_1 _4982_ (.A0(\fifo.fifo[4][45] ),
    .A1(\fifo.fifo[5][45] ),
    .A2(\fifo.fifo[6][45] ),
    .A3(\fifo.fifo[7][45] ),
    .S0(_2411_),
    .S1(_2420_),
    .X(_2453_));
 sky130_fd_sc_hd__mux4_1 _4983_ (.A0(\fifo.fifo[0][45] ),
    .A1(\fifo.fifo[1][45] ),
    .A2(\fifo.fifo[2][45] ),
    .A3(\fifo.fifo[3][45] ),
    .S0(_2432_),
    .S1(_2441_),
    .X(_2454_));
 sky130_fd_sc_hd__mux2_1 _4984_ (.A0(_2453_),
    .A1(_2454_),
    .S(_2423_),
    .X(_2455_));
 sky130_fd_sc_hd__mux2_1 _4985_ (.A0(net422),
    .A1(_2455_),
    .S(_2429_),
    .X(_2456_));
 sky130_fd_sc_hd__clkbuf_1 _4986_ (.A(_2456_),
    .X(_0143_));
 sky130_fd_sc_hd__buf_4 _4987_ (.A(\fifo.rd_ptr[0] ),
    .X(_2457_));
 sky130_fd_sc_hd__mux4_1 _4988_ (.A0(\fifo.fifo[4][46] ),
    .A1(\fifo.fifo[5][46] ),
    .A2(\fifo.fifo[6][46] ),
    .A3(\fifo.fifo[7][46] ),
    .S0(_2457_),
    .S1(_2420_),
    .X(_2458_));
 sky130_fd_sc_hd__mux4_1 _4989_ (.A0(\fifo.fifo[0][46] ),
    .A1(\fifo.fifo[1][46] ),
    .A2(\fifo.fifo[2][46] ),
    .A3(\fifo.fifo[3][46] ),
    .S0(_2432_),
    .S1(_2441_),
    .X(_2459_));
 sky130_fd_sc_hd__mux2_1 _4990_ (.A0(_2458_),
    .A1(_2459_),
    .S(_2423_),
    .X(_2460_));
 sky130_fd_sc_hd__mux2_1 _4991_ (.A0(net231),
    .A1(_2460_),
    .S(_2429_),
    .X(_2461_));
 sky130_fd_sc_hd__clkbuf_1 _4992_ (.A(_2461_),
    .X(_0144_));
 sky130_fd_sc_hd__mux4_1 _4993_ (.A0(\fifo.fifo[4][47] ),
    .A1(\fifo.fifo[5][47] ),
    .A2(\fifo.fifo[6][47] ),
    .A3(\fifo.fifo[7][47] ),
    .S0(_2457_),
    .S1(_2420_),
    .X(_2462_));
 sky130_fd_sc_hd__mux4_1 _4994_ (.A0(\fifo.fifo[0][47] ),
    .A1(\fifo.fifo[1][47] ),
    .A2(\fifo.fifo[2][47] ),
    .A3(\fifo.fifo[3][47] ),
    .S0(_2432_),
    .S1(_2441_),
    .X(_2463_));
 sky130_fd_sc_hd__mux2_1 _4995_ (.A0(_2462_),
    .A1(_2463_),
    .S(_2423_),
    .X(_2464_));
 sky130_fd_sc_hd__mux2_1 _4996_ (.A0(net418),
    .A1(_2464_),
    .S(_2429_),
    .X(_2465_));
 sky130_fd_sc_hd__clkbuf_1 _4997_ (.A(_2465_),
    .X(_0145_));
 sky130_fd_sc_hd__mux4_1 _4998_ (.A0(\fifo.fifo[4][48] ),
    .A1(\fifo.fifo[5][48] ),
    .A2(\fifo.fifo[6][48] ),
    .A3(\fifo.fifo[7][48] ),
    .S0(_2457_),
    .S1(_2247_),
    .X(_2466_));
 sky130_fd_sc_hd__mux4_1 _4999_ (.A0(\fifo.fifo[0][48] ),
    .A1(\fifo.fifo[1][48] ),
    .A2(\fifo.fifo[2][48] ),
    .A3(\fifo.fifo[3][48] ),
    .S0(_2432_),
    .S1(_2441_),
    .X(_2467_));
 sky130_fd_sc_hd__mux2_1 _5000_ (.A0(_2466_),
    .A1(_2467_),
    .S(_2284_),
    .X(_2468_));
 sky130_fd_sc_hd__mux2_1 _5001_ (.A0(net465),
    .A1(_2468_),
    .S(_2429_),
    .X(_2469_));
 sky130_fd_sc_hd__clkbuf_1 _5002_ (.A(_2469_),
    .X(_0146_));
 sky130_fd_sc_hd__mux4_1 _5003_ (.A0(\fifo.fifo[4][49] ),
    .A1(\fifo.fifo[5][49] ),
    .A2(\fifo.fifo[6][49] ),
    .A3(\fifo.fifo[7][49] ),
    .S0(_2457_),
    .S1(_2247_),
    .X(_2470_));
 sky130_fd_sc_hd__mux4_1 _5004_ (.A0(\fifo.fifo[0][49] ),
    .A1(\fifo.fifo[1][49] ),
    .A2(\fifo.fifo[2][49] ),
    .A3(\fifo.fifo[3][49] ),
    .S0(_2432_),
    .S1(_2441_),
    .X(_2471_));
 sky130_fd_sc_hd__mux2_1 _5005_ (.A0(_2470_),
    .A1(_2471_),
    .S(_2284_),
    .X(_2472_));
 sky130_fd_sc_hd__mux2_1 _5006_ (.A0(\fifo.rd_data[49] ),
    .A1(_2472_),
    .S(_2177_),
    .X(_2473_));
 sky130_fd_sc_hd__clkbuf_1 _5007_ (.A(_2473_),
    .X(_0147_));
 sky130_fd_sc_hd__mux4_1 _5008_ (.A0(\fifo.fifo[4][50] ),
    .A1(\fifo.fifo[5][50] ),
    .A2(\fifo.fifo[6][50] ),
    .A3(\fifo.fifo[7][50] ),
    .S0(_2457_),
    .S1(_2247_),
    .X(_2474_));
 sky130_fd_sc_hd__mux4_1 _5009_ (.A0(\fifo.fifo[0][50] ),
    .A1(\fifo.fifo[1][50] ),
    .A2(\fifo.fifo[2][50] ),
    .A3(\fifo.fifo[3][50] ),
    .S0(_0784_),
    .S1(_2441_),
    .X(_2475_));
 sky130_fd_sc_hd__mux2_1 _5010_ (.A0(_2474_),
    .A1(_2475_),
    .S(_2284_),
    .X(_2476_));
 sky130_fd_sc_hd__mux2_1 _5011_ (.A0(\fifo.rd_data[50] ),
    .A1(_2476_),
    .S(_2177_),
    .X(_2477_));
 sky130_fd_sc_hd__clkbuf_1 _5012_ (.A(_2477_),
    .X(_0148_));
 sky130_fd_sc_hd__mux4_1 _5013_ (.A0(\fifo.fifo[4][51] ),
    .A1(\fifo.fifo[5][51] ),
    .A2(\fifo.fifo[6][51] ),
    .A3(\fifo.fifo[7][51] ),
    .S0(_2457_),
    .S1(_2247_),
    .X(_2478_));
 sky130_fd_sc_hd__mux4_1 _5014_ (.A0(\fifo.fifo[0][51] ),
    .A1(\fifo.fifo[1][51] ),
    .A2(\fifo.fifo[2][51] ),
    .A3(\fifo.fifo[3][51] ),
    .S0(_0784_),
    .S1(_2441_),
    .X(_2479_));
 sky130_fd_sc_hd__mux2_1 _5015_ (.A0(_2478_),
    .A1(_2479_),
    .S(_2284_),
    .X(_2480_));
 sky130_fd_sc_hd__mux2_1 _5016_ (.A0(\fifo.rd_data[51] ),
    .A1(_2480_),
    .S(_2177_),
    .X(_2481_));
 sky130_fd_sc_hd__clkbuf_1 _5017_ (.A(_2481_),
    .X(_0149_));
 sky130_fd_sc_hd__mux4_1 _5018_ (.A0(\fifo.fifo[4][52] ),
    .A1(\fifo.fifo[5][52] ),
    .A2(\fifo.fifo[6][52] ),
    .A3(\fifo.fifo[7][52] ),
    .S0(_2457_),
    .S1(_2247_),
    .X(_2482_));
 sky130_fd_sc_hd__mux4_1 _5019_ (.A0(\fifo.fifo[0][52] ),
    .A1(\fifo.fifo[1][52] ),
    .A2(\fifo.fifo[2][52] ),
    .A3(\fifo.fifo[3][52] ),
    .S0(_0784_),
    .S1(_0782_),
    .X(_2483_));
 sky130_fd_sc_hd__mux2_1 _5020_ (.A0(_2482_),
    .A1(_2483_),
    .S(_2284_),
    .X(_2484_));
 sky130_fd_sc_hd__mux2_1 _5021_ (.A0(net346),
    .A1(_2484_),
    .S(_2177_),
    .X(_2485_));
 sky130_fd_sc_hd__clkbuf_1 _5022_ (.A(_2485_),
    .X(_0150_));
 sky130_fd_sc_hd__mux4_1 _5023_ (.A0(\fifo.fifo[4][53] ),
    .A1(\fifo.fifo[5][53] ),
    .A2(\fifo.fifo[6][53] ),
    .A3(\fifo.fifo[7][53] ),
    .S0(_2457_),
    .S1(_2247_),
    .X(_2486_));
 sky130_fd_sc_hd__mux4_1 _5024_ (.A0(\fifo.fifo[0][53] ),
    .A1(\fifo.fifo[1][53] ),
    .A2(\fifo.fifo[2][53] ),
    .A3(\fifo.fifo[3][53] ),
    .S0(_0784_),
    .S1(_0782_),
    .X(_2487_));
 sky130_fd_sc_hd__mux2_1 _5025_ (.A0(_2486_),
    .A1(_2487_),
    .S(_2284_),
    .X(_2488_));
 sky130_fd_sc_hd__mux2_1 _5026_ (.A0(net275),
    .A1(_2488_),
    .S(_2177_),
    .X(_2489_));
 sky130_fd_sc_hd__clkbuf_1 _5027_ (.A(_2489_),
    .X(_0151_));
 sky130_fd_sc_hd__mux4_1 _5028_ (.A0(\fifo.fifo[4][54] ),
    .A1(\fifo.fifo[5][54] ),
    .A2(\fifo.fifo[6][54] ),
    .A3(\fifo.fifo[7][54] ),
    .S0(_2457_),
    .S1(_2247_),
    .X(_2490_));
 sky130_fd_sc_hd__mux4_1 _5029_ (.A0(\fifo.fifo[0][54] ),
    .A1(\fifo.fifo[1][54] ),
    .A2(\fifo.fifo[2][54] ),
    .A3(\fifo.fifo[3][54] ),
    .S0(_0784_),
    .S1(_0782_),
    .X(_2491_));
 sky130_fd_sc_hd__mux2_1 _5030_ (.A0(_2490_),
    .A1(_2491_),
    .S(_2284_),
    .X(_2492_));
 sky130_fd_sc_hd__mux2_1 _5031_ (.A0(net651),
    .A1(_2492_),
    .S(_2177_),
    .X(_2493_));
 sky130_fd_sc_hd__clkbuf_1 _5032_ (.A(_2493_),
    .X(_0152_));
 sky130_fd_sc_hd__mux4_1 _5033_ (.A0(\fifo.fifo[4][55] ),
    .A1(\fifo.fifo[5][55] ),
    .A2(\fifo.fifo[6][55] ),
    .A3(\fifo.fifo[7][55] ),
    .S0(_2457_),
    .S1(_2247_),
    .X(_2494_));
 sky130_fd_sc_hd__mux4_1 _5034_ (.A0(\fifo.fifo[0][55] ),
    .A1(\fifo.fifo[1][55] ),
    .A2(\fifo.fifo[2][55] ),
    .A3(\fifo.fifo[3][55] ),
    .S0(_0784_),
    .S1(_0782_),
    .X(_2495_));
 sky130_fd_sc_hd__mux2_1 _5035_ (.A0(_2494_),
    .A1(_2495_),
    .S(_2284_),
    .X(_2496_));
 sky130_fd_sc_hd__mux2_1 _5036_ (.A0(net668),
    .A1(_2496_),
    .S(_2177_),
    .X(_2497_));
 sky130_fd_sc_hd__clkbuf_1 _5037_ (.A(_2497_),
    .X(_0153_));
 sky130_fd_sc_hd__and3_1 _5038_ (.A(_0772_),
    .B(\fifo.wr_ptr[1] ),
    .C(_0777_),
    .X(_2498_));
 sky130_fd_sc_hd__clkbuf_8 _5039_ (.A(_2498_),
    .X(_2499_));
 sky130_fd_sc_hd__buf_4 _5040_ (.A(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__mux2_1 _5041_ (.A0(net510),
    .A1(_1347_),
    .S(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__clkbuf_1 _5042_ (.A(_2501_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _5043_ (.A0(net513),
    .A1(_0943_),
    .S(_2500_),
    .X(_2502_));
 sky130_fd_sc_hd__clkbuf_1 _5044_ (.A(_2502_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _5045_ (.A0(net555),
    .A1(_0845_),
    .S(_2500_),
    .X(_2503_));
 sky130_fd_sc_hd__clkbuf_1 _5046_ (.A(_2503_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _5047_ (.A0(net212),
    .A1(_0705_),
    .S(_2500_),
    .X(_2504_));
 sky130_fd_sc_hd__clkbuf_1 _5048_ (.A(_2504_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _5049_ (.A0(net343),
    .A1(_0703_),
    .S(_2500_),
    .X(_2505_));
 sky130_fd_sc_hd__clkbuf_1 _5050_ (.A(_2505_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _5051_ (.A0(net535),
    .A1(_0702_),
    .S(_2500_),
    .X(_2506_));
 sky130_fd_sc_hd__clkbuf_1 _5052_ (.A(_2506_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _5053_ (.A0(net466),
    .A1(_1048_),
    .S(_2500_),
    .X(_2507_));
 sky130_fd_sc_hd__clkbuf_1 _5054_ (.A(_2507_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _5055_ (.A0(net655),
    .A1(_0847_),
    .S(_2500_),
    .X(_2508_));
 sky130_fd_sc_hd__clkbuf_1 _5056_ (.A(_2508_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(net568),
    .A1(_0713_),
    .S(_2500_),
    .X(_2509_));
 sky130_fd_sc_hd__clkbuf_1 _5058_ (.A(_2509_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _5059_ (.A0(net330),
    .A1(_0714_),
    .S(_2500_),
    .X(_2510_));
 sky130_fd_sc_hd__clkbuf_1 _5060_ (.A(_2510_),
    .X(_0163_));
 sky130_fd_sc_hd__buf_4 _5061_ (.A(_2499_),
    .X(_2511_));
 sky130_fd_sc_hd__mux2_1 _5062_ (.A0(net618),
    .A1(_1518_),
    .S(_2511_),
    .X(_2512_));
 sky130_fd_sc_hd__clkbuf_1 _5063_ (.A(_2512_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _5064_ (.A0(net355),
    .A1(_0715_),
    .S(_2511_),
    .X(_2513_));
 sky130_fd_sc_hd__clkbuf_1 _5065_ (.A(_2513_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _5066_ (.A0(net417),
    .A1(_0708_),
    .S(_2511_),
    .X(_2514_));
 sky130_fd_sc_hd__clkbuf_1 _5067_ (.A(_2514_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _5068_ (.A0(net627),
    .A1(_0711_),
    .S(_2511_),
    .X(_2515_));
 sky130_fd_sc_hd__clkbuf_1 _5069_ (.A(_2515_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(net599),
    .A1(_0710_),
    .S(_2511_),
    .X(_2516_));
 sky130_fd_sc_hd__clkbuf_1 _5071_ (.A(_2516_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5072_ (.A0(net208),
    .A1(_0709_),
    .S(_2511_),
    .X(_2517_));
 sky130_fd_sc_hd__clkbuf_1 _5073_ (.A(_2517_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _5074_ (.A0(net603),
    .A1(_0880_),
    .S(_2511_),
    .X(_2518_));
 sky130_fd_sc_hd__clkbuf_1 _5075_ (.A(_2518_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5076_ (.A0(net594),
    .A1(_0718_),
    .S(_2511_),
    .X(_2519_));
 sky130_fd_sc_hd__clkbuf_1 _5077_ (.A(_2519_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5078_ (.A0(net373),
    .A1(_1493_),
    .S(_2511_),
    .X(_2520_));
 sky130_fd_sc_hd__clkbuf_1 _5079_ (.A(_2520_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _5080_ (.A0(net524),
    .A1(_0719_),
    .S(_2511_),
    .X(_2521_));
 sky130_fd_sc_hd__clkbuf_1 _5081_ (.A(_2521_),
    .X(_0173_));
 sky130_fd_sc_hd__buf_4 _5082_ (.A(_2499_),
    .X(_2522_));
 sky130_fd_sc_hd__mux2_1 _5083_ (.A0(net276),
    .A1(_0721_),
    .S(_2522_),
    .X(_2523_));
 sky130_fd_sc_hd__clkbuf_1 _5084_ (.A(_2523_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _5085_ (.A0(net583),
    .A1(_0724_),
    .S(_2522_),
    .X(_2524_));
 sky130_fd_sc_hd__clkbuf_1 _5086_ (.A(_2524_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _5087_ (.A0(net345),
    .A1(_0723_),
    .S(_2522_),
    .X(_2525_));
 sky130_fd_sc_hd__clkbuf_1 _5088_ (.A(_2525_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _5089_ (.A0(net573),
    .A1(_0722_),
    .S(_2522_),
    .X(_2526_));
 sky130_fd_sc_hd__clkbuf_1 _5090_ (.A(_2526_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _5091_ (.A0(net237),
    .A1(_0750_),
    .S(_2522_),
    .X(_2527_));
 sky130_fd_sc_hd__clkbuf_1 _5092_ (.A(_2527_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _5093_ (.A0(net610),
    .A1(_0752_),
    .S(_2522_),
    .X(_2528_));
 sky130_fd_sc_hd__clkbuf_1 _5094_ (.A(_2528_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _5095_ (.A0(net640),
    .A1(_0751_),
    .S(_2522_),
    .X(_2529_));
 sky130_fd_sc_hd__clkbuf_1 _5096_ (.A(_2529_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _5097_ (.A0(net409),
    .A1(_1731_),
    .S(_2522_),
    .X(_2530_));
 sky130_fd_sc_hd__clkbuf_1 _5098_ (.A(_2530_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _5099_ (.A0(net427),
    .A1(_0746_),
    .S(_2522_),
    .X(_2531_));
 sky130_fd_sc_hd__clkbuf_1 _5100_ (.A(_2531_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _5101_ (.A0(net475),
    .A1(_0748_),
    .S(_2522_),
    .X(_2532_));
 sky130_fd_sc_hd__clkbuf_1 _5102_ (.A(_2532_),
    .X(_0183_));
 sky130_fd_sc_hd__buf_4 _5103_ (.A(_2499_),
    .X(_2533_));
 sky130_fd_sc_hd__mux2_1 _5104_ (.A0(net223),
    .A1(_0857_),
    .S(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__clkbuf_1 _5105_ (.A(_2534_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _5106_ (.A0(net491),
    .A1(_0747_),
    .S(_2533_),
    .X(_2535_));
 sky130_fd_sc_hd__clkbuf_1 _5107_ (.A(_2535_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _5108_ (.A0(net663),
    .A1(_0755_),
    .S(_2533_),
    .X(_2536_));
 sky130_fd_sc_hd__clkbuf_1 _5109_ (.A(_2536_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _5110_ (.A0(net432),
    .A1(_0756_),
    .S(_2533_),
    .X(_2537_));
 sky130_fd_sc_hd__clkbuf_1 _5111_ (.A(_2537_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _5112_ (.A0(net572),
    .A1(_0757_),
    .S(_2533_),
    .X(_2538_));
 sky130_fd_sc_hd__clkbuf_1 _5113_ (.A(_2538_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _5114_ (.A0(net597),
    .A1(_0758_),
    .S(_2533_),
    .X(_2539_));
 sky130_fd_sc_hd__clkbuf_1 _5115_ (.A(_2539_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _5116_ (.A0(net631),
    .A1(_0760_),
    .S(_2533_),
    .X(_2540_));
 sky130_fd_sc_hd__clkbuf_1 _5117_ (.A(_2540_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _5118_ (.A0(net576),
    .A1(_0763_),
    .S(_2533_),
    .X(_2541_));
 sky130_fd_sc_hd__clkbuf_1 _5119_ (.A(_2541_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _5120_ (.A0(net485),
    .A1(_0762_),
    .S(_2533_),
    .X(_2542_));
 sky130_fd_sc_hd__clkbuf_1 _5121_ (.A(_2542_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _5122_ (.A0(net397),
    .A1(_0761_),
    .S(_2533_),
    .X(_2543_));
 sky130_fd_sc_hd__clkbuf_1 _5123_ (.A(_2543_),
    .X(_0193_));
 sky130_fd_sc_hd__buf_4 _5124_ (.A(_2498_),
    .X(_2544_));
 sky130_fd_sc_hd__mux2_1 _5125_ (.A0(net271),
    .A1(_1038_),
    .S(_2544_),
    .X(_2545_));
 sky130_fd_sc_hd__clkbuf_1 _5126_ (.A(_2545_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _5127_ (.A0(net342),
    .A1(_0734_),
    .S(_2544_),
    .X(_2546_));
 sky130_fd_sc_hd__clkbuf_1 _5128_ (.A(_2546_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(net254),
    .A1(_0733_),
    .S(_2544_),
    .X(_2547_));
 sky130_fd_sc_hd__clkbuf_1 _5130_ (.A(_2547_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _5131_ (.A0(net424),
    .A1(_0732_),
    .S(_2544_),
    .X(_2548_));
 sky130_fd_sc_hd__clkbuf_1 _5132_ (.A(_2548_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _5133_ (.A0(net295),
    .A1(_0729_),
    .S(_2544_),
    .X(_2549_));
 sky130_fd_sc_hd__clkbuf_1 _5134_ (.A(_2549_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _5135_ (.A0(net299),
    .A1(_0730_),
    .S(_2544_),
    .X(_2550_));
 sky130_fd_sc_hd__clkbuf_1 _5136_ (.A(_2550_),
    .X(_0199_));
 sky130_fd_sc_hd__mux2_1 _5137_ (.A0(net221),
    .A1(_1426_),
    .S(_2544_),
    .X(_2551_));
 sky130_fd_sc_hd__clkbuf_1 _5138_ (.A(_2551_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _5139_ (.A0(net451),
    .A1(_0727_),
    .S(_2544_),
    .X(_2552_));
 sky130_fd_sc_hd__clkbuf_1 _5140_ (.A(_2552_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _5141_ (.A0(net196),
    .A1(_0738_),
    .S(_2544_),
    .X(_2553_));
 sky130_fd_sc_hd__clkbuf_1 _5142_ (.A(_2553_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _5143_ (.A0(net359),
    .A1(_0737_),
    .S(_2544_),
    .X(_2554_));
 sky130_fd_sc_hd__clkbuf_1 _5144_ (.A(_2554_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _5145_ (.A0(net304),
    .A1(_1227_),
    .S(_2499_),
    .X(_2555_));
 sky130_fd_sc_hd__clkbuf_1 _5146_ (.A(_2555_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _5147_ (.A0(net305),
    .A1(_0739_),
    .S(_2499_),
    .X(_2556_));
 sky130_fd_sc_hd__clkbuf_1 _5148_ (.A(_2556_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _5149_ (.A0(net248),
    .A1(_0743_),
    .S(_2499_),
    .X(_2557_));
 sky130_fd_sc_hd__clkbuf_1 _5150_ (.A(_2557_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _5151_ (.A0(net622),
    .A1(_0741_),
    .S(_2499_),
    .X(_2558_));
 sky130_fd_sc_hd__clkbuf_1 _5152_ (.A(_2558_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _5153_ (.A0(net636),
    .A1(_0742_),
    .S(_2499_),
    .X(_2559_));
 sky130_fd_sc_hd__clkbuf_1 _5154_ (.A(_2559_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _5155_ (.A0(net441),
    .A1(_1954_),
    .S(_2499_),
    .X(_2560_));
 sky130_fd_sc_hd__clkbuf_1 _5156_ (.A(_2560_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _5157_ (.A0(net205),
    .A1(_1347_),
    .S(_0774_),
    .X(_2561_));
 sky130_fd_sc_hd__clkbuf_1 _5158_ (.A(_2561_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _5159_ (.A0(net632),
    .A1(_0943_),
    .S(_0774_),
    .X(_2562_));
 sky130_fd_sc_hd__clkbuf_1 _5160_ (.A(_2562_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _5161_ (.A0(net211),
    .A1(_0845_),
    .S(_0774_),
    .X(_2563_));
 sky130_fd_sc_hd__clkbuf_1 _5162_ (.A(_2563_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _5163_ (.A0(net516),
    .A1(_0705_),
    .S(_0774_),
    .X(_2564_));
 sky130_fd_sc_hd__clkbuf_1 _5164_ (.A(_2564_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _5165_ (.A0(net486),
    .A1(_0703_),
    .S(_0774_),
    .X(_2565_));
 sky130_fd_sc_hd__clkbuf_1 _5166_ (.A(_2565_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _5167_ (.A0(net559),
    .A1(_0702_),
    .S(_0774_),
    .X(_2566_));
 sky130_fd_sc_hd__clkbuf_1 _5168_ (.A(_2566_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _5169_ (.A0(net395),
    .A1(_1048_),
    .S(_0774_),
    .X(_2567_));
 sky130_fd_sc_hd__clkbuf_1 _5170_ (.A(_2567_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _5171_ (.A0(net473),
    .A1(_0847_),
    .S(_0774_),
    .X(_2568_));
 sky130_fd_sc_hd__clkbuf_1 _5172_ (.A(_2568_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _5173_ (.A0(net249),
    .A1(_0713_),
    .S(_0774_),
    .X(_2569_));
 sky130_fd_sc_hd__clkbuf_1 _5174_ (.A(_2569_),
    .X(_0218_));
 sky130_fd_sc_hd__buf_4 _5175_ (.A(_0773_),
    .X(_2570_));
 sky130_fd_sc_hd__buf_4 _5176_ (.A(_2570_),
    .X(_2571_));
 sky130_fd_sc_hd__mux2_1 _5177_ (.A0(net650),
    .A1(_0714_),
    .S(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__clkbuf_1 _5178_ (.A(_2572_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _5179_ (.A0(net220),
    .A1(_1518_),
    .S(_2571_),
    .X(_2573_));
 sky130_fd_sc_hd__clkbuf_1 _5180_ (.A(_2573_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _5181_ (.A0(net287),
    .A1(_0715_),
    .S(_2571_),
    .X(_2574_));
 sky130_fd_sc_hd__clkbuf_1 _5182_ (.A(_2574_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _5183_ (.A0(net530),
    .A1(_0708_),
    .S(_2571_),
    .X(_2575_));
 sky130_fd_sc_hd__clkbuf_1 _5184_ (.A(_2575_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5185_ (.A0(net567),
    .A1(_0711_),
    .S(_2571_),
    .X(_2576_));
 sky130_fd_sc_hd__clkbuf_1 _5186_ (.A(_2576_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5187_ (.A0(net323),
    .A1(_0710_),
    .S(_2571_),
    .X(_2577_));
 sky130_fd_sc_hd__clkbuf_1 _5188_ (.A(_2577_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _5189_ (.A0(net350),
    .A1(_0709_),
    .S(_2571_),
    .X(_2578_));
 sky130_fd_sc_hd__clkbuf_1 _5190_ (.A(_2578_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _5191_ (.A0(net591),
    .A1(_0880_),
    .S(_2571_),
    .X(_2579_));
 sky130_fd_sc_hd__clkbuf_1 _5192_ (.A(_2579_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _5193_ (.A0(net564),
    .A1(_0718_),
    .S(_2571_),
    .X(_2580_));
 sky130_fd_sc_hd__clkbuf_1 _5194_ (.A(_2580_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _5195_ (.A0(net600),
    .A1(_1493_),
    .S(_2571_),
    .X(_2581_));
 sky130_fd_sc_hd__clkbuf_1 _5196_ (.A(_2581_),
    .X(_0228_));
 sky130_fd_sc_hd__buf_4 _5197_ (.A(_2570_),
    .X(_2582_));
 sky130_fd_sc_hd__mux2_1 _5198_ (.A0(net602),
    .A1(_0719_),
    .S(_2582_),
    .X(_2583_));
 sky130_fd_sc_hd__clkbuf_1 _5199_ (.A(_2583_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _5200_ (.A0(net335),
    .A1(_0721_),
    .S(_2582_),
    .X(_2584_));
 sky130_fd_sc_hd__clkbuf_1 _5201_ (.A(_2584_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _5202_ (.A0(net410),
    .A1(_0724_),
    .S(_2582_),
    .X(_2585_));
 sky130_fd_sc_hd__clkbuf_1 _5203_ (.A(_2585_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _5204_ (.A0(net265),
    .A1(_0723_),
    .S(_2582_),
    .X(_2586_));
 sky130_fd_sc_hd__clkbuf_1 _5205_ (.A(_2586_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _5206_ (.A0(net260),
    .A1(_0722_),
    .S(_2582_),
    .X(_2587_));
 sky130_fd_sc_hd__clkbuf_1 _5207_ (.A(_2587_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _5208_ (.A0(net391),
    .A1(_0750_),
    .S(_2582_),
    .X(_2588_));
 sky130_fd_sc_hd__clkbuf_1 _5209_ (.A(_2588_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _5210_ (.A0(net480),
    .A1(_0752_),
    .S(_2582_),
    .X(_2589_));
 sky130_fd_sc_hd__clkbuf_1 _5211_ (.A(_2589_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _5212_ (.A0(net679),
    .A1(_0751_),
    .S(_2582_),
    .X(_2590_));
 sky130_fd_sc_hd__clkbuf_1 _5213_ (.A(_2590_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _5214_ (.A0(net528),
    .A1(_1731_),
    .S(_2582_),
    .X(_2591_));
 sky130_fd_sc_hd__clkbuf_1 _5215_ (.A(_2591_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _5216_ (.A0(net243),
    .A1(_0746_),
    .S(_2582_),
    .X(_2592_));
 sky130_fd_sc_hd__clkbuf_1 _5217_ (.A(_2592_),
    .X(_0238_));
 sky130_fd_sc_hd__buf_4 _5218_ (.A(_2570_),
    .X(_2593_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(net439),
    .A1(_0748_),
    .S(_2593_),
    .X(_2594_));
 sky130_fd_sc_hd__clkbuf_1 _5220_ (.A(_2594_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _5221_ (.A0(net543),
    .A1(_0857_),
    .S(_2593_),
    .X(_2595_));
 sky130_fd_sc_hd__clkbuf_1 _5222_ (.A(_2595_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5223_ (.A0(net233),
    .A1(_0747_),
    .S(_2593_),
    .X(_2596_));
 sky130_fd_sc_hd__clkbuf_1 _5224_ (.A(_2596_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _5225_ (.A0(net455),
    .A1(_0755_),
    .S(_2593_),
    .X(_2597_));
 sky130_fd_sc_hd__clkbuf_1 _5226_ (.A(_2597_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5227_ (.A0(net216),
    .A1(_0756_),
    .S(_2593_),
    .X(_2598_));
 sky130_fd_sc_hd__clkbuf_1 _5228_ (.A(_2598_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _5229_ (.A0(net230),
    .A1(_0757_),
    .S(_2593_),
    .X(_2599_));
 sky130_fd_sc_hd__clkbuf_1 _5230_ (.A(_2599_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5231_ (.A0(net507),
    .A1(_0758_),
    .S(_2593_),
    .X(_2600_));
 sky130_fd_sc_hd__clkbuf_1 _5232_ (.A(_2600_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5233_ (.A0(net340),
    .A1(_0760_),
    .S(_2593_),
    .X(_2601_));
 sky130_fd_sc_hd__clkbuf_1 _5234_ (.A(_2601_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5235_ (.A0(net274),
    .A1(_0763_),
    .S(_2593_),
    .X(_2602_));
 sky130_fd_sc_hd__clkbuf_1 _5236_ (.A(_2602_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5237_ (.A0(net566),
    .A1(_0762_),
    .S(_2593_),
    .X(_2603_));
 sky130_fd_sc_hd__clkbuf_1 _5238_ (.A(_2603_),
    .X(_0248_));
 sky130_fd_sc_hd__buf_4 _5239_ (.A(_0773_),
    .X(_2604_));
 sky130_fd_sc_hd__mux2_1 _5240_ (.A0(net353),
    .A1(_0761_),
    .S(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__clkbuf_1 _5241_ (.A(_2605_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5242_ (.A0(net435),
    .A1(_1038_),
    .S(_2604_),
    .X(_2606_));
 sky130_fd_sc_hd__clkbuf_1 _5243_ (.A(_2606_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5244_ (.A0(net214),
    .A1(_0734_),
    .S(_2604_),
    .X(_2607_));
 sky130_fd_sc_hd__clkbuf_1 _5245_ (.A(_2607_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5246_ (.A0(net269),
    .A1(_0733_),
    .S(_2604_),
    .X(_2608_));
 sky130_fd_sc_hd__clkbuf_1 _5247_ (.A(_2608_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5248_ (.A0(net283),
    .A1(_0732_),
    .S(_2604_),
    .X(_2609_));
 sky130_fd_sc_hd__clkbuf_1 _5249_ (.A(_2609_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5250_ (.A0(net578),
    .A1(_0729_),
    .S(_2604_),
    .X(_2610_));
 sky130_fd_sc_hd__clkbuf_1 _5251_ (.A(_2610_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5252_ (.A0(net347),
    .A1(_0730_),
    .S(_2604_),
    .X(_2611_));
 sky130_fd_sc_hd__clkbuf_1 _5253_ (.A(_2611_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5254_ (.A0(net238),
    .A1(_1426_),
    .S(_2604_),
    .X(_2612_));
 sky130_fd_sc_hd__clkbuf_1 _5255_ (.A(_2612_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(net376),
    .A1(_0727_),
    .S(_2604_),
    .X(_2613_));
 sky130_fd_sc_hd__clkbuf_1 _5257_ (.A(_2613_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5258_ (.A0(net537),
    .A1(_0738_),
    .S(_2604_),
    .X(_2614_));
 sky130_fd_sc_hd__clkbuf_1 _5259_ (.A(_2614_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5260_ (.A0(net280),
    .A1(_0737_),
    .S(_2570_),
    .X(_2615_));
 sky130_fd_sc_hd__clkbuf_1 _5261_ (.A(_2615_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5262_ (.A0(net367),
    .A1(_1227_),
    .S(_2570_),
    .X(_2616_));
 sky130_fd_sc_hd__clkbuf_1 _5263_ (.A(_2616_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5264_ (.A0(net309),
    .A1(_0739_),
    .S(_2570_),
    .X(_2617_));
 sky130_fd_sc_hd__clkbuf_1 _5265_ (.A(_2617_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5266_ (.A0(net446),
    .A1(_0743_),
    .S(_2570_),
    .X(_2618_));
 sky130_fd_sc_hd__clkbuf_1 _5267_ (.A(_2618_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5268_ (.A0(net215),
    .A1(_0741_),
    .S(_2570_),
    .X(_2619_));
 sky130_fd_sc_hd__clkbuf_1 _5269_ (.A(_2619_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5270_ (.A0(net621),
    .A1(_0742_),
    .S(_2570_),
    .X(_2620_));
 sky130_fd_sc_hd__clkbuf_1 _5271_ (.A(_2620_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5272_ (.A0(net277),
    .A1(_1954_),
    .S(_2570_),
    .X(_2621_));
 sky130_fd_sc_hd__clkbuf_1 _5273_ (.A(_2621_),
    .X(_0265_));
 sky130_fd_sc_hd__and3_1 _5274_ (.A(\fifo.wr_ptr[2] ),
    .B(_0788_),
    .C(_0777_),
    .X(_2622_));
 sky130_fd_sc_hd__clkbuf_8 _5275_ (.A(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__buf_4 _5276_ (.A(_2623_),
    .X(_2624_));
 sky130_fd_sc_hd__mux2_1 _5277_ (.A0(net590),
    .A1(_1347_),
    .S(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__clkbuf_1 _5278_ (.A(_2625_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5279_ (.A0(net302),
    .A1(_0943_),
    .S(_2624_),
    .X(_2626_));
 sky130_fd_sc_hd__clkbuf_1 _5280_ (.A(_2626_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _5281_ (.A0(net372),
    .A1(_0845_),
    .S(_2624_),
    .X(_2627_));
 sky130_fd_sc_hd__clkbuf_1 _5282_ (.A(_2627_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5283_ (.A0(net582),
    .A1(_0705_),
    .S(_2624_),
    .X(_2628_));
 sky130_fd_sc_hd__clkbuf_1 _5284_ (.A(_2628_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5285_ (.A0(net606),
    .A1(_0703_),
    .S(_2624_),
    .X(_2629_));
 sky130_fd_sc_hd__clkbuf_1 _5286_ (.A(_2629_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5287_ (.A0(net312),
    .A1(_0702_),
    .S(_2624_),
    .X(_2630_));
 sky130_fd_sc_hd__clkbuf_1 _5288_ (.A(_2630_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5289_ (.A0(net239),
    .A1(_1048_),
    .S(_2624_),
    .X(_2631_));
 sky130_fd_sc_hd__clkbuf_1 _5290_ (.A(_2631_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5291_ (.A0(net363),
    .A1(_0847_),
    .S(_2624_),
    .X(_2632_));
 sky130_fd_sc_hd__clkbuf_1 _5292_ (.A(_2632_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(net411),
    .A1(_0713_),
    .S(_2624_),
    .X(_2633_));
 sky130_fd_sc_hd__clkbuf_1 _5294_ (.A(_2633_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5295_ (.A0(net365),
    .A1(_0714_),
    .S(_2624_),
    .X(_2634_));
 sky130_fd_sc_hd__clkbuf_1 _5296_ (.A(_2634_),
    .X(_0275_));
 sky130_fd_sc_hd__buf_4 _5297_ (.A(_2623_),
    .X(_2635_));
 sky130_fd_sc_hd__mux2_1 _5298_ (.A0(net317),
    .A1(_1518_),
    .S(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__clkbuf_1 _5299_ (.A(_2636_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(net259),
    .A1(_0715_),
    .S(_2635_),
    .X(_2637_));
 sky130_fd_sc_hd__clkbuf_1 _5301_ (.A(_2637_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5302_ (.A0(net558),
    .A1(_0708_),
    .S(_2635_),
    .X(_2638_));
 sky130_fd_sc_hd__clkbuf_1 _5303_ (.A(_2638_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5304_ (.A0(net400),
    .A1(_0711_),
    .S(_2635_),
    .X(_2639_));
 sky130_fd_sc_hd__clkbuf_1 _5305_ (.A(_2639_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5306_ (.A0(net474),
    .A1(_0710_),
    .S(_2635_),
    .X(_2640_));
 sky130_fd_sc_hd__clkbuf_1 _5307_ (.A(_2640_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _5308_ (.A0(net370),
    .A1(_0709_),
    .S(_2635_),
    .X(_2641_));
 sky130_fd_sc_hd__clkbuf_1 _5309_ (.A(_2641_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _5310_ (.A0(net581),
    .A1(_0880_),
    .S(_2635_),
    .X(_2642_));
 sky130_fd_sc_hd__clkbuf_1 _5311_ (.A(_2642_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _5312_ (.A0(net384),
    .A1(_0718_),
    .S(_2635_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _5313_ (.A(_2643_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _5314_ (.A0(net263),
    .A1(_1493_),
    .S(_2635_),
    .X(_2644_));
 sky130_fd_sc_hd__clkbuf_1 _5315_ (.A(_2644_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _5316_ (.A0(net338),
    .A1(_0719_),
    .S(_2635_),
    .X(_2645_));
 sky130_fd_sc_hd__clkbuf_1 _5317_ (.A(_2645_),
    .X(_0285_));
 sky130_fd_sc_hd__buf_4 _5318_ (.A(_2623_),
    .X(_2646_));
 sky130_fd_sc_hd__mux2_1 _5319_ (.A0(net387),
    .A1(_0721_),
    .S(_2646_),
    .X(_2647_));
 sky130_fd_sc_hd__clkbuf_1 _5320_ (.A(_2647_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _5321_ (.A0(net385),
    .A1(_0724_),
    .S(_2646_),
    .X(_2648_));
 sky130_fd_sc_hd__clkbuf_1 _5322_ (.A(_2648_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _5323_ (.A0(net552),
    .A1(_0723_),
    .S(_2646_),
    .X(_2649_));
 sky130_fd_sc_hd__clkbuf_1 _5324_ (.A(_2649_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _5325_ (.A0(net398),
    .A1(_0722_),
    .S(_2646_),
    .X(_2650_));
 sky130_fd_sc_hd__clkbuf_1 _5326_ (.A(_2650_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _5327_ (.A0(net412),
    .A1(_0750_),
    .S(_2646_),
    .X(_2651_));
 sky130_fd_sc_hd__clkbuf_1 _5328_ (.A(_2651_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _5329_ (.A0(net493),
    .A1(_0752_),
    .S(_2646_),
    .X(_2652_));
 sky130_fd_sc_hd__clkbuf_1 _5330_ (.A(_2652_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _5331_ (.A0(net546),
    .A1(_0751_),
    .S(_2646_),
    .X(_2653_));
 sky130_fd_sc_hd__clkbuf_1 _5332_ (.A(_2653_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _5333_ (.A0(net463),
    .A1(_1731_),
    .S(_2646_),
    .X(_2654_));
 sky130_fd_sc_hd__clkbuf_1 _5334_ (.A(_2654_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _5335_ (.A0(net539),
    .A1(_0746_),
    .S(_2646_),
    .X(_2655_));
 sky130_fd_sc_hd__clkbuf_1 _5336_ (.A(_2655_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _5337_ (.A0(net481),
    .A1(_0748_),
    .S(_2646_),
    .X(_2656_));
 sky130_fd_sc_hd__clkbuf_1 _5338_ (.A(_2656_),
    .X(_0295_));
 sky130_fd_sc_hd__buf_4 _5339_ (.A(_2623_),
    .X(_2657_));
 sky130_fd_sc_hd__mux2_1 _5340_ (.A0(net454),
    .A1(_0857_),
    .S(_2657_),
    .X(_2658_));
 sky130_fd_sc_hd__clkbuf_1 _5341_ (.A(_2658_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _5342_ (.A0(net316),
    .A1(_0747_),
    .S(_2657_),
    .X(_2659_));
 sky130_fd_sc_hd__clkbuf_1 _5343_ (.A(_2659_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _5344_ (.A0(net467),
    .A1(_0755_),
    .S(_2657_),
    .X(_2660_));
 sky130_fd_sc_hd__clkbuf_1 _5345_ (.A(_2660_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(net607),
    .A1(_0756_),
    .S(_2657_),
    .X(_2661_));
 sky130_fd_sc_hd__clkbuf_1 _5347_ (.A(_2661_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _5348_ (.A0(net619),
    .A1(_0757_),
    .S(_2657_),
    .X(_2662_));
 sky130_fd_sc_hd__clkbuf_1 _5349_ (.A(_2662_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(net492),
    .A1(_0758_),
    .S(_2657_),
    .X(_2663_));
 sky130_fd_sc_hd__clkbuf_1 _5351_ (.A(_2663_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _5352_ (.A0(net487),
    .A1(_0760_),
    .S(_2657_),
    .X(_2664_));
 sky130_fd_sc_hd__clkbuf_1 _5353_ (.A(_2664_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _5354_ (.A0(net396),
    .A1(_0763_),
    .S(_2657_),
    .X(_2665_));
 sky130_fd_sc_hd__clkbuf_1 _5355_ (.A(_2665_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _5356_ (.A0(net399),
    .A1(_0762_),
    .S(_2657_),
    .X(_2666_));
 sky130_fd_sc_hd__clkbuf_1 _5357_ (.A(_2666_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _5358_ (.A0(net428),
    .A1(_0761_),
    .S(_2657_),
    .X(_2667_));
 sky130_fd_sc_hd__clkbuf_1 _5359_ (.A(_2667_),
    .X(_0305_));
 sky130_fd_sc_hd__buf_4 _5360_ (.A(_2622_),
    .X(_2668_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(net403),
    .A1(_1038_),
    .S(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__clkbuf_1 _5362_ (.A(_2669_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _5363_ (.A0(net592),
    .A1(_0734_),
    .S(_2668_),
    .X(_2670_));
 sky130_fd_sc_hd__clkbuf_1 _5364_ (.A(_2670_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _5365_ (.A0(net364),
    .A1(_0733_),
    .S(_2668_),
    .X(_2671_));
 sky130_fd_sc_hd__clkbuf_1 _5366_ (.A(_2671_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(net554),
    .A1(_0732_),
    .S(_2668_),
    .X(_2672_));
 sky130_fd_sc_hd__clkbuf_1 _5368_ (.A(_2672_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _5369_ (.A0(net500),
    .A1(_0729_),
    .S(_2668_),
    .X(_2673_));
 sky130_fd_sc_hd__clkbuf_1 _5370_ (.A(_2673_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(net291),
    .A1(_0730_),
    .S(_2668_),
    .X(_2674_));
 sky130_fd_sc_hd__clkbuf_1 _5372_ (.A(_2674_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(net389),
    .A1(_1426_),
    .S(_2668_),
    .X(_2675_));
 sky130_fd_sc_hd__clkbuf_1 _5374_ (.A(_2675_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _5375_ (.A0(net383),
    .A1(_0727_),
    .S(_2668_),
    .X(_2676_));
 sky130_fd_sc_hd__clkbuf_1 _5376_ (.A(_2676_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _5377_ (.A0(net553),
    .A1(_0738_),
    .S(_2668_),
    .X(_2677_));
 sky130_fd_sc_hd__clkbuf_1 _5378_ (.A(_2677_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _5379_ (.A0(net585),
    .A1(_0737_),
    .S(_2668_),
    .X(_2678_));
 sky130_fd_sc_hd__clkbuf_1 _5380_ (.A(_2678_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _5381_ (.A0(net318),
    .A1(_1227_),
    .S(_2623_),
    .X(_2679_));
 sky130_fd_sc_hd__clkbuf_1 _5382_ (.A(_2679_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(net236),
    .A1(_0739_),
    .S(_2623_),
    .X(_2680_));
 sky130_fd_sc_hd__clkbuf_1 _5384_ (.A(_2680_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _5385_ (.A0(net529),
    .A1(_0743_),
    .S(_2623_),
    .X(_2681_));
 sky130_fd_sc_hd__clkbuf_1 _5386_ (.A(_2681_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _5387_ (.A0(net408),
    .A1(_0741_),
    .S(_2623_),
    .X(_2682_));
 sky130_fd_sc_hd__clkbuf_1 _5388_ (.A(_2682_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _5389_ (.A0(net264),
    .A1(_0742_),
    .S(_2623_),
    .X(_2683_));
 sky130_fd_sc_hd__clkbuf_1 _5390_ (.A(_2683_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _5391_ (.A0(net324),
    .A1(_1954_),
    .S(_2623_),
    .X(_2684_));
 sky130_fd_sc_hd__clkbuf_1 _5392_ (.A(_2684_),
    .X(_0321_));
 sky130_fd_sc_hd__and3_1 _5393_ (.A(\fifo.wr_ptr[2] ),
    .B(\fifo.wr_ptr[1] ),
    .C(_0777_),
    .X(_2685_));
 sky130_fd_sc_hd__clkbuf_8 _5394_ (.A(_2685_),
    .X(_2686_));
 sky130_fd_sc_hd__buf_4 _5395_ (.A(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__mux2_1 _5396_ (.A0(net267),
    .A1(_1347_),
    .S(_2687_),
    .X(_2688_));
 sky130_fd_sc_hd__clkbuf_1 _5397_ (.A(_2688_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _5398_ (.A0(net253),
    .A1(_0943_),
    .S(_2687_),
    .X(_2689_));
 sky130_fd_sc_hd__clkbuf_1 _5399_ (.A(_2689_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _5400_ (.A0(net575),
    .A1(_0845_),
    .S(_2687_),
    .X(_2690_));
 sky130_fd_sc_hd__clkbuf_1 _5401_ (.A(_2690_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _5402_ (.A0(net217),
    .A1(_0705_),
    .S(_2687_),
    .X(_2691_));
 sky130_fd_sc_hd__clkbuf_1 _5403_ (.A(_2691_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(net292),
    .A1(_0703_),
    .S(_2687_),
    .X(_2692_));
 sky130_fd_sc_hd__clkbuf_1 _5405_ (.A(_2692_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _5406_ (.A0(net209),
    .A1(_0702_),
    .S(_2687_),
    .X(_2693_));
 sky130_fd_sc_hd__clkbuf_1 _5407_ (.A(_2693_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _5408_ (.A0(net336),
    .A1(_1048_),
    .S(_2687_),
    .X(_2694_));
 sky130_fd_sc_hd__clkbuf_1 _5409_ (.A(_2694_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _5410_ (.A0(net348),
    .A1(_0847_),
    .S(_2687_),
    .X(_2695_));
 sky130_fd_sc_hd__clkbuf_1 _5411_ (.A(_2695_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _5412_ (.A0(net504),
    .A1(_0713_),
    .S(_2687_),
    .X(_2696_));
 sky130_fd_sc_hd__clkbuf_1 _5413_ (.A(_2696_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _5414_ (.A0(net320),
    .A1(_0714_),
    .S(_2687_),
    .X(_2697_));
 sky130_fd_sc_hd__clkbuf_1 _5415_ (.A(_2697_),
    .X(_0331_));
 sky130_fd_sc_hd__buf_4 _5416_ (.A(_2686_),
    .X(_2698_));
 sky130_fd_sc_hd__mux2_1 _5417_ (.A0(net671),
    .A1(_1518_),
    .S(_2698_),
    .X(_2699_));
 sky130_fd_sc_hd__clkbuf_1 _5418_ (.A(_2699_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _5419_ (.A0(net625),
    .A1(_0715_),
    .S(_2698_),
    .X(_2700_));
 sky130_fd_sc_hd__clkbuf_1 _5420_ (.A(_2700_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _5421_ (.A0(net378),
    .A1(_0708_),
    .S(_2698_),
    .X(_2701_));
 sky130_fd_sc_hd__clkbuf_1 _5422_ (.A(_2701_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _5423_ (.A0(net598),
    .A1(_0711_),
    .S(_2698_),
    .X(_2702_));
 sky130_fd_sc_hd__clkbuf_1 _5424_ (.A(_2702_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _5425_ (.A0(net624),
    .A1(_0710_),
    .S(_2698_),
    .X(_2703_));
 sky130_fd_sc_hd__clkbuf_1 _5426_ (.A(_2703_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _5427_ (.A0(net557),
    .A1(_0709_),
    .S(_2698_),
    .X(_2704_));
 sky130_fd_sc_hd__clkbuf_1 _5428_ (.A(_2704_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _5429_ (.A0(net623),
    .A1(_0880_),
    .S(_2698_),
    .X(_2705_));
 sky130_fd_sc_hd__clkbuf_1 _5430_ (.A(_2705_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _5431_ (.A0(net469),
    .A1(_0718_),
    .S(_2698_),
    .X(_2706_));
 sky130_fd_sc_hd__clkbuf_1 _5432_ (.A(_2706_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _5433_ (.A0(net461),
    .A1(_1493_),
    .S(_2698_),
    .X(_2707_));
 sky130_fd_sc_hd__clkbuf_1 _5434_ (.A(_2707_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _5435_ (.A0(net464),
    .A1(_0719_),
    .S(_2698_),
    .X(_2708_));
 sky130_fd_sc_hd__clkbuf_1 _5436_ (.A(_2708_),
    .X(_0341_));
 sky130_fd_sc_hd__buf_4 _5437_ (.A(_2686_),
    .X(_2709_));
 sky130_fd_sc_hd__mux2_1 _5438_ (.A0(net319),
    .A1(_0721_),
    .S(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__clkbuf_1 _5439_ (.A(_2710_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(net645),
    .A1(_0724_),
    .S(_2709_),
    .X(_2711_));
 sky130_fd_sc_hd__clkbuf_1 _5441_ (.A(_2711_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _5442_ (.A0(net298),
    .A1(_0723_),
    .S(_2709_),
    .X(_2712_));
 sky130_fd_sc_hd__clkbuf_1 _5443_ (.A(_2712_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _5444_ (.A0(net550),
    .A1(_0722_),
    .S(_2709_),
    .X(_2713_));
 sky130_fd_sc_hd__clkbuf_1 _5445_ (.A(_2713_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _5446_ (.A0(net514),
    .A1(_0750_),
    .S(_2709_),
    .X(_2714_));
 sky130_fd_sc_hd__clkbuf_1 _5447_ (.A(_2714_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _5448_ (.A0(net656),
    .A1(_0752_),
    .S(_2709_),
    .X(_2715_));
 sky130_fd_sc_hd__clkbuf_1 _5449_ (.A(_2715_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _5450_ (.A0(net680),
    .A1(_0751_),
    .S(_2709_),
    .X(_2716_));
 sky130_fd_sc_hd__clkbuf_1 _5451_ (.A(_2716_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _5452_ (.A0(net589),
    .A1(_1731_),
    .S(_2709_),
    .X(_2717_));
 sky130_fd_sc_hd__clkbuf_1 _5453_ (.A(_2717_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _5454_ (.A0(net565),
    .A1(_0746_),
    .S(_2709_),
    .X(_2718_));
 sky130_fd_sc_hd__clkbuf_1 _5455_ (.A(_2718_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _5456_ (.A0(net458),
    .A1(_0748_),
    .S(_2709_),
    .X(_2719_));
 sky130_fd_sc_hd__clkbuf_1 _5457_ (.A(_2719_),
    .X(_0351_));
 sky130_fd_sc_hd__buf_4 _5458_ (.A(_2686_),
    .X(_2720_));
 sky130_fd_sc_hd__mux2_1 _5459_ (.A0(net643),
    .A1(_0857_),
    .S(_2720_),
    .X(_2721_));
 sky130_fd_sc_hd__clkbuf_1 _5460_ (.A(_2721_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(net526),
    .A1(_0747_),
    .S(_2720_),
    .X(_2722_));
 sky130_fd_sc_hd__clkbuf_1 _5462_ (.A(_2722_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _5463_ (.A0(net406),
    .A1(_0755_),
    .S(_2720_),
    .X(_2723_));
 sky130_fd_sc_hd__clkbuf_1 _5464_ (.A(_2723_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _5465_ (.A0(net649),
    .A1(_0756_),
    .S(_2720_),
    .X(_2724_));
 sky130_fd_sc_hd__clkbuf_1 _5466_ (.A(_2724_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _5467_ (.A0(net596),
    .A1(_0757_),
    .S(_2720_),
    .X(_2725_));
 sky130_fd_sc_hd__clkbuf_1 _5468_ (.A(_2725_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _5469_ (.A0(net371),
    .A1(_0758_),
    .S(_2720_),
    .X(_2726_));
 sky130_fd_sc_hd__clkbuf_1 _5470_ (.A(_2726_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(net459),
    .A1(_0760_),
    .S(_2720_),
    .X(_2727_));
 sky130_fd_sc_hd__clkbuf_1 _5472_ (.A(_2727_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(net556),
    .A1(_0763_),
    .S(_2720_),
    .X(_2728_));
 sky130_fd_sc_hd__clkbuf_1 _5474_ (.A(_2728_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _5475_ (.A0(net691),
    .A1(_0762_),
    .S(_2720_),
    .X(_2729_));
 sky130_fd_sc_hd__clkbuf_1 _5476_ (.A(_2729_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _5477_ (.A0(net615),
    .A1(_0761_),
    .S(_2720_),
    .X(_2730_));
 sky130_fd_sc_hd__clkbuf_1 _5478_ (.A(_2730_),
    .X(_0361_));
 sky130_fd_sc_hd__buf_4 _5479_ (.A(_2685_),
    .X(_2731_));
 sky130_fd_sc_hd__mux2_1 _5480_ (.A0(net522),
    .A1(_1038_),
    .S(_2731_),
    .X(_2732_));
 sky130_fd_sc_hd__clkbuf_1 _5481_ (.A(_2732_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _5482_ (.A0(net219),
    .A1(_0734_),
    .S(_2731_),
    .X(_2733_));
 sky130_fd_sc_hd__clkbuf_1 _5483_ (.A(_2733_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _5484_ (.A0(net251),
    .A1(_0733_),
    .S(_2731_),
    .X(_2734_));
 sky130_fd_sc_hd__clkbuf_1 _5485_ (.A(_2734_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _5486_ (.A0(net407),
    .A1(_0732_),
    .S(_2731_),
    .X(_2735_));
 sky130_fd_sc_hd__clkbuf_1 _5487_ (.A(_2735_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _5488_ (.A0(net368),
    .A1(_0729_),
    .S(_2731_),
    .X(_2736_));
 sky130_fd_sc_hd__clkbuf_1 _5489_ (.A(_2736_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _5490_ (.A0(net329),
    .A1(_0730_),
    .S(_2731_),
    .X(_2737_));
 sky130_fd_sc_hd__clkbuf_1 _5491_ (.A(_2737_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _5492_ (.A0(net285),
    .A1(_1426_),
    .S(_2731_),
    .X(_2738_));
 sky130_fd_sc_hd__clkbuf_1 _5493_ (.A(_2738_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(net245),
    .A1(_0727_),
    .S(_2731_),
    .X(_2739_));
 sky130_fd_sc_hd__clkbuf_1 _5495_ (.A(_2739_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _5496_ (.A0(net438),
    .A1(_0738_),
    .S(_2731_),
    .X(_2740_));
 sky130_fd_sc_hd__clkbuf_1 _5497_ (.A(_2740_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _5498_ (.A0(net531),
    .A1(_0737_),
    .S(_2731_),
    .X(_2741_));
 sky130_fd_sc_hd__clkbuf_1 _5499_ (.A(_2741_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _5500_ (.A0(net213),
    .A1(_1227_),
    .S(_2686_),
    .X(_2742_));
 sky130_fd_sc_hd__clkbuf_1 _5501_ (.A(_2742_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _5502_ (.A0(net536),
    .A1(_0739_),
    .S(_2686_),
    .X(_2743_));
 sky130_fd_sc_hd__clkbuf_1 _5503_ (.A(_2743_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _5504_ (.A0(net545),
    .A1(_0743_),
    .S(_2686_),
    .X(_2744_));
 sky130_fd_sc_hd__clkbuf_1 _5505_ (.A(_2744_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _5506_ (.A0(net532),
    .A1(_0741_),
    .S(_2686_),
    .X(_2745_));
 sky130_fd_sc_hd__clkbuf_1 _5507_ (.A(_2745_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _5508_ (.A0(net326),
    .A1(_0742_),
    .S(_2686_),
    .X(_2746_));
 sky130_fd_sc_hd__clkbuf_1 _5509_ (.A(_2746_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _5510_ (.A0(net635),
    .A1(_1954_),
    .S(_2686_),
    .X(_2747_));
 sky130_fd_sc_hd__clkbuf_1 _5511_ (.A(_2747_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_8 _5512_ (.A(net123),
    .X(_2748_));
 sky130_fd_sc_hd__clkbuf_8 _5513_ (.A(_2748_),
    .X(_2749_));
 sky130_fd_sc_hd__inv_2 _5514_ (.A(_2749_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _5515_ (.A(_2749_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _5516_ (.A(_2749_),
    .Y(_0002_));
 sky130_fd_sc_hd__and3_1 _5517_ (.A(_0772_),
    .B(_0788_),
    .C(_0770_),
    .X(_2750_));
 sky130_fd_sc_hd__clkbuf_8 _5518_ (.A(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__buf_4 _5519_ (.A(_2751_),
    .X(_2752_));
 sky130_fd_sc_hd__mux2_1 _5520_ (.A0(net495),
    .A1(_1347_),
    .S(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__clkbuf_1 _5521_ (.A(_2753_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _5522_ (.A0(net444),
    .A1(_0943_),
    .S(_2752_),
    .X(_2754_));
 sky130_fd_sc_hd__clkbuf_1 _5523_ (.A(_2754_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _5524_ (.A0(net300),
    .A1(_0845_),
    .S(_2752_),
    .X(_2755_));
 sky130_fd_sc_hd__clkbuf_1 _5525_ (.A(_2755_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _5526_ (.A0(net628),
    .A1(_0705_),
    .S(_2752_),
    .X(_2756_));
 sky130_fd_sc_hd__clkbuf_1 _5527_ (.A(_2756_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _5528_ (.A0(net601),
    .A1(_0703_),
    .S(_2752_),
    .X(_2757_));
 sky130_fd_sc_hd__clkbuf_1 _5529_ (.A(_2757_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _5530_ (.A0(net322),
    .A1(_0702_),
    .S(_2752_),
    .X(_2758_));
 sky130_fd_sc_hd__clkbuf_1 _5531_ (.A(_2758_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(net527),
    .A1(_1048_),
    .S(_2752_),
    .X(_2759_));
 sky130_fd_sc_hd__clkbuf_1 _5533_ (.A(_2759_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(net333),
    .A1(_0847_),
    .S(_2752_),
    .X(_2760_));
 sky130_fd_sc_hd__clkbuf_1 _5535_ (.A(_2760_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _5536_ (.A0(net678),
    .A1(_0713_),
    .S(_2752_),
    .X(_2761_));
 sky130_fd_sc_hd__clkbuf_1 _5537_ (.A(_2761_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _5538_ (.A0(net362),
    .A1(_0714_),
    .S(_2752_),
    .X(_2762_));
 sky130_fd_sc_hd__clkbuf_1 _5539_ (.A(_2762_),
    .X(_0390_));
 sky130_fd_sc_hd__buf_4 _5540_ (.A(_2751_),
    .X(_2763_));
 sky130_fd_sc_hd__mux2_1 _5541_ (.A0(net521),
    .A1(_1518_),
    .S(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__clkbuf_1 _5542_ (.A(_2764_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(net199),
    .A1(_0715_),
    .S(_2763_),
    .X(_2765_));
 sky130_fd_sc_hd__clkbuf_1 _5544_ (.A(_2765_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _5545_ (.A0(net270),
    .A1(_0708_),
    .S(_2763_),
    .X(_2766_));
 sky130_fd_sc_hd__clkbuf_1 _5546_ (.A(_2766_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(net247),
    .A1(_0711_),
    .S(_2763_),
    .X(_2767_));
 sky130_fd_sc_hd__clkbuf_1 _5548_ (.A(_2767_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _5549_ (.A0(net321),
    .A1(_0710_),
    .S(_2763_),
    .X(_2768_));
 sky130_fd_sc_hd__clkbuf_1 _5550_ (.A(_2768_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _5551_ (.A0(net393),
    .A1(_0709_),
    .S(_2763_),
    .X(_2769_));
 sky130_fd_sc_hd__clkbuf_1 _5552_ (.A(_2769_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _5553_ (.A0(net273),
    .A1(_0880_),
    .S(_2763_),
    .X(_2770_));
 sky130_fd_sc_hd__clkbuf_1 _5554_ (.A(_2770_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _5555_ (.A0(net440),
    .A1(_0718_),
    .S(_2763_),
    .X(_2771_));
 sky130_fd_sc_hd__clkbuf_1 _5556_ (.A(_2771_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _5557_ (.A0(net246),
    .A1(_1493_),
    .S(_2763_),
    .X(_2772_));
 sky130_fd_sc_hd__clkbuf_1 _5558_ (.A(_2772_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _5559_ (.A0(net289),
    .A1(_0719_),
    .S(_2763_),
    .X(_2773_));
 sky130_fd_sc_hd__clkbuf_1 _5560_ (.A(_2773_),
    .X(_0400_));
 sky130_fd_sc_hd__buf_4 _5561_ (.A(_2751_),
    .X(_2774_));
 sky130_fd_sc_hd__mux2_1 _5562_ (.A0(net515),
    .A1(_0721_),
    .S(_2774_),
    .X(_2775_));
 sky130_fd_sc_hd__clkbuf_1 _5563_ (.A(_2775_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _5564_ (.A0(net352),
    .A1(_0724_),
    .S(_2774_),
    .X(_2776_));
 sky130_fd_sc_hd__clkbuf_1 _5565_ (.A(_2776_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _5566_ (.A0(net534),
    .A1(_0723_),
    .S(_2774_),
    .X(_2777_));
 sky130_fd_sc_hd__clkbuf_1 _5567_ (.A(_2777_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _5568_ (.A0(net296),
    .A1(_0722_),
    .S(_2774_),
    .X(_2778_));
 sky130_fd_sc_hd__clkbuf_1 _5569_ (.A(_2778_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _5570_ (.A0(net646),
    .A1(_0750_),
    .S(_2774_),
    .X(_2779_));
 sky130_fd_sc_hd__clkbuf_1 _5571_ (.A(_2779_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _5572_ (.A0(net386),
    .A1(_0752_),
    .S(_2774_),
    .X(_2780_));
 sky130_fd_sc_hd__clkbuf_1 _5573_ (.A(_2780_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(net225),
    .A1(_0751_),
    .S(_2774_),
    .X(_2781_));
 sky130_fd_sc_hd__clkbuf_1 _5575_ (.A(_2781_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _5576_ (.A0(net195),
    .A1(_1731_),
    .S(_2774_),
    .X(_2782_));
 sky130_fd_sc_hd__clkbuf_1 _5577_ (.A(_2782_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _5578_ (.A0(net431),
    .A1(_0746_),
    .S(_2774_),
    .X(_2783_));
 sky130_fd_sc_hd__clkbuf_1 _5579_ (.A(_2783_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _5580_ (.A0(net268),
    .A1(_0748_),
    .S(_2774_),
    .X(_2784_));
 sky130_fd_sc_hd__clkbuf_1 _5581_ (.A(_2784_),
    .X(_0410_));
 sky130_fd_sc_hd__buf_4 _5582_ (.A(_2751_),
    .X(_2785_));
 sky130_fd_sc_hd__mux2_1 _5583_ (.A0(net327),
    .A1(_0857_),
    .S(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__clkbuf_1 _5584_ (.A(_2786_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _5585_ (.A0(net659),
    .A1(_0747_),
    .S(_2785_),
    .X(_2787_));
 sky130_fd_sc_hd__clkbuf_1 _5586_ (.A(_2787_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _5587_ (.A0(net468),
    .A1(_0755_),
    .S(_2785_),
    .X(_2788_));
 sky130_fd_sc_hd__clkbuf_1 _5588_ (.A(_2788_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _5589_ (.A0(net226),
    .A1(_0756_),
    .S(_2785_),
    .X(_2789_));
 sky130_fd_sc_hd__clkbuf_1 _5590_ (.A(_2789_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _5591_ (.A0(net331),
    .A1(_0757_),
    .S(_2785_),
    .X(_2790_));
 sky130_fd_sc_hd__clkbuf_1 _5592_ (.A(_2790_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _5593_ (.A0(net228),
    .A1(_0758_),
    .S(_2785_),
    .X(_2791_));
 sky130_fd_sc_hd__clkbuf_1 _5594_ (.A(_2791_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _5595_ (.A0(net311),
    .A1(_0760_),
    .S(_2785_),
    .X(_2792_));
 sky130_fd_sc_hd__clkbuf_1 _5596_ (.A(_2792_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(net250),
    .A1(_0763_),
    .S(_2785_),
    .X(_2793_));
 sky130_fd_sc_hd__clkbuf_1 _5598_ (.A(_2793_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(net579),
    .A1(_0762_),
    .S(_2785_),
    .X(_2794_));
 sky130_fd_sc_hd__clkbuf_1 _5600_ (.A(_2794_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _5601_ (.A0(net489),
    .A1(_0761_),
    .S(_2785_),
    .X(_2795_));
 sky130_fd_sc_hd__clkbuf_1 _5602_ (.A(_2795_),
    .X(_0420_));
 sky130_fd_sc_hd__buf_4 _5603_ (.A(_2750_),
    .X(_2796_));
 sky130_fd_sc_hd__mux2_1 _5604_ (.A0(net586),
    .A1(_1038_),
    .S(_2796_),
    .X(_2797_));
 sky130_fd_sc_hd__clkbuf_1 _5605_ (.A(_2797_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _5606_ (.A0(net198),
    .A1(_0734_),
    .S(_2796_),
    .X(_2798_));
 sky130_fd_sc_hd__clkbuf_1 _5607_ (.A(_2798_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _5608_ (.A0(net496),
    .A1(_0733_),
    .S(_2796_),
    .X(_2799_));
 sky130_fd_sc_hd__clkbuf_1 _5609_ (.A(_2799_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _5610_ (.A0(net341),
    .A1(_0732_),
    .S(_2796_),
    .X(_2800_));
 sky130_fd_sc_hd__clkbuf_1 _5611_ (.A(_2800_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _5612_ (.A0(net498),
    .A1(_0729_),
    .S(_2796_),
    .X(_2801_));
 sky130_fd_sc_hd__clkbuf_1 _5613_ (.A(_2801_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _5614_ (.A0(net339),
    .A1(_0730_),
    .S(_2796_),
    .X(_2802_));
 sky130_fd_sc_hd__clkbuf_1 _5615_ (.A(_2802_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _5616_ (.A0(net479),
    .A1(_1426_),
    .S(_2796_),
    .X(_2803_));
 sky130_fd_sc_hd__clkbuf_1 _5617_ (.A(_2803_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _5618_ (.A0(net234),
    .A1(_0727_),
    .S(_2796_),
    .X(_2804_));
 sky130_fd_sc_hd__clkbuf_1 _5619_ (.A(_2804_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _5620_ (.A0(net642),
    .A1(_0738_),
    .S(_2796_),
    .X(_2805_));
 sky130_fd_sc_hd__clkbuf_1 _5621_ (.A(_2805_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _5622_ (.A0(net293),
    .A1(_0737_),
    .S(_2796_),
    .X(_2806_));
 sky130_fd_sc_hd__clkbuf_1 _5623_ (.A(_2806_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _5624_ (.A0(net374),
    .A1(_1227_),
    .S(_2751_),
    .X(_2807_));
 sky130_fd_sc_hd__clkbuf_1 _5625_ (.A(_2807_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _5626_ (.A0(net388),
    .A1(_0739_),
    .S(_2751_),
    .X(_2808_));
 sky130_fd_sc_hd__clkbuf_1 _5627_ (.A(_2808_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _5628_ (.A0(net462),
    .A1(_0743_),
    .S(_2751_),
    .X(_2809_));
 sky130_fd_sc_hd__clkbuf_1 _5629_ (.A(_2809_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _5630_ (.A0(net519),
    .A1(_0741_),
    .S(_2751_),
    .X(_2810_));
 sky130_fd_sc_hd__clkbuf_1 _5631_ (.A(_2810_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _5632_ (.A0(net310),
    .A1(_0742_),
    .S(_2751_),
    .X(_2811_));
 sky130_fd_sc_hd__clkbuf_1 _5633_ (.A(_2811_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _5634_ (.A0(net415),
    .A1(_1954_),
    .S(_2751_),
    .X(_2812_));
 sky130_fd_sc_hd__clkbuf_1 _5635_ (.A(_2812_),
    .X(_0436_));
 sky130_fd_sc_hd__and3_1 _5636_ (.A(_0772_),
    .B(_0788_),
    .C(_0777_),
    .X(_2813_));
 sky130_fd_sc_hd__clkbuf_8 _5637_ (.A(_2813_),
    .X(_2814_));
 sky130_fd_sc_hd__buf_4 _5638_ (.A(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__mux2_1 _5639_ (.A0(net470),
    .A1(_1347_),
    .S(_2815_),
    .X(_2816_));
 sky130_fd_sc_hd__clkbuf_1 _5640_ (.A(_2816_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _5641_ (.A0(net301),
    .A1(_0943_),
    .S(_2815_),
    .X(_2817_));
 sky130_fd_sc_hd__clkbuf_1 _5642_ (.A(_2817_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _5643_ (.A0(net361),
    .A1(_0845_),
    .S(_2815_),
    .X(_2818_));
 sky130_fd_sc_hd__clkbuf_1 _5644_ (.A(_2818_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _5645_ (.A0(net229),
    .A1(_0705_),
    .S(_2815_),
    .X(_2819_));
 sky130_fd_sc_hd__clkbuf_1 _5646_ (.A(_2819_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _5647_ (.A0(net256),
    .A1(_0703_),
    .S(_2815_),
    .X(_2820_));
 sky130_fd_sc_hd__clkbuf_1 _5648_ (.A(_2820_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _5649_ (.A0(net210),
    .A1(_0702_),
    .S(_2815_),
    .X(_2821_));
 sky130_fd_sc_hd__clkbuf_1 _5650_ (.A(_2821_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _5651_ (.A0(net240),
    .A1(_1048_),
    .S(_2815_),
    .X(_2822_));
 sky130_fd_sc_hd__clkbuf_1 _5652_ (.A(_2822_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _5653_ (.A0(net670),
    .A1(_0847_),
    .S(_2815_),
    .X(_2823_));
 sky130_fd_sc_hd__clkbuf_1 _5654_ (.A(_2823_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _5655_ (.A0(net541),
    .A1(_0713_),
    .S(_2815_),
    .X(_2824_));
 sky130_fd_sc_hd__clkbuf_1 _5656_ (.A(_2824_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _5657_ (.A0(net282),
    .A1(_0714_),
    .S(_2815_),
    .X(_2825_));
 sky130_fd_sc_hd__clkbuf_1 _5658_ (.A(_2825_),
    .X(_0446_));
 sky130_fd_sc_hd__buf_4 _5659_ (.A(_2814_),
    .X(_2826_));
 sky130_fd_sc_hd__mux2_1 _5660_ (.A0(net402),
    .A1(_1518_),
    .S(_2826_),
    .X(_2827_));
 sky130_fd_sc_hd__clkbuf_1 _5661_ (.A(_2827_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _5662_ (.A0(net620),
    .A1(_0715_),
    .S(_2826_),
    .X(_2828_));
 sky130_fd_sc_hd__clkbuf_1 _5663_ (.A(_2828_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _5664_ (.A0(net290),
    .A1(_0708_),
    .S(_2826_),
    .X(_2829_));
 sky130_fd_sc_hd__clkbuf_1 _5665_ (.A(_2829_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _5666_ (.A0(net506),
    .A1(_0711_),
    .S(_2826_),
    .X(_2830_));
 sky130_fd_sc_hd__clkbuf_1 _5667_ (.A(_2830_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _5668_ (.A0(net584),
    .A1(_0710_),
    .S(_2826_),
    .X(_2831_));
 sky130_fd_sc_hd__clkbuf_1 _5669_ (.A(_2831_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _5670_ (.A0(net337),
    .A1(_0709_),
    .S(_2826_),
    .X(_2832_));
 sky130_fd_sc_hd__clkbuf_1 _5671_ (.A(_2832_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _5672_ (.A0(net577),
    .A1(_0880_),
    .S(_2826_),
    .X(_2833_));
 sky130_fd_sc_hd__clkbuf_1 _5673_ (.A(_2833_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _5674_ (.A0(net392),
    .A1(_0718_),
    .S(_2826_),
    .X(_2834_));
 sky130_fd_sc_hd__clkbuf_1 _5675_ (.A(_2834_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _5676_ (.A0(net297),
    .A1(_1493_),
    .S(_2826_),
    .X(_2835_));
 sky130_fd_sc_hd__clkbuf_1 _5677_ (.A(_2835_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _5678_ (.A0(net505),
    .A1(_0719_),
    .S(_2826_),
    .X(_2836_));
 sky130_fd_sc_hd__clkbuf_1 _5679_ (.A(_2836_),
    .X(_0456_));
 sky130_fd_sc_hd__buf_4 _5680_ (.A(_2814_),
    .X(_2837_));
 sky130_fd_sc_hd__mux2_1 _5681_ (.A0(net261),
    .A1(_0721_),
    .S(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__clkbuf_1 _5682_ (.A(_2838_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _5683_ (.A0(net278),
    .A1(_0724_),
    .S(_2837_),
    .X(_2839_));
 sky130_fd_sc_hd__clkbuf_1 _5684_ (.A(_2839_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _5685_ (.A0(net294),
    .A1(_0723_),
    .S(_2837_),
    .X(_2840_));
 sky130_fd_sc_hd__clkbuf_1 _5686_ (.A(_2840_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _5687_ (.A0(net562),
    .A1(_0722_),
    .S(_2837_),
    .X(_2841_));
 sky130_fd_sc_hd__clkbuf_1 _5688_ (.A(_2841_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _5689_ (.A0(net452),
    .A1(_0750_),
    .S(_2837_),
    .X(_2842_));
 sky130_fd_sc_hd__clkbuf_1 _5690_ (.A(_2842_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _5691_ (.A0(net366),
    .A1(_0752_),
    .S(_2837_),
    .X(_2843_));
 sky130_fd_sc_hd__clkbuf_1 _5692_ (.A(_2843_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _5693_ (.A0(net613),
    .A1(_0751_),
    .S(_2837_),
    .X(_2844_));
 sky130_fd_sc_hd__clkbuf_1 _5694_ (.A(_2844_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _5695_ (.A0(net262),
    .A1(_1731_),
    .S(_2837_),
    .X(_2845_));
 sky130_fd_sc_hd__clkbuf_1 _5696_ (.A(_2845_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _5697_ (.A0(net548),
    .A1(_0746_),
    .S(_2837_),
    .X(_2846_));
 sky130_fd_sc_hd__clkbuf_1 _5698_ (.A(_2846_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _5699_ (.A0(net423),
    .A1(_0748_),
    .S(_2837_),
    .X(_2847_));
 sky130_fd_sc_hd__clkbuf_1 _5700_ (.A(_2847_),
    .X(_0466_));
 sky130_fd_sc_hd__buf_4 _5701_ (.A(_2814_),
    .X(_2848_));
 sky130_fd_sc_hd__mux2_1 _5702_ (.A0(net380),
    .A1(_0857_),
    .S(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__clkbuf_1 _5703_ (.A(_2849_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _5704_ (.A0(net472),
    .A1(_0747_),
    .S(_2848_),
    .X(_2850_));
 sky130_fd_sc_hd__clkbuf_1 _5705_ (.A(_2850_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _5706_ (.A0(net421),
    .A1(_0755_),
    .S(_2848_),
    .X(_2851_));
 sky130_fd_sc_hd__clkbuf_1 _5707_ (.A(_2851_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _5708_ (.A0(net593),
    .A1(_0756_),
    .S(_2848_),
    .X(_2852_));
 sky130_fd_sc_hd__clkbuf_1 _5709_ (.A(_2852_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _5710_ (.A0(net281),
    .A1(_0757_),
    .S(_2848_),
    .X(_2853_));
 sky130_fd_sc_hd__clkbuf_1 _5711_ (.A(_2853_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _5712_ (.A0(net258),
    .A1(_0758_),
    .S(_2848_),
    .X(_2854_));
 sky130_fd_sc_hd__clkbuf_1 _5713_ (.A(_2854_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _5714_ (.A0(net614),
    .A1(_0760_),
    .S(_2848_),
    .X(_2855_));
 sky130_fd_sc_hd__clkbuf_1 _5715_ (.A(_2855_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _5716_ (.A0(net448),
    .A1(_0763_),
    .S(_2848_),
    .X(_2856_));
 sky130_fd_sc_hd__clkbuf_1 _5717_ (.A(_2856_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(net272),
    .A1(_0762_),
    .S(_2848_),
    .X(_2857_));
 sky130_fd_sc_hd__clkbuf_1 _5719_ (.A(_2857_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _5720_ (.A0(net630),
    .A1(_0761_),
    .S(_2848_),
    .X(_2858_));
 sky130_fd_sc_hd__clkbuf_1 _5721_ (.A(_2858_),
    .X(_0476_));
 sky130_fd_sc_hd__buf_4 _5722_ (.A(_2813_),
    .X(_2859_));
 sky130_fd_sc_hd__mux2_1 _5723_ (.A0(net200),
    .A1(_1038_),
    .S(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__clkbuf_1 _5724_ (.A(_2860_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _5725_ (.A0(net334),
    .A1(_0734_),
    .S(_2859_),
    .X(_2861_));
 sky130_fd_sc_hd__clkbuf_1 _5726_ (.A(_2861_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _5727_ (.A0(net203),
    .A1(_0733_),
    .S(_2859_),
    .X(_2862_));
 sky130_fd_sc_hd__clkbuf_1 _5728_ (.A(_2862_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _5729_ (.A0(net626),
    .A1(_0732_),
    .S(_2859_),
    .X(_2863_));
 sky130_fd_sc_hd__clkbuf_1 _5730_ (.A(_2863_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _5731_ (.A0(net638),
    .A1(_0729_),
    .S(_2859_),
    .X(_2864_));
 sky130_fd_sc_hd__clkbuf_1 _5732_ (.A(_2864_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _5733_ (.A0(net674),
    .A1(_0730_),
    .S(_2859_),
    .X(_2865_));
 sky130_fd_sc_hd__clkbuf_1 _5734_ (.A(_2865_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _5735_ (.A0(net242),
    .A1(_1426_),
    .S(_2859_),
    .X(_2866_));
 sky130_fd_sc_hd__clkbuf_1 _5736_ (.A(_2866_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _5737_ (.A0(net244),
    .A1(_0727_),
    .S(_2859_),
    .X(_2867_));
 sky130_fd_sc_hd__clkbuf_1 _5738_ (.A(_2867_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _5739_ (.A0(net443),
    .A1(_0738_),
    .S(_2859_),
    .X(_2868_));
 sky130_fd_sc_hd__clkbuf_1 _5740_ (.A(_2868_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _5741_ (.A0(net549),
    .A1(_0737_),
    .S(_2859_),
    .X(_2869_));
 sky130_fd_sc_hd__clkbuf_1 _5742_ (.A(_2869_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _5743_ (.A0(net375),
    .A1(_1227_),
    .S(_2814_),
    .X(_2870_));
 sky130_fd_sc_hd__clkbuf_1 _5744_ (.A(_2870_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _5745_ (.A0(net587),
    .A1(_0739_),
    .S(_2814_),
    .X(_2871_));
 sky130_fd_sc_hd__clkbuf_1 _5746_ (.A(_2871_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _5747_ (.A0(net325),
    .A1(_0743_),
    .S(_2814_),
    .X(_2872_));
 sky130_fd_sc_hd__clkbuf_1 _5748_ (.A(_2872_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _5749_ (.A0(net478),
    .A1(_0741_),
    .S(_2814_),
    .X(_2873_));
 sky130_fd_sc_hd__clkbuf_1 _5750_ (.A(_2873_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _5751_ (.A0(net460),
    .A1(_0742_),
    .S(_2814_),
    .X(_2874_));
 sky130_fd_sc_hd__clkbuf_1 _5752_ (.A(_2874_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _5753_ (.A0(net255),
    .A1(_1954_),
    .S(_2814_),
    .X(_2875_));
 sky130_fd_sc_hd__clkbuf_1 _5754_ (.A(_2875_),
    .X(_0492_));
 sky130_fd_sc_hd__or2_1 _5755_ (.A(_0772_),
    .B(_0771_),
    .X(_2876_));
 sky130_fd_sc_hd__clkbuf_8 _5756_ (.A(_2876_),
    .X(_2877_));
 sky130_fd_sc_hd__buf_4 _5757_ (.A(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__mux2_1 _5758_ (.A0(_1347_),
    .A1(net308),
    .S(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__clkbuf_1 _5759_ (.A(_2879_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _5760_ (.A0(_0943_),
    .A1(net523),
    .S(_2878_),
    .X(_2880_));
 sky130_fd_sc_hd__clkbuf_1 _5761_ (.A(_2880_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _5762_ (.A0(_0845_),
    .A1(net390),
    .S(_2878_),
    .X(_2881_));
 sky130_fd_sc_hd__clkbuf_1 _5763_ (.A(_2881_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _5764_ (.A0(_0705_),
    .A1(net551),
    .S(_2878_),
    .X(_2882_));
 sky130_fd_sc_hd__clkbuf_1 _5765_ (.A(_2882_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _5766_ (.A0(_0703_),
    .A1(net608),
    .S(_2878_),
    .X(_2883_));
 sky130_fd_sc_hd__clkbuf_1 _5767_ (.A(_2883_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _5768_ (.A0(_0702_),
    .A1(net471),
    .S(_2878_),
    .X(_2884_));
 sky130_fd_sc_hd__clkbuf_1 _5769_ (.A(_2884_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _5770_ (.A0(_1048_),
    .A1(net560),
    .S(_2878_),
    .X(_2885_));
 sky130_fd_sc_hd__clkbuf_1 _5771_ (.A(_2885_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _5772_ (.A0(_0847_),
    .A1(net667),
    .S(_2878_),
    .X(_2886_));
 sky130_fd_sc_hd__clkbuf_1 _5773_ (.A(_2886_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _5774_ (.A0(_0713_),
    .A1(net647),
    .S(_2878_),
    .X(_2887_));
 sky130_fd_sc_hd__clkbuf_1 _5775_ (.A(_2887_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _5776_ (.A0(_0714_),
    .A1(net540),
    .S(_2878_),
    .X(_2888_));
 sky130_fd_sc_hd__clkbuf_1 _5777_ (.A(_2888_),
    .X(_0502_));
 sky130_fd_sc_hd__buf_4 _5778_ (.A(_2877_),
    .X(_2889_));
 sky130_fd_sc_hd__mux2_1 _5779_ (.A0(_1518_),
    .A1(net476),
    .S(_2889_),
    .X(_2890_));
 sky130_fd_sc_hd__clkbuf_1 _5780_ (.A(_2890_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(_0715_),
    .A1(net657),
    .S(_2889_),
    .X(_2891_));
 sky130_fd_sc_hd__clkbuf_1 _5782_ (.A(_2891_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _5783_ (.A0(_0708_),
    .A1(net457),
    .S(_2889_),
    .X(_2892_));
 sky130_fd_sc_hd__clkbuf_1 _5784_ (.A(_2892_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _5785_ (.A0(_0711_),
    .A1(net413),
    .S(_2889_),
    .X(_2893_));
 sky130_fd_sc_hd__clkbuf_1 _5786_ (.A(_2893_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(_0710_),
    .A1(net490),
    .S(_2889_),
    .X(_2894_));
 sky130_fd_sc_hd__clkbuf_1 _5788_ (.A(_2894_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(_0709_),
    .A1(net313),
    .S(_2889_),
    .X(_2895_));
 sky130_fd_sc_hd__clkbuf_1 _5790_ (.A(_2895_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _5791_ (.A0(_0880_),
    .A1(net482),
    .S(_2889_),
    .X(_2896_));
 sky130_fd_sc_hd__clkbuf_1 _5792_ (.A(_2896_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _5793_ (.A0(_0718_),
    .A1(net616),
    .S(_2889_),
    .X(_2897_));
 sky130_fd_sc_hd__clkbuf_1 _5794_ (.A(_2897_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _5795_ (.A0(_1493_),
    .A1(net544),
    .S(_2889_),
    .X(_2898_));
 sky130_fd_sc_hd__clkbuf_1 _5796_ (.A(_2898_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(_0719_),
    .A1(net641),
    .S(_2889_),
    .X(_2899_));
 sky130_fd_sc_hd__clkbuf_1 _5798_ (.A(_2899_),
    .X(_0512_));
 sky130_fd_sc_hd__buf_4 _5799_ (.A(_2877_),
    .X(_2900_));
 sky130_fd_sc_hd__mux2_1 _5800_ (.A0(_0721_),
    .A1(net571),
    .S(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__clkbuf_1 _5801_ (.A(_2901_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _5802_ (.A0(_0724_),
    .A1(net637),
    .S(_2900_),
    .X(_2902_));
 sky130_fd_sc_hd__clkbuf_1 _5803_ (.A(_2902_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _5804_ (.A0(_0723_),
    .A1(net449),
    .S(_2900_),
    .X(_2903_));
 sky130_fd_sc_hd__clkbuf_1 _5805_ (.A(_2903_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _5806_ (.A0(_0722_),
    .A1(net665),
    .S(_2900_),
    .X(_2904_));
 sky130_fd_sc_hd__clkbuf_1 _5807_ (.A(_2904_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _5808_ (.A0(_0750_),
    .A1(net639),
    .S(_2900_),
    .X(_2905_));
 sky130_fd_sc_hd__clkbuf_1 _5809_ (.A(_2905_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _5810_ (.A0(_0752_),
    .A1(net633),
    .S(_2900_),
    .X(_2906_));
 sky130_fd_sc_hd__clkbuf_1 _5811_ (.A(_2906_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _5812_ (.A0(_0751_),
    .A1(net660),
    .S(_2900_),
    .X(_2907_));
 sky130_fd_sc_hd__clkbuf_1 _5813_ (.A(_2907_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _5814_ (.A0(_1731_),
    .A1(net580),
    .S(_2900_),
    .X(_2908_));
 sky130_fd_sc_hd__clkbuf_1 _5815_ (.A(_2908_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _5816_ (.A0(_0746_),
    .A1(net654),
    .S(_2900_),
    .X(_2909_));
 sky130_fd_sc_hd__clkbuf_1 _5817_ (.A(_2909_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _5818_ (.A0(_0748_),
    .A1(net617),
    .S(_2900_),
    .X(_2910_));
 sky130_fd_sc_hd__clkbuf_1 _5819_ (.A(_2910_),
    .X(_0522_));
 sky130_fd_sc_hd__buf_4 _5820_ (.A(_2877_),
    .X(_2911_));
 sky130_fd_sc_hd__mux2_1 _5821_ (.A0(_0857_),
    .A1(net416),
    .S(_2911_),
    .X(_2912_));
 sky130_fd_sc_hd__clkbuf_1 _5822_ (.A(_2912_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _5823_ (.A0(_0747_),
    .A1(net533),
    .S(_2911_),
    .X(_2913_));
 sky130_fd_sc_hd__clkbuf_1 _5824_ (.A(_2913_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _5825_ (.A0(_0755_),
    .A1(net414),
    .S(_2911_),
    .X(_2914_));
 sky130_fd_sc_hd__clkbuf_1 _5826_ (.A(_2914_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _5827_ (.A0(_0756_),
    .A1(net538),
    .S(_2911_),
    .X(_2915_));
 sky130_fd_sc_hd__clkbuf_1 _5828_ (.A(_2915_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _5829_ (.A0(_0757_),
    .A1(net570),
    .S(_2911_),
    .X(_2916_));
 sky130_fd_sc_hd__clkbuf_1 _5830_ (.A(_2916_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _5831_ (.A0(_0758_),
    .A1(net483),
    .S(_2911_),
    .X(_2917_));
 sky130_fd_sc_hd__clkbuf_1 _5832_ (.A(_2917_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _5833_ (.A0(_0760_),
    .A1(net588),
    .S(_2911_),
    .X(_2918_));
 sky130_fd_sc_hd__clkbuf_1 _5834_ (.A(_2918_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _5835_ (.A0(_0763_),
    .A1(net426),
    .S(_2911_),
    .X(_2919_));
 sky130_fd_sc_hd__clkbuf_1 _5836_ (.A(_2919_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _5837_ (.A0(_0762_),
    .A1(net525),
    .S(_2911_),
    .X(_2920_));
 sky130_fd_sc_hd__clkbuf_1 _5838_ (.A(_2920_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _5839_ (.A0(_0761_),
    .A1(net503),
    .S(_2911_),
    .X(_2921_));
 sky130_fd_sc_hd__clkbuf_1 _5840_ (.A(_2921_),
    .X(_0532_));
 sky130_fd_sc_hd__buf_4 _5841_ (.A(_2876_),
    .X(_2922_));
 sky130_fd_sc_hd__mux2_1 _5842_ (.A0(_1038_),
    .A1(net419),
    .S(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__clkbuf_1 _5843_ (.A(_2923_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _5844_ (.A0(_0734_),
    .A1(net634),
    .S(_2922_),
    .X(_2924_));
 sky130_fd_sc_hd__clkbuf_1 _5845_ (.A(_2924_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _5846_ (.A0(_0733_),
    .A1(net517),
    .S(_2922_),
    .X(_2925_));
 sky130_fd_sc_hd__clkbuf_1 _5847_ (.A(_2925_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _5848_ (.A0(_0732_),
    .A1(net612),
    .S(_2922_),
    .X(_2926_));
 sky130_fd_sc_hd__clkbuf_1 _5849_ (.A(_2926_),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _5850_ (.A0(_0729_),
    .A1(net658),
    .S(_2922_),
    .X(_2927_));
 sky130_fd_sc_hd__clkbuf_1 _5851_ (.A(_2927_),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _5852_ (.A0(_0730_),
    .A1(net676),
    .S(_2922_),
    .X(_2928_));
 sky130_fd_sc_hd__clkbuf_1 _5853_ (.A(_2928_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _5854_ (.A0(_1426_),
    .A1(net644),
    .S(_2922_),
    .X(_2929_));
 sky130_fd_sc_hd__clkbuf_1 _5855_ (.A(_2929_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _5856_ (.A0(_0727_),
    .A1(net677),
    .S(_2922_),
    .X(_2930_));
 sky130_fd_sc_hd__clkbuf_1 _5857_ (.A(_2930_),
    .X(_0540_));
 sky130_fd_sc_hd__mux2_1 _5858_ (.A0(_0738_),
    .A1(net609),
    .S(_2922_),
    .X(_2931_));
 sky130_fd_sc_hd__clkbuf_1 _5859_ (.A(_2931_),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _5860_ (.A0(_0737_),
    .A1(net430),
    .S(_2922_),
    .X(_2932_));
 sky130_fd_sc_hd__clkbuf_1 _5861_ (.A(_2932_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _5862_ (.A0(_1227_),
    .A1(net445),
    .S(_2877_),
    .X(_2933_));
 sky130_fd_sc_hd__clkbuf_1 _5863_ (.A(_2933_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _5864_ (.A0(_0739_),
    .A1(net456),
    .S(_2877_),
    .X(_2934_));
 sky130_fd_sc_hd__clkbuf_1 _5865_ (.A(_2934_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _5866_ (.A0(_0743_),
    .A1(net404),
    .S(_2877_),
    .X(_2935_));
 sky130_fd_sc_hd__clkbuf_1 _5867_ (.A(_2935_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _5868_ (.A0(_0741_),
    .A1(net664),
    .S(_2877_),
    .X(_2936_));
 sky130_fd_sc_hd__clkbuf_1 _5869_ (.A(_2936_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _5870_ (.A0(_0742_),
    .A1(net358),
    .S(_2877_),
    .X(_2937_));
 sky130_fd_sc_hd__clkbuf_1 _5871_ (.A(_2937_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _5872_ (.A0(_1954_),
    .A1(net369),
    .S(_2877_),
    .X(_2938_));
 sky130_fd_sc_hd__clkbuf_1 _5873_ (.A(_2938_),
    .X(_0548_));
 sky130_fd_sc_hd__inv_2 _5874_ (.A(_2749_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _5875_ (.A(_2749_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _5876_ (.A(_2749_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _5877_ (.A(_2749_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _5878_ (.A(_2749_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _5879_ (.A(_2749_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _5880_ (.A(_2749_),
    .Y(_0009_));
 sky130_fd_sc_hd__clkbuf_8 _5881_ (.A(_2748_),
    .X(_2939_));
 sky130_fd_sc_hd__inv_2 _5882_ (.A(_2939_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _5883_ (.A(_2939_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _5884_ (.A(_2939_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _5885_ (.A(_2939_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _5886_ (.A(_2939_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _5887_ (.A(_2939_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _5888_ (.A(_2939_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _5889_ (.A(_2939_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _5890_ (.A(_2939_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _5891_ (.A(_2939_),
    .Y(_0019_));
 sky130_fd_sc_hd__clkbuf_8 _5892_ (.A(_2748_),
    .X(_2940_));
 sky130_fd_sc_hd__inv_2 _5893_ (.A(_2940_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _5894_ (.A(_2940_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _5895_ (.A(_2940_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _5896_ (.A(_2940_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _5897_ (.A(_2940_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _5898_ (.A(_2940_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _5899_ (.A(_2940_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _5900_ (.A(_2940_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _5901_ (.A(_2940_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _5902_ (.A(_2940_),
    .Y(_0029_));
 sky130_fd_sc_hd__buf_6 _5903_ (.A(net123),
    .X(_2941_));
 sky130_fd_sc_hd__inv_2 _5904_ (.A(_2941_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _5905_ (.A(_2941_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _5906_ (.A(_2941_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _5907_ (.A(_2941_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _5908_ (.A(_2941_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _5909_ (.A(_2941_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _5910_ (.A(_2941_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _5911_ (.A(_2941_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _5912_ (.A(_2941_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _5913_ (.A(_2941_),
    .Y(_0039_));
 sky130_fd_sc_hd__clkbuf_8 _5914_ (.A(net123),
    .X(_2942_));
 sky130_fd_sc_hd__inv_2 _5915_ (.A(_2942_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _5916_ (.A(_2942_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _5917_ (.A(_2942_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _5918_ (.A(_2942_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _5919_ (.A(_2942_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _5920_ (.A(_2942_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _5921_ (.A(_2942_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _5922_ (.A(_2942_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _5923_ (.A(_2942_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _5924_ (.A(_2942_),
    .Y(_0049_));
 sky130_fd_sc_hd__clkbuf_8 _5925_ (.A(net123),
    .X(_2943_));
 sky130_fd_sc_hd__inv_2 _5926_ (.A(_2943_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _5927_ (.A(_2943_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _5928_ (.A(_2943_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _5929_ (.A(_2943_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _5930_ (.A(_2943_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _5931_ (.A(_2943_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _5932_ (.A(_2943_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _5933_ (.A(_2943_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _5934_ (.A(_2943_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _5935_ (.A(_2943_),
    .Y(_0059_));
 sky130_fd_sc_hd__clkbuf_8 _5936_ (.A(net123),
    .X(_2944_));
 sky130_fd_sc_hd__inv_2 _5937_ (.A(_2944_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _5938_ (.A(_2944_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _5939_ (.A(_2944_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _5940_ (.A(_2944_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _5941_ (.A(_2944_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _5942_ (.A(_2944_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _5943_ (.A(_2944_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _5944_ (.A(_2944_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _5945_ (.A(_2944_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _5946_ (.A(_2944_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _5947_ (.A(_2748_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _5948_ (.A(_2748_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _5949_ (.A(_2748_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _5950_ (.A(_2748_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _5951_ (.A(_2748_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _5952_ (.A(_2748_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _5953_ (.A(_2748_),
    .Y(_0076_));
 sky130_fd_sc_hd__dfxtp_1 _5954_ (.CLK(clknet_leaf_32_clk),
    .D(_0623_),
    .Q(\fifo.fifo[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5955_ (.CLK(clknet_leaf_26_clk),
    .D(_0624_),
    .Q(\fifo.fifo[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5956_ (.CLK(clknet_leaf_27_clk),
    .D(_0625_),
    .Q(\fifo.fifo[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5957_ (.CLK(clknet_leaf_28_clk),
    .D(_0626_),
    .Q(\fifo.fifo[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5958_ (.CLK(clknet_leaf_30_clk),
    .D(_0627_),
    .Q(\fifo.fifo[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5959_ (.CLK(clknet_leaf_30_clk),
    .D(_0628_),
    .Q(\fifo.fifo[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5960_ (.CLK(clknet_leaf_27_clk),
    .D(_0629_),
    .Q(\fifo.fifo[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5961_ (.CLK(clknet_leaf_18_clk),
    .D(_0630_),
    .Q(\fifo.fifo[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5962_ (.CLK(clknet_leaf_17_clk),
    .D(_0631_),
    .Q(\fifo.fifo[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _5963_ (.CLK(clknet_leaf_20_clk),
    .D(_0632_),
    .Q(\fifo.fifo[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _5964_ (.CLK(clknet_leaf_15_clk),
    .D(_0633_),
    .Q(\fifo.fifo[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _5965_ (.CLK(clknet_leaf_17_clk),
    .D(_0634_),
    .Q(\fifo.fifo[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _5966_ (.CLK(clknet_leaf_15_clk),
    .D(_0635_),
    .Q(\fifo.fifo[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _5967_ (.CLK(clknet_leaf_12_clk),
    .D(_0636_),
    .Q(\fifo.fifo[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _5968_ (.CLK(clknet_leaf_13_clk),
    .D(_0637_),
    .Q(\fifo.fifo[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _5969_ (.CLK(clknet_leaf_16_clk),
    .D(_0638_),
    .Q(\fifo.fifo[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _5970_ (.CLK(clknet_leaf_12_clk),
    .D(_0639_),
    .Q(\fifo.fifo[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _5971_ (.CLK(clknet_leaf_9_clk),
    .D(_0640_),
    .Q(\fifo.fifo[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _5972_ (.CLK(clknet_leaf_9_clk),
    .D(_0641_),
    .Q(\fifo.fifo[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _5973_ (.CLK(clknet_leaf_10_clk),
    .D(_0642_),
    .Q(\fifo.fifo[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _5974_ (.CLK(clknet_leaf_1_clk),
    .D(_0643_),
    .Q(\fifo.fifo[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _5975_ (.CLK(clknet_leaf_0_clk),
    .D(_0644_),
    .Q(\fifo.fifo[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _5976_ (.CLK(clknet_leaf_69_clk),
    .D(_0645_),
    .Q(\fifo.fifo[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _5977_ (.CLK(clknet_leaf_0_clk),
    .D(_0646_),
    .Q(\fifo.fifo[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _5978_ (.CLK(clknet_leaf_2_clk),
    .D(_0647_),
    .Q(\fifo.fifo[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _5979_ (.CLK(clknet_leaf_0_clk),
    .D(_0648_),
    .Q(\fifo.fifo[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _5980_ (.CLK(clknet_leaf_3_clk),
    .D(_0649_),
    .Q(\fifo.fifo[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _5981_ (.CLK(clknet_leaf_2_clk),
    .D(_0650_),
    .Q(\fifo.fifo[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _5982_ (.CLK(clknet_leaf_68_clk),
    .D(_0651_),
    .Q(\fifo.fifo[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _5983_ (.CLK(clknet_leaf_3_clk),
    .D(_0652_),
    .Q(\fifo.fifo[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _5984_ (.CLK(clknet_leaf_66_clk),
    .D(_0653_),
    .Q(\fifo.fifo[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _5985_ (.CLK(clknet_leaf_65_clk),
    .D(_0654_),
    .Q(\fifo.fifo[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _5986_ (.CLK(clknet_leaf_64_clk),
    .D(_0655_),
    .Q(\fifo.fifo[5][32] ));
 sky130_fd_sc_hd__dfxtp_1 _5987_ (.CLK(clknet_leaf_64_clk),
    .D(_0656_),
    .Q(\fifo.fifo[5][33] ));
 sky130_fd_sc_hd__dfxtp_1 _5988_ (.CLK(clknet_leaf_64_clk),
    .D(_0657_),
    .Q(\fifo.fifo[5][34] ));
 sky130_fd_sc_hd__dfxtp_1 _5989_ (.CLK(clknet_leaf_67_clk),
    .D(_0077_),
    .Q(\fifo.fifo[5][35] ));
 sky130_fd_sc_hd__dfxtp_1 _5990_ (.CLK(clknet_leaf_62_clk),
    .D(_0078_),
    .Q(\fifo.fifo[5][36] ));
 sky130_fd_sc_hd__dfxtp_1 _5991_ (.CLK(clknet_leaf_63_clk),
    .D(_0079_),
    .Q(\fifo.fifo[5][37] ));
 sky130_fd_sc_hd__dfxtp_1 _5992_ (.CLK(clknet_leaf_62_clk),
    .D(_0080_),
    .Q(\fifo.fifo[5][38] ));
 sky130_fd_sc_hd__dfxtp_1 _5993_ (.CLK(clknet_leaf_62_clk),
    .D(_0081_),
    .Q(\fifo.fifo[5][39] ));
 sky130_fd_sc_hd__dfxtp_1 _5994_ (.CLK(clknet_leaf_52_clk),
    .D(_0082_),
    .Q(\fifo.fifo[5][40] ));
 sky130_fd_sc_hd__dfxtp_1 _5995_ (.CLK(clknet_leaf_51_clk),
    .D(_0083_),
    .Q(\fifo.fifo[5][41] ));
 sky130_fd_sc_hd__dfxtp_1 _5996_ (.CLK(clknet_leaf_49_clk),
    .D(_0084_),
    .Q(\fifo.fifo[5][42] ));
 sky130_fd_sc_hd__dfxtp_1 _5997_ (.CLK(clknet_leaf_48_clk),
    .D(_0085_),
    .Q(\fifo.fifo[5][43] ));
 sky130_fd_sc_hd__dfxtp_1 _5998_ (.CLK(clknet_leaf_48_clk),
    .D(_0086_),
    .Q(\fifo.fifo[5][44] ));
 sky130_fd_sc_hd__dfxtp_1 _5999_ (.CLK(clknet_leaf_47_clk),
    .D(_0087_),
    .Q(\fifo.fifo[5][45] ));
 sky130_fd_sc_hd__dfxtp_1 _6000_ (.CLK(clknet_leaf_44_clk),
    .D(_0088_),
    .Q(\fifo.fifo[5][46] ));
 sky130_fd_sc_hd__dfxtp_1 _6001_ (.CLK(clknet_leaf_44_clk),
    .D(_0089_),
    .Q(\fifo.fifo[5][47] ));
 sky130_fd_sc_hd__dfxtp_1 _6002_ (.CLK(clknet_leaf_49_clk),
    .D(_0090_),
    .Q(\fifo.fifo[5][48] ));
 sky130_fd_sc_hd__dfxtp_1 _6003_ (.CLK(clknet_leaf_50_clk),
    .D(_0091_),
    .Q(\fifo.fifo[5][49] ));
 sky130_fd_sc_hd__dfxtp_1 _6004_ (.CLK(clknet_leaf_54_clk),
    .D(_0092_),
    .Q(\fifo.fifo[5][50] ));
 sky130_fd_sc_hd__dfxtp_1 _6005_ (.CLK(clknet_leaf_56_clk),
    .D(_0093_),
    .Q(\fifo.fifo[5][51] ));
 sky130_fd_sc_hd__dfxtp_1 _6006_ (.CLK(clknet_leaf_55_clk),
    .D(_0094_),
    .Q(\fifo.fifo[5][52] ));
 sky130_fd_sc_hd__dfxtp_1 _6007_ (.CLK(clknet_leaf_58_clk),
    .D(_0095_),
    .Q(\fifo.fifo[5][53] ));
 sky130_fd_sc_hd__dfxtp_1 _6008_ (.CLK(clknet_leaf_62_clk),
    .D(_0096_),
    .Q(\fifo.fifo[5][54] ));
 sky130_fd_sc_hd__dfxtp_1 _6009_ (.CLK(clknet_leaf_61_clk),
    .D(_0097_),
    .Q(\fifo.fifo[5][55] ));
 sky130_fd_sc_hd__dfxtp_1 _6010_ (.CLK(clknet_leaf_31_clk),
    .D(_0098_),
    .Q(\fifo.rd_data[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6011_ (.CLK(clknet_leaf_26_clk),
    .D(_0099_),
    .Q(\fifo.rd_data[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6012_ (.CLK(clknet_leaf_32_clk),
    .D(_0100_),
    .Q(\fifo.rd_data[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6013_ (.CLK(clknet_leaf_27_clk),
    .D(_0101_),
    .Q(\fifo.rd_data[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6014_ (.CLK(clknet_leaf_32_clk),
    .D(_0102_),
    .Q(\fifo.rd_data[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6015_ (.CLK(clknet_leaf_32_clk),
    .D(_0103_),
    .Q(\fifo.rd_data[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6016_ (.CLK(clknet_leaf_19_clk),
    .D(_0104_),
    .Q(\fifo.rd_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6017_ (.CLK(clknet_leaf_18_clk),
    .D(_0105_),
    .Q(\fifo.rd_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6018_ (.CLK(clknet_leaf_18_clk),
    .D(_0106_),
    .Q(\fifo.rd_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6019_ (.CLK(clknet_leaf_20_clk),
    .D(_0107_),
    .Q(\fifo.rd_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6020_ (.CLK(clknet_leaf_17_clk),
    .D(_0108_),
    .Q(\fifo.rd_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6021_ (.CLK(clknet_leaf_16_clk),
    .D(_0109_),
    .Q(\fifo.rd_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6022_ (.CLK(clknet_leaf_16_clk),
    .D(_0110_),
    .Q(\fifo.rd_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6023_ (.CLK(clknet_leaf_21_clk),
    .D(_0111_),
    .Q(\fifo.rd_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6024_ (.CLK(clknet_leaf_20_clk),
    .D(_0112_),
    .Q(\fifo.rd_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6025_ (.CLK(clknet_leaf_20_clk),
    .D(_0113_),
    .Q(\fifo.rd_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6026_ (.CLK(clknet_leaf_8_clk),
    .D(_0114_),
    .Q(\fifo.rd_data[16] ));
 sky130_fd_sc_hd__dfxtp_1 _6027_ (.CLK(clknet_leaf_8_clk),
    .D(_0115_),
    .Q(\fifo.rd_data[17] ));
 sky130_fd_sc_hd__dfxtp_1 _6028_ (.CLK(clknet_leaf_8_clk),
    .D(_0116_),
    .Q(\fifo.rd_data[18] ));
 sky130_fd_sc_hd__dfxtp_1 _6029_ (.CLK(clknet_leaf_9_clk),
    .D(_0117_),
    .Q(\fifo.rd_data[19] ));
 sky130_fd_sc_hd__dfxtp_1 _6030_ (.CLK(clknet_leaf_10_clk),
    .D(_0118_),
    .Q(\fifo.rd_data[20] ));
 sky130_fd_sc_hd__dfxtp_1 _6031_ (.CLK(clknet_leaf_10_clk),
    .D(_0119_),
    .Q(\fifo.rd_data[21] ));
 sky130_fd_sc_hd__dfxtp_1 _6032_ (.CLK(clknet_leaf_9_clk),
    .D(_0120_),
    .Q(\fifo.rd_data[22] ));
 sky130_fd_sc_hd__dfxtp_1 _6033_ (.CLK(clknet_leaf_10_clk),
    .D(_0121_),
    .Q(\fifo.rd_data[23] ));
 sky130_fd_sc_hd__dfxtp_1 _6034_ (.CLK(clknet_leaf_9_clk),
    .D(_0122_),
    .Q(\fifo.rd_data[24] ));
 sky130_fd_sc_hd__dfxtp_1 _6035_ (.CLK(clknet_leaf_10_clk),
    .D(_0123_),
    .Q(\fifo.rd_data[25] ));
 sky130_fd_sc_hd__dfxtp_1 _6036_ (.CLK(clknet_leaf_6_clk),
    .D(_0124_),
    .Q(\fifo.rd_data[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6037_ (.CLK(clknet_leaf_4_clk),
    .D(_0125_),
    .Q(\fifo.rd_data[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6038_ (.CLK(clknet_leaf_2_clk),
    .D(_0126_),
    .Q(\fifo.rd_data[28] ));
 sky130_fd_sc_hd__dfxtp_1 _6039_ (.CLK(clknet_leaf_60_clk),
    .D(_0127_),
    .Q(\fifo.rd_data[29] ));
 sky130_fd_sc_hd__dfxtp_1 _6040_ (.CLK(clknet_leaf_66_clk),
    .D(_0128_),
    .Q(\fifo.rd_data[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6041_ (.CLK(clknet_leaf_60_clk),
    .D(_0129_),
    .Q(\fifo.rd_data[31] ));
 sky130_fd_sc_hd__dfxtp_1 _6042_ (.CLK(clknet_leaf_61_clk),
    .D(_0130_),
    .Q(\fifo.rd_data[32] ));
 sky130_fd_sc_hd__dfxtp_1 _6043_ (.CLK(clknet_leaf_60_clk),
    .D(_0131_),
    .Q(\fifo.rd_data[33] ));
 sky130_fd_sc_hd__dfxtp_1 _6044_ (.CLK(clknet_leaf_59_clk),
    .D(_0132_),
    .Q(\fifo.rd_data[34] ));
 sky130_fd_sc_hd__dfxtp_1 _6045_ (.CLK(clknet_leaf_60_clk),
    .D(_0133_),
    .Q(\fifo.rd_data[35] ));
 sky130_fd_sc_hd__dfxtp_1 _6046_ (.CLK(clknet_leaf_57_clk),
    .D(_0134_),
    .Q(\fifo.rd_data[36] ));
 sky130_fd_sc_hd__dfxtp_1 _6047_ (.CLK(clknet_leaf_57_clk),
    .D(_0135_),
    .Q(\fifo.rd_data[37] ));
 sky130_fd_sc_hd__dfxtp_1 _6048_ (.CLK(clknet_leaf_57_clk),
    .D(_0136_),
    .Q(\fifo.rd_data[38] ));
 sky130_fd_sc_hd__dfxtp_1 _6049_ (.CLK(clknet_leaf_42_clk),
    .D(_0137_),
    .Q(\fifo.rd_data[39] ));
 sky130_fd_sc_hd__dfxtp_1 _6050_ (.CLK(clknet_leaf_42_clk),
    .D(_0138_),
    .Q(\fifo.rd_data[40] ));
 sky130_fd_sc_hd__dfxtp_1 _6051_ (.CLK(clknet_leaf_44_clk),
    .D(_0139_),
    .Q(\fifo.rd_data[41] ));
 sky130_fd_sc_hd__dfxtp_1 _6052_ (.CLK(clknet_leaf_42_clk),
    .D(_0140_),
    .Q(\fifo.rd_data[42] ));
 sky130_fd_sc_hd__dfxtp_1 _6053_ (.CLK(clknet_leaf_42_clk),
    .D(_0141_),
    .Q(\fifo.rd_data[43] ));
 sky130_fd_sc_hd__dfxtp_1 _6054_ (.CLK(clknet_leaf_43_clk),
    .D(_0142_),
    .Q(\fifo.rd_data[44] ));
 sky130_fd_sc_hd__dfxtp_1 _6055_ (.CLK(clknet_leaf_41_clk),
    .D(_0143_),
    .Q(\fifo.rd_data[45] ));
 sky130_fd_sc_hd__dfxtp_1 _6056_ (.CLK(clknet_leaf_42_clk),
    .D(_0144_),
    .Q(\fifo.rd_data[46] ));
 sky130_fd_sc_hd__dfxtp_1 _6057_ (.CLK(clknet_leaf_42_clk),
    .D(_0145_),
    .Q(\fifo.rd_data[47] ));
 sky130_fd_sc_hd__dfxtp_1 _6058_ (.CLK(clknet_leaf_43_clk),
    .D(_0146_),
    .Q(\fifo.rd_data[48] ));
 sky130_fd_sc_hd__dfxtp_1 _6059_ (.CLK(clknet_leaf_50_clk),
    .D(_0147_),
    .Q(\fifo.rd_data[49] ));
 sky130_fd_sc_hd__dfxtp_1 _6060_ (.CLK(clknet_leaf_44_clk),
    .D(_0148_),
    .Q(\fifo.rd_data[50] ));
 sky130_fd_sc_hd__dfxtp_1 _6061_ (.CLK(clknet_leaf_50_clk),
    .D(_0149_),
    .Q(\fifo.rd_data[51] ));
 sky130_fd_sc_hd__dfxtp_1 _6062_ (.CLK(clknet_leaf_38_clk),
    .D(_0150_),
    .Q(\fifo.rd_data[52] ));
 sky130_fd_sc_hd__dfxtp_1 _6063_ (.CLK(clknet_leaf_38_clk),
    .D(_0151_),
    .Q(\fifo.rd_data[53] ));
 sky130_fd_sc_hd__dfxtp_1 _6064_ (.CLK(clknet_leaf_56_clk),
    .D(_0152_),
    .Q(\fifo.rd_data[54] ));
 sky130_fd_sc_hd__dfxtp_1 _6065_ (.CLK(clknet_leaf_38_clk),
    .D(_0153_),
    .Q(\fifo.rd_data[55] ));
 sky130_fd_sc_hd__dfxtp_1 _6066_ (.CLK(clknet_leaf_26_clk),
    .D(_0154_),
    .Q(\fifo.fifo[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6067_ (.CLK(clknet_leaf_19_clk),
    .D(_0155_),
    .Q(\fifo.fifo[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6068_ (.CLK(clknet_leaf_28_clk),
    .D(_0156_),
    .Q(\fifo.fifo[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6069_ (.CLK(clknet_leaf_28_clk),
    .D(_0157_),
    .Q(\fifo.fifo[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6070_ (.CLK(clknet_leaf_29_clk),
    .D(_0158_),
    .Q(\fifo.fifo[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6071_ (.CLK(clknet_leaf_29_clk),
    .D(_0159_),
    .Q(\fifo.fifo[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6072_ (.CLK(clknet_leaf_18_clk),
    .D(_0160_),
    .Q(\fifo.fifo[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6073_ (.CLK(clknet_leaf_18_clk),
    .D(_0161_),
    .Q(\fifo.fifo[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6074_ (.CLK(clknet_leaf_17_clk),
    .D(_0162_),
    .Q(\fifo.fifo[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6075_ (.CLK(clknet_leaf_20_clk),
    .D(_0163_),
    .Q(\fifo.fifo[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6076_ (.CLK(clknet_leaf_15_clk),
    .D(_0164_),
    .Q(\fifo.fifo[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6077_ (.CLK(clknet_leaf_15_clk),
    .D(_0165_),
    .Q(\fifo.fifo[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6078_ (.CLK(clknet_leaf_14_clk),
    .D(_0166_),
    .Q(\fifo.fifo[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6079_ (.CLK(clknet_leaf_12_clk),
    .D(_0167_),
    .Q(\fifo.fifo[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6080_ (.CLK(clknet_leaf_14_clk),
    .D(_0168_),
    .Q(\fifo.fifo[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6081_ (.CLK(clknet_leaf_13_clk),
    .D(_0169_),
    .Q(\fifo.fifo[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _6082_ (.CLK(clknet_leaf_11_clk),
    .D(_0170_),
    .Q(\fifo.fifo[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _6083_ (.CLK(clknet_leaf_11_clk),
    .D(_0171_),
    .Q(\fifo.fifo[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _6084_ (.CLK(clknet_leaf_11_clk),
    .D(_0172_),
    .Q(\fifo.fifo[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _6085_ (.CLK(clknet_leaf_10_clk),
    .D(_0173_),
    .Q(\fifo.fifo[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _6086_ (.CLK(clknet_leaf_1_clk),
    .D(_0174_),
    .Q(\fifo.fifo[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _6087_ (.CLK(clknet_leaf_0_clk),
    .D(_0175_),
    .Q(\fifo.fifo[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _6088_ (.CLK(clknet_leaf_69_clk),
    .D(_0176_),
    .Q(\fifo.fifo[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _6089_ (.CLK(clknet_leaf_69_clk),
    .D(_0177_),
    .Q(\fifo.fifo[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _6090_ (.CLK(clknet_leaf_2_clk),
    .D(_0178_),
    .Q(\fifo.fifo[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _6091_ (.CLK(clknet_leaf_0_clk),
    .D(_0179_),
    .Q(\fifo.fifo[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _6092_ (.CLK(clknet_leaf_3_clk),
    .D(_0180_),
    .Q(\fifo.fifo[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _6093_ (.CLK(clknet_leaf_2_clk),
    .D(_0181_),
    .Q(\fifo.fifo[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _6094_ (.CLK(clknet_leaf_68_clk),
    .D(_0182_),
    .Q(\fifo.fifo[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _6095_ (.CLK(clknet_leaf_68_clk),
    .D(_0183_),
    .Q(\fifo.fifo[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _6096_ (.CLK(clknet_leaf_66_clk),
    .D(_0184_),
    .Q(\fifo.fifo[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _6097_ (.CLK(clknet_leaf_66_clk),
    .D(_0185_),
    .Q(\fifo.fifo[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _6098_ (.CLK(clknet_leaf_60_clk),
    .D(_0186_),
    .Q(\fifo.fifo[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _6099_ (.CLK(clknet_leaf_65_clk),
    .D(_0187_),
    .Q(\fifo.fifo[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _6100_ (.CLK(clknet_leaf_64_clk),
    .D(_0188_),
    .Q(\fifo.fifo[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _6101_ (.CLK(clknet_leaf_67_clk),
    .D(_0189_),
    .Q(\fifo.fifo[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _6102_ (.CLK(clknet_leaf_61_clk),
    .D(_0190_),
    .Q(\fifo.fifo[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _6103_ (.CLK(clknet_leaf_63_clk),
    .D(_0191_),
    .Q(\fifo.fifo[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _6104_ (.CLK(clknet_leaf_53_clk),
    .D(_0192_),
    .Q(\fifo.fifo[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _6105_ (.CLK(clknet_leaf_53_clk),
    .D(_0193_),
    .Q(\fifo.fifo[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _6106_ (.CLK(clknet_leaf_52_clk),
    .D(_0194_),
    .Q(\fifo.fifo[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _6107_ (.CLK(clknet_leaf_51_clk),
    .D(_0195_),
    .Q(\fifo.fifo[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _6108_ (.CLK(clknet_leaf_46_clk),
    .D(_0196_),
    .Q(\fifo.fifo[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _6109_ (.CLK(clknet_leaf_48_clk),
    .D(_0197_),
    .Q(\fifo.fifo[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _6110_ (.CLK(clknet_leaf_48_clk),
    .D(_0198_),
    .Q(\fifo.fifo[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _6111_ (.CLK(clknet_leaf_47_clk),
    .D(_0199_),
    .Q(\fifo.fifo[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _6112_ (.CLK(clknet_leaf_45_clk),
    .D(_0200_),
    .Q(\fifo.fifo[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _6113_ (.CLK(clknet_leaf_45_clk),
    .D(_0201_),
    .Q(\fifo.fifo[2][47] ));
 sky130_fd_sc_hd__dfxtp_1 _6114_ (.CLK(clknet_leaf_49_clk),
    .D(_0202_),
    .Q(\fifo.fifo[2][48] ));
 sky130_fd_sc_hd__dfxtp_1 _6115_ (.CLK(clknet_leaf_51_clk),
    .D(_0203_),
    .Q(\fifo.fifo[2][49] ));
 sky130_fd_sc_hd__dfxtp_1 _6116_ (.CLK(clknet_leaf_54_clk),
    .D(_0204_),
    .Q(\fifo.fifo[2][50] ));
 sky130_fd_sc_hd__dfxtp_1 _6117_ (.CLK(clknet_leaf_55_clk),
    .D(_0205_),
    .Q(\fifo.fifo[2][51] ));
 sky130_fd_sc_hd__dfxtp_1 _6118_ (.CLK(clknet_leaf_58_clk),
    .D(_0206_),
    .Q(\fifo.fifo[2][52] ));
 sky130_fd_sc_hd__dfxtp_1 _6119_ (.CLK(clknet_leaf_59_clk),
    .D(_0207_),
    .Q(\fifo.fifo[2][53] ));
 sky130_fd_sc_hd__dfxtp_1 _6120_ (.CLK(clknet_leaf_61_clk),
    .D(_0208_),
    .Q(\fifo.fifo[2][54] ));
 sky130_fd_sc_hd__dfxtp_1 _6121_ (.CLK(clknet_leaf_55_clk),
    .D(_0209_),
    .Q(\fifo.fifo[2][55] ));
 sky130_fd_sc_hd__dfxtp_1 _6122_ (.CLK(clknet_leaf_26_clk),
    .D(_0210_),
    .Q(\fifo.fifo[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6123_ (.CLK(clknet_leaf_19_clk),
    .D(_0211_),
    .Q(\fifo.fifo[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6124_ (.CLK(clknet_leaf_29_clk),
    .D(_0212_),
    .Q(\fifo.fifo[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6125_ (.CLK(clknet_leaf_28_clk),
    .D(_0213_),
    .Q(\fifo.fifo[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6126_ (.CLK(clknet_leaf_28_clk),
    .D(_0214_),
    .Q(\fifo.fifo[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6127_ (.CLK(clknet_leaf_29_clk),
    .D(_0215_),
    .Q(\fifo.fifo[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6128_ (.CLK(clknet_leaf_18_clk),
    .D(_0216_),
    .Q(\fifo.fifo[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6129_ (.CLK(clknet_leaf_18_clk),
    .D(_0217_),
    .Q(\fifo.fifo[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6130_ (.CLK(clknet_leaf_17_clk),
    .D(_0218_),
    .Q(\fifo.fifo[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6131_ (.CLK(clknet_leaf_20_clk),
    .D(_0219_),
    .Q(\fifo.fifo[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6132_ (.CLK(clknet_leaf_15_clk),
    .D(_0220_),
    .Q(\fifo.fifo[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6133_ (.CLK(clknet_leaf_16_clk),
    .D(_0221_),
    .Q(\fifo.fifo[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6134_ (.CLK(clknet_leaf_14_clk),
    .D(_0222_),
    .Q(\fifo.fifo[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6135_ (.CLK(clknet_leaf_14_clk),
    .D(_0223_),
    .Q(\fifo.fifo[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6136_ (.CLK(clknet_leaf_14_clk),
    .D(_0224_),
    .Q(\fifo.fifo[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6137_ (.CLK(clknet_leaf_8_clk),
    .D(_0225_),
    .Q(\fifo.fifo[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _6138_ (.CLK(clknet_leaf_11_clk),
    .D(_0226_),
    .Q(\fifo.fifo[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _6139_ (.CLK(clknet_leaf_11_clk),
    .D(_0227_),
    .Q(\fifo.fifo[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _6140_ (.CLK(clknet_leaf_11_clk),
    .D(_0228_),
    .Q(\fifo.fifo[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _6141_ (.CLK(clknet_leaf_10_clk),
    .D(_0229_),
    .Q(\fifo.fifo[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _6142_ (.CLK(clknet_leaf_1_clk),
    .D(_0230_),
    .Q(\fifo.fifo[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _6143_ (.CLK(clknet_leaf_0_clk),
    .D(_0231_),
    .Q(\fifo.fifo[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _6144_ (.CLK(clknet_leaf_69_clk),
    .D(_0232_),
    .Q(\fifo.fifo[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _6145_ (.CLK(clknet_leaf_69_clk),
    .D(_0233_),
    .Q(\fifo.fifo[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _6146_ (.CLK(clknet_leaf_2_clk),
    .D(_0234_),
    .Q(\fifo.fifo[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _6147_ (.CLK(clknet_leaf_0_clk),
    .D(_0235_),
    .Q(\fifo.fifo[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _6148_ (.CLK(clknet_leaf_3_clk),
    .D(_0236_),
    .Q(\fifo.fifo[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _6149_ (.CLK(clknet_leaf_2_clk),
    .D(_0237_),
    .Q(\fifo.fifo[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _6150_ (.CLK(clknet_leaf_68_clk),
    .D(_0238_),
    .Q(\fifo.fifo[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _6151_ (.CLK(clknet_leaf_68_clk),
    .D(_0239_),
    .Q(\fifo.fifo[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _6152_ (.CLK(clknet_leaf_66_clk),
    .D(_0240_),
    .Q(\fifo.fifo[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _6153_ (.CLK(clknet_leaf_66_clk),
    .D(_0241_),
    .Q(\fifo.fifo[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _6154_ (.CLK(clknet_leaf_60_clk),
    .D(_0242_),
    .Q(\fifo.fifo[3][32] ));
 sky130_fd_sc_hd__dfxtp_1 _6155_ (.CLK(clknet_leaf_65_clk),
    .D(_0243_),
    .Q(\fifo.fifo[3][33] ));
 sky130_fd_sc_hd__dfxtp_1 _6156_ (.CLK(clknet_leaf_64_clk),
    .D(_0244_),
    .Q(\fifo.fifo[3][34] ));
 sky130_fd_sc_hd__dfxtp_1 _6157_ (.CLK(clknet_leaf_67_clk),
    .D(_0245_),
    .Q(\fifo.fifo[3][35] ));
 sky130_fd_sc_hd__dfxtp_1 _6158_ (.CLK(clknet_leaf_61_clk),
    .D(_0246_),
    .Q(\fifo.fifo[3][36] ));
 sky130_fd_sc_hd__dfxtp_1 _6159_ (.CLK(clknet_leaf_63_clk),
    .D(_0247_),
    .Q(\fifo.fifo[3][37] ));
 sky130_fd_sc_hd__dfxtp_1 _6160_ (.CLK(clknet_leaf_53_clk),
    .D(_0248_),
    .Q(\fifo.fifo[3][38] ));
 sky130_fd_sc_hd__dfxtp_1 _6161_ (.CLK(clknet_leaf_52_clk),
    .D(_0249_),
    .Q(\fifo.fifo[3][39] ));
 sky130_fd_sc_hd__dfxtp_1 _6162_ (.CLK(clknet_leaf_52_clk),
    .D(_0250_),
    .Q(\fifo.fifo[3][40] ));
 sky130_fd_sc_hd__dfxtp_1 _6163_ (.CLK(clknet_leaf_51_clk),
    .D(_0251_),
    .Q(\fifo.fifo[3][41] ));
 sky130_fd_sc_hd__dfxtp_1 _6164_ (.CLK(clknet_leaf_46_clk),
    .D(_0252_),
    .Q(\fifo.fifo[3][42] ));
 sky130_fd_sc_hd__dfxtp_1 _6165_ (.CLK(clknet_leaf_47_clk),
    .D(_0253_),
    .Q(\fifo.fifo[3][43] ));
 sky130_fd_sc_hd__dfxtp_1 _6166_ (.CLK(clknet_leaf_48_clk),
    .D(_0254_),
    .Q(\fifo.fifo[3][44] ));
 sky130_fd_sc_hd__dfxtp_1 _6167_ (.CLK(clknet_leaf_47_clk),
    .D(_0255_),
    .Q(\fifo.fifo[3][45] ));
 sky130_fd_sc_hd__dfxtp_1 _6168_ (.CLK(clknet_leaf_46_clk),
    .D(_0256_),
    .Q(\fifo.fifo[3][46] ));
 sky130_fd_sc_hd__dfxtp_1 _6169_ (.CLK(clknet_leaf_45_clk),
    .D(_0257_),
    .Q(\fifo.fifo[3][47] ));
 sky130_fd_sc_hd__dfxtp_1 _6170_ (.CLK(clknet_leaf_49_clk),
    .D(_0258_),
    .Q(\fifo.fifo[3][48] ));
 sky130_fd_sc_hd__dfxtp_1 _6171_ (.CLK(clknet_leaf_51_clk),
    .D(_0259_),
    .Q(\fifo.fifo[3][49] ));
 sky130_fd_sc_hd__dfxtp_1 _6172_ (.CLK(clknet_leaf_54_clk),
    .D(_0260_),
    .Q(\fifo.fifo[3][50] ));
 sky130_fd_sc_hd__dfxtp_1 _6173_ (.CLK(clknet_leaf_55_clk),
    .D(_0261_),
    .Q(\fifo.fifo[3][51] ));
 sky130_fd_sc_hd__dfxtp_1 _6174_ (.CLK(clknet_leaf_58_clk),
    .D(_0262_),
    .Q(\fifo.fifo[3][52] ));
 sky130_fd_sc_hd__dfxtp_1 _6175_ (.CLK(clknet_leaf_59_clk),
    .D(_0263_),
    .Q(\fifo.fifo[3][53] ));
 sky130_fd_sc_hd__dfxtp_1 _6176_ (.CLK(clknet_leaf_61_clk),
    .D(_0264_),
    .Q(\fifo.fifo[3][54] ));
 sky130_fd_sc_hd__dfxtp_1 _6177_ (.CLK(clknet_leaf_58_clk),
    .D(_0265_),
    .Q(\fifo.fifo[3][55] ));
 sky130_fd_sc_hd__dfxtp_1 _6178_ (.CLK(clknet_leaf_32_clk),
    .D(_0266_),
    .Q(\fifo.fifo[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6179_ (.CLK(clknet_leaf_26_clk),
    .D(_0267_),
    .Q(\fifo.fifo[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6180_ (.CLK(clknet_leaf_27_clk),
    .D(_0268_),
    .Q(\fifo.fifo[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6181_ (.CLK(clknet_leaf_29_clk),
    .D(_0269_),
    .Q(\fifo.fifo[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6182_ (.CLK(clknet_leaf_32_clk),
    .D(_0270_),
    .Q(\fifo.fifo[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6183_ (.CLK(clknet_leaf_32_clk),
    .D(_0271_),
    .Q(\fifo.fifo[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6184_ (.CLK(clknet_leaf_27_clk),
    .D(_0272_),
    .Q(\fifo.fifo[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6185_ (.CLK(clknet_leaf_18_clk),
    .D(_0273_),
    .Q(\fifo.fifo[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6186_ (.CLK(clknet_leaf_19_clk),
    .D(_0274_),
    .Q(\fifo.fifo[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6187_ (.CLK(clknet_leaf_19_clk),
    .D(_0275_),
    .Q(\fifo.fifo[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6188_ (.CLK(clknet_leaf_15_clk),
    .D(_0276_),
    .Q(\fifo.fifo[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6189_ (.CLK(clknet_leaf_17_clk),
    .D(_0277_),
    .Q(\fifo.fifo[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6190_ (.CLK(clknet_leaf_15_clk),
    .D(_0278_),
    .Q(\fifo.fifo[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6191_ (.CLK(clknet_leaf_13_clk),
    .D(_0279_),
    .Q(\fifo.fifo[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6192_ (.CLK(clknet_leaf_13_clk),
    .D(_0280_),
    .Q(\fifo.fifo[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6193_ (.CLK(clknet_leaf_20_clk),
    .D(_0281_),
    .Q(\fifo.fifo[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _6194_ (.CLK(clknet_leaf_12_clk),
    .D(_0282_),
    .Q(\fifo.fifo[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _6195_ (.CLK(clknet_leaf_8_clk),
    .D(_0283_),
    .Q(\fifo.fifo[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _6196_ (.CLK(clknet_leaf_9_clk),
    .D(_0284_),
    .Q(\fifo.fifo[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _6197_ (.CLK(clknet_leaf_9_clk),
    .D(_0285_),
    .Q(\fifo.fifo[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _6198_ (.CLK(clknet_leaf_1_clk),
    .D(_0286_),
    .Q(\fifo.fifo[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _6199_ (.CLK(clknet_leaf_1_clk),
    .D(_0287_),
    .Q(\fifo.fifo[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _6200_ (.CLK(clknet_leaf_69_clk),
    .D(_0288_),
    .Q(\fifo.fifo[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _6201_ (.CLK(clknet_leaf_69_clk),
    .D(_0289_),
    .Q(\fifo.fifo[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _6202_ (.CLK(clknet_leaf_2_clk),
    .D(_0290_),
    .Q(\fifo.fifo[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _6203_ (.CLK(clknet_leaf_0_clk),
    .D(_0291_),
    .Q(\fifo.fifo[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _6204_ (.CLK(clknet_leaf_3_clk),
    .D(_0292_),
    .Q(\fifo.fifo[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _6205_ (.CLK(clknet_leaf_3_clk),
    .D(_0293_),
    .Q(\fifo.fifo[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _6206_ (.CLK(clknet_leaf_3_clk),
    .D(_0294_),
    .Q(\fifo.fifo[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _6207_ (.CLK(clknet_leaf_3_clk),
    .D(_0295_),
    .Q(\fifo.fifo[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _6208_ (.CLK(clknet_leaf_66_clk),
    .D(_0296_),
    .Q(\fifo.fifo[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _6209_ (.CLK(clknet_leaf_64_clk),
    .D(_0297_),
    .Q(\fifo.fifo[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _6210_ (.CLK(clknet_leaf_64_clk),
    .D(_0298_),
    .Q(\fifo.fifo[4][32] ));
 sky130_fd_sc_hd__dfxtp_1 _6211_ (.CLK(clknet_leaf_64_clk),
    .D(_0299_),
    .Q(\fifo.fifo[4][33] ));
 sky130_fd_sc_hd__dfxtp_1 _6212_ (.CLK(clknet_leaf_63_clk),
    .D(_0300_),
    .Q(\fifo.fifo[4][34] ));
 sky130_fd_sc_hd__dfxtp_1 _6213_ (.CLK(clknet_leaf_65_clk),
    .D(_0301_),
    .Q(\fifo.fifo[4][35] ));
 sky130_fd_sc_hd__dfxtp_1 _6214_ (.CLK(clknet_leaf_62_clk),
    .D(_0302_),
    .Q(\fifo.fifo[4][36] ));
 sky130_fd_sc_hd__dfxtp_1 _6215_ (.CLK(clknet_leaf_62_clk),
    .D(_0303_),
    .Q(\fifo.fifo[4][37] ));
 sky130_fd_sc_hd__dfxtp_1 _6216_ (.CLK(clknet_leaf_53_clk),
    .D(_0304_),
    .Q(\fifo.fifo[4][38] ));
 sky130_fd_sc_hd__dfxtp_1 _6217_ (.CLK(clknet_leaf_53_clk),
    .D(_0305_),
    .Q(\fifo.fifo[4][39] ));
 sky130_fd_sc_hd__dfxtp_1 _6218_ (.CLK(clknet_leaf_52_clk),
    .D(_0306_),
    .Q(\fifo.fifo[4][40] ));
 sky130_fd_sc_hd__dfxtp_1 _6219_ (.CLK(clknet_leaf_52_clk),
    .D(_0307_),
    .Q(\fifo.fifo[4][41] ));
 sky130_fd_sc_hd__dfxtp_1 _6220_ (.CLK(clknet_leaf_45_clk),
    .D(_0308_),
    .Q(\fifo.fifo[4][42] ));
 sky130_fd_sc_hd__dfxtp_1 _6221_ (.CLK(clknet_leaf_47_clk),
    .D(_0309_),
    .Q(\fifo.fifo[4][43] ));
 sky130_fd_sc_hd__dfxtp_1 _6222_ (.CLK(clknet_leaf_48_clk),
    .D(_0310_),
    .Q(\fifo.fifo[4][44] ));
 sky130_fd_sc_hd__dfxtp_1 _6223_ (.CLK(clknet_leaf_47_clk),
    .D(_0311_),
    .Q(\fifo.fifo[4][45] ));
 sky130_fd_sc_hd__dfxtp_1 _6224_ (.CLK(clknet_leaf_45_clk),
    .D(_0312_),
    .Q(\fifo.fifo[4][46] ));
 sky130_fd_sc_hd__dfxtp_1 _6225_ (.CLK(clknet_leaf_45_clk),
    .D(_0313_),
    .Q(\fifo.fifo[4][47] ));
 sky130_fd_sc_hd__dfxtp_1 _6226_ (.CLK(clknet_leaf_44_clk),
    .D(_0314_),
    .Q(\fifo.fifo[4][48] ));
 sky130_fd_sc_hd__dfxtp_1 _6227_ (.CLK(clknet_leaf_50_clk),
    .D(_0315_),
    .Q(\fifo.fifo[4][49] ));
 sky130_fd_sc_hd__dfxtp_1 _6228_ (.CLK(clknet_leaf_54_clk),
    .D(_0316_),
    .Q(\fifo.fifo[4][50] ));
 sky130_fd_sc_hd__dfxtp_1 _6229_ (.CLK(clknet_leaf_56_clk),
    .D(_0317_),
    .Q(\fifo.fifo[4][51] ));
 sky130_fd_sc_hd__dfxtp_1 _6230_ (.CLK(clknet_leaf_55_clk),
    .D(_0318_),
    .Q(\fifo.fifo[4][52] ));
 sky130_fd_sc_hd__dfxtp_1 _6231_ (.CLK(clknet_leaf_58_clk),
    .D(_0319_),
    .Q(\fifo.fifo[4][53] ));
 sky130_fd_sc_hd__dfxtp_1 _6232_ (.CLK(clknet_leaf_54_clk),
    .D(_0320_),
    .Q(\fifo.fifo[4][54] ));
 sky130_fd_sc_hd__dfxtp_1 _6233_ (.CLK(clknet_leaf_58_clk),
    .D(_0321_),
    .Q(\fifo.fifo[4][55] ));
 sky130_fd_sc_hd__dfxtp_1 _6234_ (.CLK(clknet_leaf_31_clk),
    .D(_0322_),
    .Q(\fifo.fifo[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6235_ (.CLK(clknet_leaf_26_clk),
    .D(_0323_),
    .Q(\fifo.fifo[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6236_ (.CLK(clknet_leaf_26_clk),
    .D(_0324_),
    .Q(\fifo.fifo[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6237_ (.CLK(clknet_leaf_27_clk),
    .D(_0325_),
    .Q(\fifo.fifo[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6238_ (.CLK(clknet_leaf_30_clk),
    .D(_0326_),
    .Q(\fifo.fifo[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6239_ (.CLK(clknet_leaf_30_clk),
    .D(_0327_),
    .Q(\fifo.fifo[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6240_ (.CLK(clknet_leaf_18_clk),
    .D(_0328_),
    .Q(\fifo.fifo[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6241_ (.CLK(clknet_leaf_18_clk),
    .D(_0329_),
    .Q(\fifo.fifo[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6242_ (.CLK(clknet_leaf_17_clk),
    .D(_0330_),
    .Q(\fifo.fifo[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6243_ (.CLK(clknet_leaf_17_clk),
    .D(_0331_),
    .Q(\fifo.fifo[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6244_ (.CLK(clknet_leaf_15_clk),
    .D(_0332_),
    .Q(\fifo.fifo[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6245_ (.CLK(clknet_leaf_17_clk),
    .D(_0333_),
    .Q(\fifo.fifo[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6246_ (.CLK(clknet_leaf_14_clk),
    .D(_0334_),
    .Q(\fifo.fifo[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6247_ (.CLK(clknet_leaf_12_clk),
    .D(_0335_),
    .Q(\fifo.fifo[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6248_ (.CLK(clknet_leaf_13_clk),
    .D(_0336_),
    .Q(\fifo.fifo[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6249_ (.CLK(clknet_leaf_16_clk),
    .D(_0337_),
    .Q(\fifo.fifo[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _6250_ (.CLK(clknet_leaf_12_clk),
    .D(_0338_),
    .Q(\fifo.fifo[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _6251_ (.CLK(clknet_leaf_12_clk),
    .D(_0339_),
    .Q(\fifo.fifo[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _6252_ (.CLK(clknet_leaf_10_clk),
    .D(_0340_),
    .Q(\fifo.fifo[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _6253_ (.CLK(clknet_leaf_10_clk),
    .D(_0341_),
    .Q(\fifo.fifo[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _6254_ (.CLK(clknet_leaf_1_clk),
    .D(_0342_),
    .Q(\fifo.fifo[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _6255_ (.CLK(clknet_leaf_0_clk),
    .D(_0343_),
    .Q(\fifo.fifo[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _6256_ (.CLK(clknet_leaf_69_clk),
    .D(_0344_),
    .Q(\fifo.fifo[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _6257_ (.CLK(clknet_leaf_0_clk),
    .D(_0345_),
    .Q(\fifo.fifo[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _6258_ (.CLK(clknet_leaf_2_clk),
    .D(_0346_),
    .Q(\fifo.fifo[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _6259_ (.CLK(clknet_leaf_0_clk),
    .D(_0347_),
    .Q(\fifo.fifo[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _6260_ (.CLK(clknet_leaf_3_clk),
    .D(_0348_),
    .Q(\fifo.fifo[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _6261_ (.CLK(clknet_leaf_2_clk),
    .D(_0349_),
    .Q(\fifo.fifo[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _6262_ (.CLK(clknet_leaf_68_clk),
    .D(_0350_),
    .Q(\fifo.fifo[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _6263_ (.CLK(clknet_leaf_3_clk),
    .D(_0351_),
    .Q(\fifo.fifo[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _6264_ (.CLK(clknet_leaf_66_clk),
    .D(_0352_),
    .Q(\fifo.fifo[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _6265_ (.CLK(clknet_leaf_65_clk),
    .D(_0353_),
    .Q(\fifo.fifo[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _6266_ (.CLK(clknet_leaf_60_clk),
    .D(_0354_),
    .Q(\fifo.fifo[6][32] ));
 sky130_fd_sc_hd__dfxtp_1 _6267_ (.CLK(clknet_leaf_65_clk),
    .D(_0355_),
    .Q(\fifo.fifo[6][33] ));
 sky130_fd_sc_hd__dfxtp_1 _6268_ (.CLK(clknet_leaf_64_clk),
    .D(_0356_),
    .Q(\fifo.fifo[6][34] ));
 sky130_fd_sc_hd__dfxtp_1 _6269_ (.CLK(clknet_leaf_67_clk),
    .D(_0357_),
    .Q(\fifo.fifo[6][35] ));
 sky130_fd_sc_hd__dfxtp_1 _6270_ (.CLK(clknet_leaf_62_clk),
    .D(_0358_),
    .Q(\fifo.fifo[6][36] ));
 sky130_fd_sc_hd__dfxtp_1 _6271_ (.CLK(clknet_leaf_63_clk),
    .D(_0359_),
    .Q(\fifo.fifo[6][37] ));
 sky130_fd_sc_hd__dfxtp_1 _6272_ (.CLK(clknet_leaf_62_clk),
    .D(_0360_),
    .Q(\fifo.fifo[6][38] ));
 sky130_fd_sc_hd__dfxtp_1 _6273_ (.CLK(clknet_leaf_62_clk),
    .D(_0361_),
    .Q(\fifo.fifo[6][39] ));
 sky130_fd_sc_hd__dfxtp_1 _6274_ (.CLK(clknet_leaf_52_clk),
    .D(_0362_),
    .Q(\fifo.fifo[6][40] ));
 sky130_fd_sc_hd__dfxtp_1 _6275_ (.CLK(clknet_leaf_52_clk),
    .D(_0363_),
    .Q(\fifo.fifo[6][41] ));
 sky130_fd_sc_hd__dfxtp_1 _6276_ (.CLK(clknet_leaf_49_clk),
    .D(_0364_),
    .Q(\fifo.fifo[6][42] ));
 sky130_fd_sc_hd__dfxtp_1 _6277_ (.CLK(clknet_leaf_48_clk),
    .D(_0365_),
    .Q(\fifo.fifo[6][43] ));
 sky130_fd_sc_hd__dfxtp_1 _6278_ (.CLK(clknet_leaf_48_clk),
    .D(_0366_),
    .Q(\fifo.fifo[6][44] ));
 sky130_fd_sc_hd__dfxtp_1 _6279_ (.CLK(clknet_leaf_48_clk),
    .D(_0367_),
    .Q(\fifo.fifo[6][45] ));
 sky130_fd_sc_hd__dfxtp_1 _6280_ (.CLK(clknet_leaf_44_clk),
    .D(_0368_),
    .Q(\fifo.fifo[6][46] ));
 sky130_fd_sc_hd__dfxtp_1 _6281_ (.CLK(clknet_leaf_44_clk),
    .D(_0369_),
    .Q(\fifo.fifo[6][47] ));
 sky130_fd_sc_hd__dfxtp_1 _6282_ (.CLK(clknet_leaf_50_clk),
    .D(_0370_),
    .Q(\fifo.fifo[6][48] ));
 sky130_fd_sc_hd__dfxtp_1 _6283_ (.CLK(clknet_leaf_50_clk),
    .D(_0371_),
    .Q(\fifo.fifo[6][49] ));
 sky130_fd_sc_hd__dfxtp_1 _6284_ (.CLK(clknet_leaf_54_clk),
    .D(_0372_),
    .Q(\fifo.fifo[6][50] ));
 sky130_fd_sc_hd__dfxtp_1 _6285_ (.CLK(clknet_leaf_53_clk),
    .D(_0373_),
    .Q(\fifo.fifo[6][51] ));
 sky130_fd_sc_hd__dfxtp_1 _6286_ (.CLK(clknet_leaf_55_clk),
    .D(_0374_),
    .Q(\fifo.fifo[6][52] ));
 sky130_fd_sc_hd__dfxtp_1 _6287_ (.CLK(clknet_leaf_58_clk),
    .D(_0375_),
    .Q(\fifo.fifo[6][53] ));
 sky130_fd_sc_hd__dfxtp_1 _6288_ (.CLK(clknet_leaf_62_clk),
    .D(_0376_),
    .Q(\fifo.fifo[6][54] ));
 sky130_fd_sc_hd__dfxtp_1 _6289_ (.CLK(clknet_leaf_61_clk),
    .D(_0377_),
    .Q(\fifo.fifo[6][55] ));
 sky130_fd_sc_hd__dfrtp_4 _6290_ (.CLK(clknet_leaf_25_clk),
    .D(_0378_),
    .RESET_B(_0000_),
    .Q(\fifo.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6291_ (.CLK(clknet_leaf_24_clk),
    .D(_0379_),
    .RESET_B(_0001_),
    .Q(\fifo.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6292_ (.CLK(clknet_leaf_24_clk),
    .D(_0380_),
    .RESET_B(_0002_),
    .Q(\fifo.rd_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6293_ (.CLK(clknet_leaf_31_clk),
    .D(_0381_),
    .Q(\fifo.fifo[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6294_ (.CLK(clknet_leaf_19_clk),
    .D(_0382_),
    .Q(\fifo.fifo[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6295_ (.CLK(clknet_leaf_29_clk),
    .D(_0383_),
    .Q(\fifo.fifo[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6296_ (.CLK(clknet_leaf_28_clk),
    .D(_0384_),
    .Q(\fifo.fifo[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6297_ (.CLK(clknet_leaf_29_clk),
    .D(_0385_),
    .Q(\fifo.fifo[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6298_ (.CLK(clknet_leaf_30_clk),
    .D(_0386_),
    .Q(\fifo.fifo[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6299_ (.CLK(clknet_leaf_28_clk),
    .D(_0387_),
    .Q(\fifo.fifo[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6300_ (.CLK(clknet_leaf_18_clk),
    .D(_0388_),
    .Q(\fifo.fifo[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6301_ (.CLK(clknet_leaf_18_clk),
    .D(_0389_),
    .Q(\fifo.fifo[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6302_ (.CLK(clknet_leaf_20_clk),
    .D(_0390_),
    .Q(\fifo.fifo[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6303_ (.CLK(clknet_leaf_15_clk),
    .D(_0391_),
    .Q(\fifo.fifo[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6304_ (.CLK(clknet_leaf_16_clk),
    .D(_0392_),
    .Q(\fifo.fifo[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6305_ (.CLK(clknet_leaf_14_clk),
    .D(_0393_),
    .Q(\fifo.fifo[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6306_ (.CLK(clknet_leaf_12_clk),
    .D(_0394_),
    .Q(\fifo.fifo[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6307_ (.CLK(clknet_leaf_14_clk),
    .D(_0395_),
    .Q(\fifo.fifo[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6308_ (.CLK(clknet_leaf_8_clk),
    .D(_0396_),
    .Q(\fifo.fifo[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _6309_ (.CLK(clknet_leaf_11_clk),
    .D(_0397_),
    .Q(\fifo.fifo[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _6310_ (.CLK(clknet_leaf_11_clk),
    .D(_0398_),
    .Q(\fifo.fifo[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _6311_ (.CLK(clknet_leaf_11_clk),
    .D(_0399_),
    .Q(\fifo.fifo[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _6312_ (.CLK(clknet_leaf_10_clk),
    .D(_0400_),
    .Q(\fifo.fifo[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _6313_ (.CLK(clknet_leaf_1_clk),
    .D(_0401_),
    .Q(\fifo.fifo[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _6314_ (.CLK(clknet_leaf_1_clk),
    .D(_0402_),
    .Q(\fifo.fifo[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _6315_ (.CLK(clknet_leaf_69_clk),
    .D(_0403_),
    .Q(\fifo.fifo[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _6316_ (.CLK(clknet_leaf_68_clk),
    .D(_0404_),
    .Q(\fifo.fifo[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _6317_ (.CLK(clknet_leaf_2_clk),
    .D(_0405_),
    .Q(\fifo.fifo[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _6318_ (.CLK(clknet_leaf_69_clk),
    .D(_0406_),
    .Q(\fifo.fifo[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _6319_ (.CLK(clknet_leaf_3_clk),
    .D(_0407_),
    .Q(\fifo.fifo[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _6320_ (.CLK(clknet_leaf_4_clk),
    .D(_0408_),
    .Q(\fifo.fifo[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _6321_ (.CLK(clknet_leaf_68_clk),
    .D(_0409_),
    .Q(\fifo.fifo[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _6322_ (.CLK(clknet_leaf_68_clk),
    .D(_0410_),
    .Q(\fifo.fifo[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _6323_ (.CLK(clknet_leaf_66_clk),
    .D(_0411_),
    .Q(\fifo.fifo[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _6324_ (.CLK(clknet_leaf_60_clk),
    .D(_0412_),
    .Q(\fifo.fifo[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _6325_ (.CLK(clknet_leaf_61_clk),
    .D(_0413_),
    .Q(\fifo.fifo[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _6326_ (.CLK(clknet_leaf_65_clk),
    .D(_0414_),
    .Q(\fifo.fifo[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _6327_ (.CLK(clknet_leaf_63_clk),
    .D(_0415_),
    .Q(\fifo.fifo[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _6328_ (.CLK(clknet_leaf_67_clk),
    .D(_0416_),
    .Q(\fifo.fifo[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _6329_ (.CLK(clknet_leaf_62_clk),
    .D(_0417_),
    .Q(\fifo.fifo[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _6330_ (.CLK(clknet_leaf_63_clk),
    .D(_0418_),
    .Q(\fifo.fifo[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _6331_ (.CLK(clknet_leaf_53_clk),
    .D(_0419_),
    .Q(\fifo.fifo[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _6332_ (.CLK(clknet_leaf_52_clk),
    .D(_0420_),
    .Q(\fifo.fifo[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _6333_ (.CLK(clknet_leaf_52_clk),
    .D(_0421_),
    .Q(\fifo.fifo[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _6334_ (.CLK(clknet_leaf_51_clk),
    .D(_0422_),
    .Q(\fifo.fifo[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _6335_ (.CLK(clknet_leaf_47_clk),
    .D(_0423_),
    .Q(\fifo.fifo[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _6336_ (.CLK(clknet_leaf_47_clk),
    .D(_0424_),
    .Q(\fifo.fifo[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _6337_ (.CLK(clknet_leaf_48_clk),
    .D(_0425_),
    .Q(\fifo.fifo[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _6338_ (.CLK(clknet_leaf_47_clk),
    .D(_0426_),
    .Q(\fifo.fifo[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _6339_ (.CLK(clknet_leaf_46_clk),
    .D(_0427_),
    .Q(\fifo.fifo[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _6340_ (.CLK(clknet_leaf_46_clk),
    .D(_0428_),
    .Q(\fifo.fifo[1][47] ));
 sky130_fd_sc_hd__dfxtp_1 _6341_ (.CLK(clknet_leaf_49_clk),
    .D(_0429_),
    .Q(\fifo.fifo[1][48] ));
 sky130_fd_sc_hd__dfxtp_1 _6342_ (.CLK(clknet_leaf_50_clk),
    .D(_0430_),
    .Q(\fifo.fifo[1][49] ));
 sky130_fd_sc_hd__dfxtp_1 _6343_ (.CLK(clknet_leaf_54_clk),
    .D(_0431_),
    .Q(\fifo.fifo[1][50] ));
 sky130_fd_sc_hd__dfxtp_1 _6344_ (.CLK(clknet_leaf_56_clk),
    .D(_0432_),
    .Q(\fifo.fifo[1][51] ));
 sky130_fd_sc_hd__dfxtp_1 _6345_ (.CLK(clknet_leaf_57_clk),
    .D(_0433_),
    .Q(\fifo.fifo[1][52] ));
 sky130_fd_sc_hd__dfxtp_1 _6346_ (.CLK(clknet_leaf_59_clk),
    .D(_0434_),
    .Q(\fifo.fifo[1][53] ));
 sky130_fd_sc_hd__dfxtp_1 _6347_ (.CLK(clknet_leaf_61_clk),
    .D(_0435_),
    .Q(\fifo.fifo[1][54] ));
 sky130_fd_sc_hd__dfxtp_1 _6348_ (.CLK(clknet_leaf_58_clk),
    .D(_0436_),
    .Q(\fifo.fifo[1][55] ));
 sky130_fd_sc_hd__dfxtp_1 _6349_ (.CLK(clknet_leaf_25_clk),
    .D(_0437_),
    .Q(\fifo.fifo[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6350_ (.CLK(clknet_leaf_19_clk),
    .D(_0438_),
    .Q(\fifo.fifo[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6351_ (.CLK(clknet_leaf_29_clk),
    .D(_0439_),
    .Q(\fifo.fifo[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6352_ (.CLK(clknet_leaf_29_clk),
    .D(_0440_),
    .Q(\fifo.fifo[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6353_ (.CLK(clknet_leaf_29_clk),
    .D(_0441_),
    .Q(\fifo.fifo[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6354_ (.CLK(clknet_leaf_30_clk),
    .D(_0442_),
    .Q(\fifo.fifo[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6355_ (.CLK(clknet_leaf_28_clk),
    .D(_0443_),
    .Q(\fifo.fifo[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6356_ (.CLK(clknet_leaf_18_clk),
    .D(_0444_),
    .Q(\fifo.fifo[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6357_ (.CLK(clknet_leaf_18_clk),
    .D(_0445_),
    .Q(\fifo.fifo[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6358_ (.CLK(clknet_leaf_19_clk),
    .D(_0446_),
    .Q(\fifo.fifo[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6359_ (.CLK(clknet_leaf_15_clk),
    .D(_0447_),
    .Q(\fifo.fifo[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6360_ (.CLK(clknet_leaf_16_clk),
    .D(_0448_),
    .Q(\fifo.fifo[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6361_ (.CLK(clknet_leaf_13_clk),
    .D(_0449_),
    .Q(\fifo.fifo[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6362_ (.CLK(clknet_leaf_12_clk),
    .D(_0450_),
    .Q(\fifo.fifo[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6363_ (.CLK(clknet_leaf_13_clk),
    .D(_0451_),
    .Q(\fifo.fifo[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6364_ (.CLK(clknet_leaf_21_clk),
    .D(_0452_),
    .Q(\fifo.fifo[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _6365_ (.CLK(clknet_leaf_12_clk),
    .D(_0453_),
    .Q(\fifo.fifo[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _6366_ (.CLK(clknet_leaf_11_clk),
    .D(_0454_),
    .Q(\fifo.fifo[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _6367_ (.CLK(clknet_leaf_11_clk),
    .D(_0455_),
    .Q(\fifo.fifo[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _6368_ (.CLK(clknet_leaf_10_clk),
    .D(_0456_),
    .Q(\fifo.fifo[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _6369_ (.CLK(clknet_leaf_1_clk),
    .D(_0457_),
    .Q(\fifo.fifo[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _6370_ (.CLK(clknet_leaf_1_clk),
    .D(_0458_),
    .Q(\fifo.fifo[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _6371_ (.CLK(clknet_leaf_69_clk),
    .D(_0459_),
    .Q(\fifo.fifo[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _6372_ (.CLK(clknet_leaf_68_clk),
    .D(_0460_),
    .Q(\fifo.fifo[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _6373_ (.CLK(clknet_leaf_2_clk),
    .D(_0461_),
    .Q(\fifo.fifo[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _6374_ (.CLK(clknet_leaf_3_clk),
    .D(_0462_),
    .Q(\fifo.fifo[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _6375_ (.CLK(clknet_leaf_3_clk),
    .D(_0463_),
    .Q(\fifo.fifo[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _6376_ (.CLK(clknet_leaf_4_clk),
    .D(_0464_),
    .Q(\fifo.fifo[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _6377_ (.CLK(clknet_leaf_68_clk),
    .D(_0465_),
    .Q(\fifo.fifo[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _6378_ (.CLK(clknet_leaf_60_clk),
    .D(_0466_),
    .Q(\fifo.fifo[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _6379_ (.CLK(clknet_leaf_66_clk),
    .D(_0467_),
    .Q(\fifo.fifo[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _6380_ (.CLK(clknet_leaf_66_clk),
    .D(_0468_),
    .Q(\fifo.fifo[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _6381_ (.CLK(clknet_leaf_61_clk),
    .D(_0469_),
    .Q(\fifo.fifo[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _6382_ (.CLK(clknet_leaf_64_clk),
    .D(_0470_),
    .Q(\fifo.fifo[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _6383_ (.CLK(clknet_leaf_63_clk),
    .D(_0471_),
    .Q(\fifo.fifo[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _6384_ (.CLK(clknet_leaf_65_clk),
    .D(_0472_),
    .Q(\fifo.fifo[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _6385_ (.CLK(clknet_leaf_62_clk),
    .D(_0473_),
    .Q(\fifo.fifo[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _6386_ (.CLK(clknet_leaf_63_clk),
    .D(_0474_),
    .Q(\fifo.fifo[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _6387_ (.CLK(clknet_leaf_53_clk),
    .D(_0475_),
    .Q(\fifo.fifo[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _6388_ (.CLK(clknet_leaf_53_clk),
    .D(_0476_),
    .Q(\fifo.fifo[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _6389_ (.CLK(clknet_leaf_51_clk),
    .D(_0477_),
    .Q(\fifo.fifo[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _6390_ (.CLK(clknet_leaf_48_clk),
    .D(_0478_),
    .Q(\fifo.fifo[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _6391_ (.CLK(clknet_leaf_46_clk),
    .D(_0479_),
    .Q(\fifo.fifo[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _6392_ (.CLK(clknet_leaf_47_clk),
    .D(_0480_),
    .Q(\fifo.fifo[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _6393_ (.CLK(clknet_leaf_48_clk),
    .D(_0481_),
    .Q(\fifo.fifo[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _6394_ (.CLK(clknet_leaf_47_clk),
    .D(_0482_),
    .Q(\fifo.fifo[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _6395_ (.CLK(clknet_leaf_46_clk),
    .D(_0483_),
    .Q(\fifo.fifo[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _6396_ (.CLK(clknet_leaf_46_clk),
    .D(_0484_),
    .Q(\fifo.fifo[0][47] ));
 sky130_fd_sc_hd__dfxtp_1 _6397_ (.CLK(clknet_leaf_49_clk),
    .D(_0485_),
    .Q(\fifo.fifo[0][48] ));
 sky130_fd_sc_hd__dfxtp_1 _6398_ (.CLK(clknet_leaf_50_clk),
    .D(_0486_),
    .Q(\fifo.fifo[0][49] ));
 sky130_fd_sc_hd__dfxtp_1 _6399_ (.CLK(clknet_leaf_55_clk),
    .D(_0487_),
    .Q(\fifo.fifo[0][50] ));
 sky130_fd_sc_hd__dfxtp_1 _6400_ (.CLK(clknet_leaf_56_clk),
    .D(_0488_),
    .Q(\fifo.fifo[0][51] ));
 sky130_fd_sc_hd__dfxtp_1 _6401_ (.CLK(clknet_leaf_57_clk),
    .D(_0489_),
    .Q(\fifo.fifo[0][52] ));
 sky130_fd_sc_hd__dfxtp_1 _6402_ (.CLK(clknet_leaf_59_clk),
    .D(_0490_),
    .Q(\fifo.fifo[0][53] ));
 sky130_fd_sc_hd__dfxtp_1 _6403_ (.CLK(clknet_leaf_54_clk),
    .D(_0491_),
    .Q(\fifo.fifo[0][54] ));
 sky130_fd_sc_hd__dfxtp_1 _6404_ (.CLK(clknet_leaf_55_clk),
    .D(_0492_),
    .Q(\fifo.fifo[0][55] ));
 sky130_fd_sc_hd__dfxtp_1 _6405_ (.CLK(clknet_leaf_31_clk),
    .D(_0493_),
    .Q(\fifo.fifo[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6406_ (.CLK(clknet_leaf_26_clk),
    .D(_0494_),
    .Q(\fifo.fifo[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6407_ (.CLK(clknet_leaf_27_clk),
    .D(_0495_),
    .Q(\fifo.fifo[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6408_ (.CLK(clknet_leaf_28_clk),
    .D(_0496_),
    .Q(\fifo.fifo[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6409_ (.CLK(clknet_leaf_29_clk),
    .D(_0497_),
    .Q(\fifo.fifo[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6410_ (.CLK(clknet_leaf_30_clk),
    .D(_0498_),
    .Q(\fifo.fifo[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6411_ (.CLK(clknet_leaf_18_clk),
    .D(_0499_),
    .Q(\fifo.fifo[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6412_ (.CLK(clknet_leaf_18_clk),
    .D(_0500_),
    .Q(\fifo.fifo[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6413_ (.CLK(clknet_leaf_17_clk),
    .D(_0501_),
    .Q(\fifo.fifo[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _6414_ (.CLK(clknet_leaf_17_clk),
    .D(_0502_),
    .Q(\fifo.fifo[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _6415_ (.CLK(clknet_leaf_15_clk),
    .D(_0503_),
    .Q(\fifo.fifo[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _6416_ (.CLK(clknet_leaf_17_clk),
    .D(_0504_),
    .Q(\fifo.fifo[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _6417_ (.CLK(clknet_leaf_14_clk),
    .D(_0505_),
    .Q(\fifo.fifo[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _6418_ (.CLK(clknet_leaf_12_clk),
    .D(_0506_),
    .Q(\fifo.fifo[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _6419_ (.CLK(clknet_leaf_13_clk),
    .D(_0507_),
    .Q(\fifo.fifo[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _6420_ (.CLK(clknet_leaf_16_clk),
    .D(_0508_),
    .Q(\fifo.fifo[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _6421_ (.CLK(clknet_leaf_12_clk),
    .D(_0509_),
    .Q(\fifo.fifo[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _6422_ (.CLK(clknet_leaf_12_clk),
    .D(_0510_),
    .Q(\fifo.fifo[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _6423_ (.CLK(clknet_leaf_10_clk),
    .D(_0511_),
    .Q(\fifo.fifo[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _6424_ (.CLK(clknet_leaf_10_clk),
    .D(_0512_),
    .Q(\fifo.fifo[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _6425_ (.CLK(clknet_leaf_1_clk),
    .D(_0513_),
    .Q(\fifo.fifo[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _6426_ (.CLK(clknet_leaf_0_clk),
    .D(_0514_),
    .Q(\fifo.fifo[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _6427_ (.CLK(clknet_leaf_69_clk),
    .D(_0515_),
    .Q(\fifo.fifo[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _6428_ (.CLK(clknet_leaf_0_clk),
    .D(_0516_),
    .Q(\fifo.fifo[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _6429_ (.CLK(clknet_leaf_2_clk),
    .D(_0517_),
    .Q(\fifo.fifo[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _6430_ (.CLK(clknet_leaf_0_clk),
    .D(_0518_),
    .Q(\fifo.fifo[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _6431_ (.CLK(clknet_leaf_3_clk),
    .D(_0519_),
    .Q(\fifo.fifo[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _6432_ (.CLK(clknet_leaf_2_clk),
    .D(_0520_),
    .Q(\fifo.fifo[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _6433_ (.CLK(clknet_leaf_68_clk),
    .D(_0521_),
    .Q(\fifo.fifo[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _6434_ (.CLK(clknet_leaf_3_clk),
    .D(_0522_),
    .Q(\fifo.fifo[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _6435_ (.CLK(clknet_leaf_66_clk),
    .D(_0523_),
    .Q(\fifo.fifo[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _6436_ (.CLK(clknet_leaf_65_clk),
    .D(_0524_),
    .Q(\fifo.fifo[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _6437_ (.CLK(clknet_leaf_60_clk),
    .D(_0525_),
    .Q(\fifo.fifo[7][32] ));
 sky130_fd_sc_hd__dfxtp_1 _6438_ (.CLK(clknet_leaf_65_clk),
    .D(_0526_),
    .Q(\fifo.fifo[7][33] ));
 sky130_fd_sc_hd__dfxtp_1 _6439_ (.CLK(clknet_leaf_64_clk),
    .D(_0527_),
    .Q(\fifo.fifo[7][34] ));
 sky130_fd_sc_hd__dfxtp_1 _6440_ (.CLK(clknet_leaf_67_clk),
    .D(_0528_),
    .Q(\fifo.fifo[7][35] ));
 sky130_fd_sc_hd__dfxtp_1 _6441_ (.CLK(clknet_leaf_62_clk),
    .D(_0529_),
    .Q(\fifo.fifo[7][36] ));
 sky130_fd_sc_hd__dfxtp_1 _6442_ (.CLK(clknet_leaf_63_clk),
    .D(_0530_),
    .Q(\fifo.fifo[7][37] ));
 sky130_fd_sc_hd__dfxtp_1 _6443_ (.CLK(clknet_leaf_53_clk),
    .D(_0531_),
    .Q(\fifo.fifo[7][38] ));
 sky130_fd_sc_hd__dfxtp_1 _6444_ (.CLK(clknet_leaf_62_clk),
    .D(_0532_),
    .Q(\fifo.fifo[7][39] ));
 sky130_fd_sc_hd__dfxtp_1 _6445_ (.CLK(clknet_leaf_52_clk),
    .D(_0533_),
    .Q(\fifo.fifo[7][40] ));
 sky130_fd_sc_hd__dfxtp_1 _6446_ (.CLK(clknet_leaf_51_clk),
    .D(_0534_),
    .Q(\fifo.fifo[7][41] ));
 sky130_fd_sc_hd__dfxtp_1 _6447_ (.CLK(clknet_leaf_49_clk),
    .D(_0535_),
    .Q(\fifo.fifo[7][42] ));
 sky130_fd_sc_hd__dfxtp_1 _6448_ (.CLK(clknet_leaf_47_clk),
    .D(_0536_),
    .Q(\fifo.fifo[7][43] ));
 sky130_fd_sc_hd__dfxtp_1 _6449_ (.CLK(clknet_leaf_48_clk),
    .D(_0537_),
    .Q(\fifo.fifo[7][44] ));
 sky130_fd_sc_hd__dfxtp_1 _6450_ (.CLK(clknet_leaf_48_clk),
    .D(_0538_),
    .Q(\fifo.fifo[7][45] ));
 sky130_fd_sc_hd__dfxtp_1 _6451_ (.CLK(clknet_leaf_44_clk),
    .D(_0539_),
    .Q(\fifo.fifo[7][46] ));
 sky130_fd_sc_hd__dfxtp_1 _6452_ (.CLK(clknet_leaf_44_clk),
    .D(_0540_),
    .Q(\fifo.fifo[7][47] ));
 sky130_fd_sc_hd__dfxtp_1 _6453_ (.CLK(clknet_leaf_49_clk),
    .D(_0541_),
    .Q(\fifo.fifo[7][48] ));
 sky130_fd_sc_hd__dfxtp_1 _6454_ (.CLK(clknet_leaf_56_clk),
    .D(_0542_),
    .Q(\fifo.fifo[7][49] ));
 sky130_fd_sc_hd__dfxtp_1 _6455_ (.CLK(clknet_leaf_54_clk),
    .D(_0543_),
    .Q(\fifo.fifo[7][50] ));
 sky130_fd_sc_hd__dfxtp_1 _6456_ (.CLK(clknet_leaf_54_clk),
    .D(_0544_),
    .Q(\fifo.fifo[7][51] ));
 sky130_fd_sc_hd__dfxtp_1 _6457_ (.CLK(clknet_leaf_55_clk),
    .D(_0545_),
    .Q(\fifo.fifo[7][52] ));
 sky130_fd_sc_hd__dfxtp_1 _6458_ (.CLK(clknet_leaf_59_clk),
    .D(_0546_),
    .Q(\fifo.fifo[7][53] ));
 sky130_fd_sc_hd__dfxtp_1 _6459_ (.CLK(clknet_leaf_61_clk),
    .D(_0547_),
    .Q(\fifo.fifo[7][54] ));
 sky130_fd_sc_hd__dfxtp_1 _6460_ (.CLK(clknet_leaf_58_clk),
    .D(_0548_),
    .Q(\fifo.fifo[7][55] ));
 sky130_fd_sc_hd__dfrtp_4 _6461_ (.CLK(clknet_leaf_31_clk),
    .D(_0549_),
    .RESET_B(_0003_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_4 _6462_ (.CLK(clknet_leaf_25_clk),
    .D(_0550_),
    .RESET_B(_0004_),
    .Q(net135));
 sky130_fd_sc_hd__dfrtp_4 _6463_ (.CLK(clknet_leaf_33_clk),
    .D(_0551_),
    .RESET_B(_0005_),
    .Q(net146));
 sky130_fd_sc_hd__dfrtp_4 _6464_ (.CLK(clknet_leaf_26_clk),
    .D(_0552_),
    .RESET_B(_0006_),
    .Q(net157));
 sky130_fd_sc_hd__dfrtp_4 _6465_ (.CLK(clknet_leaf_33_clk),
    .D(_0553_),
    .RESET_B(_0007_),
    .Q(net168));
 sky130_fd_sc_hd__dfrtp_2 _6466_ (.CLK(clknet_leaf_32_clk),
    .D(_0554_),
    .RESET_B(_0008_),
    .Q(net179));
 sky130_fd_sc_hd__dfrtp_4 _6467_ (.CLK(clknet_leaf_24_clk),
    .D(_0555_),
    .RESET_B(_0009_),
    .Q(net184));
 sky130_fd_sc_hd__dfrtp_4 _6468_ (.CLK(clknet_leaf_32_clk),
    .D(_0556_),
    .RESET_B(_0010_),
    .Q(net185));
 sky130_fd_sc_hd__dfrtp_4 _6469_ (.CLK(clknet_leaf_19_clk),
    .D(_0557_),
    .RESET_B(_0011_),
    .Q(net186));
 sky130_fd_sc_hd__dfrtp_2 _6470_ (.CLK(clknet_leaf_32_clk),
    .D(_0558_),
    .RESET_B(_0012_),
    .Q(net187));
 sky130_fd_sc_hd__dfrtp_4 _6471_ (.CLK(clknet_leaf_32_clk),
    .D(_0559_),
    .RESET_B(_0013_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_4 _6472_ (.CLK(clknet_leaf_32_clk),
    .D(_0560_),
    .RESET_B(_0014_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_4 _6473_ (.CLK(clknet_leaf_20_clk),
    .D(_0561_),
    .RESET_B(_0015_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_4 _6474_ (.CLK(clknet_leaf_21_clk),
    .D(_0562_),
    .RESET_B(_0016_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_4 _6475_ (.CLK(clknet_leaf_20_clk),
    .D(_0563_),
    .RESET_B(_0017_),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_4 _6476_ (.CLK(clknet_leaf_20_clk),
    .D(_0564_),
    .RESET_B(_0018_),
    .Q(net130));
 sky130_fd_sc_hd__dfrtp_2 _6477_ (.CLK(clknet_leaf_7_clk),
    .D(_0565_),
    .RESET_B(_0019_),
    .Q(net131));
 sky130_fd_sc_hd__dfrtp_4 _6478_ (.CLK(clknet_leaf_8_clk),
    .D(_0566_),
    .RESET_B(_0020_),
    .Q(net132));
 sky130_fd_sc_hd__dfrtp_4 _6479_ (.CLK(clknet_leaf_8_clk),
    .D(_0567_),
    .RESET_B(_0021_),
    .Q(net133));
 sky130_fd_sc_hd__dfrtp_2 _6480_ (.CLK(clknet_leaf_12_clk),
    .D(net193),
    .RESET_B(_0022_),
    .Q(net134));
 sky130_fd_sc_hd__dfrtp_4 _6481_ (.CLK(clknet_leaf_9_clk),
    .D(_0569_),
    .RESET_B(_0023_),
    .Q(net136));
 sky130_fd_sc_hd__dfrtp_2 _6482_ (.CLK(clknet_leaf_9_clk),
    .D(_0570_),
    .RESET_B(_0024_),
    .Q(net137));
 sky130_fd_sc_hd__dfrtp_2 _6483_ (.CLK(clknet_leaf_9_clk),
    .D(_0571_),
    .RESET_B(_0025_),
    .Q(net138));
 sky130_fd_sc_hd__dfrtp_4 _6484_ (.CLK(clknet_leaf_6_clk),
    .D(_0572_),
    .RESET_B(_0026_),
    .Q(net139));
 sky130_fd_sc_hd__dfrtp_2 _6485_ (.CLK(clknet_leaf_21_clk),
    .D(net688),
    .RESET_B(_0027_),
    .Q(net140));
 sky130_fd_sc_hd__dfrtp_4 _6486_ (.CLK(clknet_leaf_9_clk),
    .D(_0574_),
    .RESET_B(_0028_),
    .Q(net141));
 sky130_fd_sc_hd__dfrtp_4 _6487_ (.CLK(clknet_leaf_21_clk),
    .D(_0575_),
    .RESET_B(_0029_),
    .Q(net142));
 sky130_fd_sc_hd__dfrtp_4 _6488_ (.CLK(clknet_leaf_59_clk),
    .D(_0576_),
    .RESET_B(_0030_),
    .Q(net143));
 sky130_fd_sc_hd__dfrtp_2 _6489_ (.CLK(clknet_leaf_6_clk),
    .D(_0577_),
    .RESET_B(_0031_),
    .Q(net144));
 sky130_fd_sc_hd__dfrtp_4 _6490_ (.CLK(clknet_leaf_7_clk),
    .D(_0578_),
    .RESET_B(_0032_),
    .Q(net145));
 sky130_fd_sc_hd__dfrtp_4 _6491_ (.CLK(clknet_leaf_60_clk),
    .D(_0579_),
    .RESET_B(_0033_),
    .Q(net147));
 sky130_fd_sc_hd__dfrtp_2 _6492_ (.CLK(clknet_leaf_59_clk),
    .D(_0580_),
    .RESET_B(_0034_),
    .Q(net148));
 sky130_fd_sc_hd__dfrtp_4 _6493_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0581_),
    .RESET_B(_0035_),
    .Q(net149));
 sky130_fd_sc_hd__dfrtp_4 _6494_ (.CLK(clknet_leaf_59_clk),
    .D(_0582_),
    .RESET_B(_0036_),
    .Q(net150));
 sky130_fd_sc_hd__dfrtp_2 _6495_ (.CLK(clknet_leaf_59_clk),
    .D(_0583_),
    .RESET_B(_0037_),
    .Q(net151));
 sky130_fd_sc_hd__dfrtp_4 _6496_ (.CLK(clknet_leaf_42_clk),
    .D(_0584_),
    .RESET_B(_0038_),
    .Q(net152));
 sky130_fd_sc_hd__dfrtp_4 _6497_ (.CLK(clknet_leaf_42_clk),
    .D(_0585_),
    .RESET_B(_0039_),
    .Q(net153));
 sky130_fd_sc_hd__dfrtp_2 _6498_ (.CLK(clknet_leaf_43_clk),
    .D(_0586_),
    .RESET_B(_0040_),
    .Q(net154));
 sky130_fd_sc_hd__dfrtp_2 _6499_ (.CLK(clknet_leaf_34_clk),
    .D(_0587_),
    .RESET_B(_0041_),
    .Q(net155));
 sky130_fd_sc_hd__dfrtp_4 _6500_ (.CLK(clknet_leaf_34_clk),
    .D(_0588_),
    .RESET_B(_0042_),
    .Q(net156));
 sky130_fd_sc_hd__dfrtp_4 _6501_ (.CLK(clknet_leaf_34_clk),
    .D(_0589_),
    .RESET_B(_0043_),
    .Q(net158));
 sky130_fd_sc_hd__dfrtp_4 _6502_ (.CLK(clknet_leaf_42_clk),
    .D(_0590_),
    .RESET_B(_0044_),
    .Q(net159));
 sky130_fd_sc_hd__dfrtp_4 _6503_ (.CLK(clknet_leaf_33_clk),
    .D(_0591_),
    .RESET_B(_0045_),
    .Q(net160));
 sky130_fd_sc_hd__dfrtp_4 _6504_ (.CLK(clknet_leaf_42_clk),
    .D(_0592_),
    .RESET_B(_0046_),
    .Q(net161));
 sky130_fd_sc_hd__dfrtp_4 _6505_ (.CLK(clknet_leaf_43_clk),
    .D(_0593_),
    .RESET_B(_0047_),
    .Q(net162));
 sky130_fd_sc_hd__dfrtp_4 _6506_ (.CLK(clknet_leaf_41_clk),
    .D(_0594_),
    .RESET_B(_0048_),
    .Q(net163));
 sky130_fd_sc_hd__dfrtp_4 _6507_ (.CLK(clknet_leaf_41_clk),
    .D(_0595_),
    .RESET_B(_0049_),
    .Q(net164));
 sky130_fd_sc_hd__dfrtp_2 _6508_ (.CLK(clknet_leaf_41_clk),
    .D(_0596_),
    .RESET_B(_0050_),
    .Q(net165));
 sky130_fd_sc_hd__dfrtp_4 _6509_ (.CLK(clknet_leaf_38_clk),
    .D(_0597_),
    .RESET_B(_0051_),
    .Q(net166));
 sky130_fd_sc_hd__dfrtp_2 _6510_ (.CLK(clknet_leaf_35_clk),
    .D(_0598_),
    .RESET_B(_0052_),
    .Q(net167));
 sky130_fd_sc_hd__dfrtp_4 _6511_ (.CLK(clknet_leaf_35_clk),
    .D(_0599_),
    .RESET_B(_0053_),
    .Q(net169));
 sky130_fd_sc_hd__dfrtp_4 _6512_ (.CLK(clknet_leaf_35_clk),
    .D(_0600_),
    .RESET_B(_0054_),
    .Q(net170));
 sky130_fd_sc_hd__dfrtp_2 _6513_ (.CLK(clknet_leaf_38_clk),
    .D(_0601_),
    .RESET_B(_0055_),
    .Q(net171));
 sky130_fd_sc_hd__dfrtp_4 _6514_ (.CLK(clknet_leaf_38_clk),
    .D(_0602_),
    .RESET_B(_0056_),
    .Q(net172));
 sky130_fd_sc_hd__dfrtp_4 _6515_ (.CLK(clknet_leaf_25_clk),
    .D(_0603_),
    .RESET_B(_0057_),
    .Q(net173));
 sky130_fd_sc_hd__dfrtp_2 _6516_ (.CLK(clknet_leaf_41_clk),
    .D(_0604_),
    .RESET_B(_0058_),
    .Q(net174));
 sky130_fd_sc_hd__dfrtp_4 _6517_ (.CLK(clknet_leaf_41_clk),
    .D(_0605_),
    .RESET_B(_0059_),
    .Q(net175));
 sky130_fd_sc_hd__dfrtp_4 _6518_ (.CLK(clknet_leaf_34_clk),
    .D(_0606_),
    .RESET_B(_0060_),
    .Q(net176));
 sky130_fd_sc_hd__dfrtp_2 _6519_ (.CLK(clknet_leaf_41_clk),
    .D(_0607_),
    .RESET_B(_0061_),
    .Q(net177));
 sky130_fd_sc_hd__dfrtp_4 _6520_ (.CLK(clknet_leaf_34_clk),
    .D(_0608_),
    .RESET_B(_0062_),
    .Q(net178));
 sky130_fd_sc_hd__dfrtp_4 _6521_ (.CLK(clknet_leaf_34_clk),
    .D(_0609_),
    .RESET_B(_0063_),
    .Q(net180));
 sky130_fd_sc_hd__dfrtp_4 _6522_ (.CLK(clknet_leaf_34_clk),
    .D(_0610_),
    .RESET_B(_0064_),
    .Q(net181));
 sky130_fd_sc_hd__dfrtp_4 _6523_ (.CLK(clknet_leaf_42_clk),
    .D(_0611_),
    .RESET_B(_0065_),
    .Q(net182));
 sky130_fd_sc_hd__dfrtp_4 _6524_ (.CLK(clknet_leaf_41_clk),
    .D(_0612_),
    .RESET_B(_0066_),
    .Q(net183));
 sky130_fd_sc_hd__dfstp_1 _6525_ (.CLK(clknet_leaf_37_clk),
    .D(_0613_),
    .SET_B(_0067_),
    .Q(\fifo.fifo_empty ));
 sky130_fd_sc_hd__dfrtp_1 _6526_ (.CLK(clknet_leaf_38_clk),
    .D(_0614_),
    .RESET_B(_0068_),
    .Q(\fifo.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6527_ (.CLK(clknet_leaf_57_clk),
    .D(_0615_),
    .RESET_B(_0069_),
    .Q(\fifo.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6528_ (.CLK(clknet_leaf_57_clk),
    .D(_0616_),
    .RESET_B(_0070_),
    .Q(\fifo.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6529_ (.CLK(clknet_leaf_37_clk),
    .D(_0617_),
    .RESET_B(_0071_),
    .Q(net188));
 sky130_fd_sc_hd__dfrtp_1 _6530_ (.CLK(clknet_leaf_37_clk),
    .D(_0618_),
    .RESET_B(_0072_),
    .Q(\counter_inst.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6531_ (.CLK(clknet_leaf_25_clk),
    .D(_0619_),
    .RESET_B(_0073_),
    .Q(\counter_inst.count[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6532_ (.CLK(clknet_leaf_25_clk),
    .D(_0620_),
    .RESET_B(_0074_),
    .Q(\counter_inst.count[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6533_ (.CLK(clknet_leaf_25_clk),
    .D(_0621_),
    .RESET_B(_0075_),
    .Q(\counter_inst.count[3] ));
 sky130_fd_sc_hd__dfstp_1 _6534_ (.CLK(clknet_leaf_25_clk),
    .D(_0622_),
    .SET_B(_0076_),
    .Q(\counter_inst.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6535_ (.CLK(clknet_leaf_33_clk),
    .D(\u0.E[1] ),
    .Q(\L[32] ));
 sky130_fd_sc_hd__dfxtp_1 _6536_ (.CLK(clknet_leaf_35_clk),
    .D(\u0.E[46] ),
    .Q(\L[31] ));
 sky130_fd_sc_hd__dfxtp_1 _6537_ (.CLK(clknet_leaf_34_clk),
    .D(\u0.E[45] ),
    .Q(\L[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6538_ (.CLK(clknet_leaf_5_clk),
    .D(\u0.E[42] ),
    .Q(\L[29] ));
 sky130_fd_sc_hd__dfxtp_1 _6539_ (.CLK(clknet_leaf_21_clk),
    .D(\u0.E[41] ),
    .Q(\L[28] ));
 sky130_fd_sc_hd__dfxtp_1 _6540_ (.CLK(clknet_leaf_7_clk),
    .D(\u0.E[40] ),
    .Q(\L[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6541_ (.CLK(clknet_leaf_22_clk),
    .D(\u0.E[39] ),
    .Q(\L[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6542_ (.CLK(clknet_leaf_20_clk),
    .D(\u0.E[36] ),
    .Q(\L[25] ));
 sky130_fd_sc_hd__dfxtp_1 _6543_ (.CLK(clknet_leaf_35_clk),
    .D(\u0.E[35] ),
    .Q(\L[24] ));
 sky130_fd_sc_hd__dfxtp_1 _6544_ (.CLK(clknet_leaf_36_clk),
    .D(\u0.E[34] ),
    .Q(\L[23] ));
 sky130_fd_sc_hd__dfxtp_1 _6545_ (.CLK(clknet_leaf_33_clk),
    .D(\u0.E[33] ),
    .Q(\L[22] ));
 sky130_fd_sc_hd__dfxtp_1 _6546_ (.CLK(clknet_leaf_7_clk),
    .D(\u0.E[30] ),
    .Q(\L[21] ));
 sky130_fd_sc_hd__dfxtp_1 _6547_ (.CLK(clknet_leaf_22_clk),
    .D(\u0.E[29] ),
    .Q(\L[20] ));
 sky130_fd_sc_hd__dfxtp_1 _6548_ (.CLK(clknet_leaf_7_clk),
    .D(\u0.E[28] ),
    .Q(\L[19] ));
 sky130_fd_sc_hd__dfxtp_1 _6549_ (.CLK(clknet_leaf_19_clk),
    .D(\u0.E[27] ),
    .Q(\L[18] ));
 sky130_fd_sc_hd__dfxtp_1 _6550_ (.CLK(clknet_leaf_31_clk),
    .D(\u0.E[24] ),
    .Q(\L[17] ));
 sky130_fd_sc_hd__dfxtp_1 _6551_ (.CLK(clknet_leaf_41_clk),
    .D(\u0.E[23] ),
    .Q(\L[16] ));
 sky130_fd_sc_hd__dfxtp_1 _6552_ (.CLK(clknet_leaf_37_clk),
    .D(\u0.E[22] ),
    .Q(\L[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6553_ (.CLK(clknet_leaf_38_clk),
    .D(\u0.E[21] ),
    .Q(\L[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6554_ (.CLK(clknet_leaf_36_clk),
    .D(\u0.E[18] ),
    .Q(\L[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6555_ (.CLK(clknet_leaf_21_clk),
    .D(\u0.E[17] ),
    .Q(\L[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6556_ (.CLK(clknet_leaf_6_clk),
    .D(\u0.E[16] ),
    .Q(\L[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6557_ (.CLK(clknet_leaf_21_clk),
    .D(\u0.E[15] ),
    .Q(\L[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6558_ (.CLK(clknet_leaf_32_clk),
    .D(\u0.E[12] ),
    .Q(\L[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6559_ (.CLK(clknet_leaf_39_clk),
    .D(\u0.E[11] ),
    .Q(\L[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6560_ (.CLK(clknet_leaf_25_clk),
    .D(\u0.E[10] ),
    .Q(\L[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6561_ (.CLK(clknet_leaf_39_clk),
    .D(\u0.E[9] ),
    .Q(\L[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6562_ (.CLK(clknet_leaf_34_clk),
    .D(\u0.E[6] ),
    .Q(\L[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6563_ (.CLK(clknet_leaf_7_clk),
    .D(\u0.E[5] ),
    .Q(\L[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6564_ (.CLK(clknet_leaf_6_clk),
    .D(\u0.E[4] ),
    .Q(\L[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6565_ (.CLK(clknet_leaf_21_clk),
    .D(\u0.E[3] ),
    .Q(\L[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6566_ (.CLK(clknet_leaf_24_clk),
    .D(\u0.E[2] ),
    .Q(\L[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6567_ (.CLK(clknet_leaf_35_clk),
    .D(\FP[32] ),
    .Q(\R[32] ));
 sky130_fd_sc_hd__dfxtp_1 _6568_ (.CLK(clknet_leaf_39_clk),
    .D(\FP[31] ),
    .Q(\R[31] ));
 sky130_fd_sc_hd__dfxtp_1 _6569_ (.CLK(clknet_leaf_35_clk),
    .D(\FP[30] ),
    .Q(\R[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6570_ (.CLK(clknet_leaf_5_clk),
    .D(\FP[29] ),
    .Q(\R[29] ));
 sky130_fd_sc_hd__dfxtp_1 _6571_ (.CLK(clknet_leaf_21_clk),
    .D(\FP[28] ),
    .Q(\R[28] ));
 sky130_fd_sc_hd__dfxtp_1 _6572_ (.CLK(clknet_leaf_7_clk),
    .D(\FP[27] ),
    .Q(\R[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6573_ (.CLK(clknet_leaf_19_clk),
    .D(\FP[26] ),
    .Q(\R[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6574_ (.CLK(clknet_leaf_19_clk),
    .D(\FP[25] ),
    .Q(\R[25] ));
 sky130_fd_sc_hd__dfxtp_1 _6575_ (.CLK(clknet_3_3__leaf_clk),
    .D(\FP[24] ),
    .Q(\R[24] ));
 sky130_fd_sc_hd__dfxtp_1 _6576_ (.CLK(clknet_leaf_36_clk),
    .D(\FP[23] ),
    .Q(\R[23] ));
 sky130_fd_sc_hd__dfxtp_1 _6577_ (.CLK(clknet_leaf_25_clk),
    .D(\FP[22] ),
    .Q(\R[22] ));
 sky130_fd_sc_hd__dfxtp_1 _6578_ (.CLK(clknet_leaf_5_clk),
    .D(\FP[21] ),
    .Q(\R[21] ));
 sky130_fd_sc_hd__dfxtp_1 _6579_ (.CLK(clknet_leaf_21_clk),
    .D(\FP[20] ),
    .Q(\R[20] ));
 sky130_fd_sc_hd__dfxtp_1 _6580_ (.CLK(clknet_leaf_7_clk),
    .D(\FP[19] ),
    .Q(\R[19] ));
 sky130_fd_sc_hd__dfxtp_1 _6581_ (.CLK(clknet_leaf_19_clk),
    .D(\FP[18] ),
    .Q(\R[18] ));
 sky130_fd_sc_hd__dfxtp_1 _6582_ (.CLK(clknet_leaf_32_clk),
    .D(\FP[17] ),
    .Q(\R[17] ));
 sky130_fd_sc_hd__dfxtp_1 _6583_ (.CLK(clknet_leaf_35_clk),
    .D(\FP[16] ),
    .Q(\R[16] ));
 sky130_fd_sc_hd__dfxtp_1 _6584_ (.CLK(clknet_leaf_37_clk),
    .D(\FP[15] ),
    .Q(\R[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6585_ (.CLK(clknet_leaf_43_clk),
    .D(\FP[14] ),
    .Q(\R[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6586_ (.CLK(clknet_leaf_43_clk),
    .D(\FP[13] ),
    .Q(\R[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6587_ (.CLK(clknet_leaf_21_clk),
    .D(\FP[12] ),
    .Q(\R[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6588_ (.CLK(clknet_leaf_6_clk),
    .D(\FP[11] ),
    .Q(\R[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6589_ (.CLK(clknet_leaf_21_clk),
    .D(\FP[10] ),
    .Q(\R[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6590_ (.CLK(clknet_leaf_33_clk),
    .D(\FP[9] ),
    .Q(\R[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6591_ (.CLK(clknet_leaf_41_clk),
    .D(\FP[8] ),
    .Q(\R[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6592_ (.CLK(clknet_leaf_25_clk),
    .D(\FP[7] ),
    .Q(\R[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6593_ (.CLK(clknet_leaf_41_clk),
    .D(\FP[6] ),
    .Q(\R[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6594_ (.CLK(clknet_leaf_34_clk),
    .D(\FP[5] ),
    .Q(\R[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6595_ (.CLK(clknet_leaf_4_clk),
    .D(\FP[4] ),
    .Q(\R[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6596_ (.CLK(clknet_leaf_6_clk),
    .D(\FP[3] ),
    .Q(\R[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6597_ (.CLK(clknet_leaf_21_clk),
    .D(\FP[2] ),
    .Q(\R[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6598_ (.CLK(clknet_leaf_24_clk),
    .D(\FP[1] ),
    .Q(\R[1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\R[24] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\fifo.fifo[1][41] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\fifo.fifo[5][31] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\fifo.fifo[1][19] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\fifo.fifo[0][12] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\fifo.fifo[4][45] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\fifo.fifo[6][4] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\fifo.fifo[1][49] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\fifo.fifo[0][22] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\fifo.fifo[2][44] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\fifo.fifo[1][23] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\fifo.fifo[0][18] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\fifo.fifo[1][11] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\fifo.fifo[6][22] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\fifo.fifo[2][45] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\fifo.fifo[1][2] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\fifo.fifo[0][1] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\fifo.fifo[4][1] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\fifo.fifo[5][24] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\fifo.fifo[2][50] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\fifo.fifo[2][51] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\fifo.fifo[5][32] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\fifo.fifo[5][4] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\fifo.fifo[0][40] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\fifo.fifo[7][0] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\fifo.fifo[3][51] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\fifo.fifo[1][54] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\fifo.fifo[1][36] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\fifo.fifo[4][5] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\fifo.fifo[7][15] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\fifo.fifo[5][2] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\fifo.fifo[5][28] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\fifo.fifo[4][31] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\fifo.fifo[4][10] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\fifo.fifo[5][35] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\fifo.fifo[4][50] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\fifo.fifo[6][20] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\fifo.fifo[6][9] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\fifo.fifo[1][14] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\fifo.fifo[1][5] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\fifo.fifo[3][14] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\fifo.fifo[4][55] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\fifo.fifo[0][52] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\fifo.fifo[6][54] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\fifo.fifo[1][30] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\fifo.rd_data[34] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\fifo.fifo[5][42] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\fifo.fifo[6][45] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\fifo.fifo[2][9] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\fifo.fifo[1][34] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\fifo.fifo[5][43] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\fifo.fifo[1][7] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\fifo.fifo[0][41] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\fifo.fifo[3][20] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\fifo.fifo[6][6] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\fifo.fifo[0][15] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\fifo.fifo[0][42] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\fifo.fifo[4][19] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\fifo.fifo[1][45] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\fifo.fifo[3][36] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\fifo.fifo[1][43] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\fifo.fifo[2][41] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\fifo.fifo[2][4] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\fifo.fifo[5][15] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\fifo.fifo[2][22] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\fifo.rd_data[52] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\fifo.fifo[3][45] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\fifo.fifo[5][6] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\fifo.fifo[6][7] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\fifo.fifo[5][33] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\fifo.fifo[3][15] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\fifo.fifo[5][5] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\fifo.fifo[1][21] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\fifo.fifo[3][39] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\fifo.fifo[5][10] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\fifo.fifo[2][11] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\fifo.fifo[5][23] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\fifo.fifo[5][3] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\fifo.fifo[3][0] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\fifo.fifo[7][54] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\fifo.fifo[2][49] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\fifo.fifo[5][55] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\fifo.fifo[0][2] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\fifo.fifo[1][9] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\fifo.fifo[4][7] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\fifo.fifo[4][42] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\fifo.fifo[4][9] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\fifo.fifo[0][25] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\fifo.fifo[3][50] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\fifo.fifo[5][41] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\fifo.fifo[6][44] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\fifo.fifo[7][55] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\fifo.fifo[4][15] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\fifo.fifo[6][35] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\fifo.fifo[4][2] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\fifo.fifo[2][18] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\fifo.fifo[1][50] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\fifo.fifo[0][50] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\fifo.fifo[3][47] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\fifo.fifo[5][50] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\fifo.rd_data[12] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\fifo.fifo[6][12] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\fifo.fifo[5][19] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\fifo.fifo[0][30] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\fifo.rd_data[16] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\fifo.fifo[5][39] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\fifo.fifo[4][47] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\fifo.fifo[4][17] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\fifo.fifo[4][21] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\fifo.fifo[1][25] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\fifo.fifo[4][20] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\L[20] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\fifo.fifo[2][15] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\fifo.fifo[1][51] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\fifo.fifo[4][46] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\fifo.fifo[7][2] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\fifo.fifo[3][24] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\fifo.fifo[0][17] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\fifo.fifo[1][15] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\fifo.rd_data[33] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\fifo.fifo[3][6] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\fifo.fifo[4][37] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\fifo.fifo[2][39] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\fifo.fifo[6][5] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\fifo.fifo[4][23] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\fifo.fifo[4][38] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\fifo.fifo[4][13] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\fifo.fifo[5][22] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\fifo.fifo[0][10] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\fifo.fifo[4][40] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\fifo.fifo[7][52] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\fifo.rd_data[17] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\fifo.fifo[6][32] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\fifo.fifo[6][43] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\fifo.fifo[0][5] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\fifo.fifo[4][53] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\fifo.fifo[2][27] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\fifo.fifo[3][21] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\fifo.fifo[4][8] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\fifo.fifo[4][24] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\fifo.fifo[7][13] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\fifo.fifo[7][32] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\fifo.fifo[1][55] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\fifo.fifo[7][30] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\fifo.fifo[2][12] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\fifo.fifo[3][2] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\fifo.rd_data[47] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\fifo.fifo[7][40] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\fifo.rd_data[1] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\fifo.fifo[0][32] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\fifo.rd_data[45] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\fifo.fifo[0][29] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\fifo.fifo[2][43] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\fifo.fifo[5][54] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\fifo.fifo[7][37] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\fifo.fifo[2][28] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\fifo.fifo[2][3] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\fifo.fifo[4][39] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\fifo.fifo[5][26] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\fifo.fifo[7][49] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\fifo.fifo[1][28] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\fifo.fifo[2][33] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\fifo.rd_data[14] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\L[26] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\fifo.fifo[3][40] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\fifo.rd_data[43] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\fifo.fifo[5][40] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\fifo.fifo[6][50] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\fifo.fifo[6][48] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\fifo.fifo[3][29] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\fifo.fifo[1][17] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\fifo.fifo[2][55] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\fifo.fifo[5][16] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\fifo.fifo[0][48] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\fifo.fifo[1][1] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\fifo.fifo[7][50] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\fifo.fifo[3][52] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\fifo.fifo[5][30] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\fifo.fifo[3][41] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\fifo.fifo[0][37] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\fifo.fifo[7][22] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\fifo.fifo[5][9] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\fifo.fifo[2][47] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\fifo.fifo[0][24] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\fifo.fifo[5][0] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\fifo.fifo[4][30] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\fifo.fifo[3][32] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\fifo.fifo[7][51] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\fifo.fifo[7][12] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\fifo.fifo[3][53] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\fifo.fifo[6][29] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\fifo.fifo[6][36] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\fifo.fifo[0][54] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\fifo.fifo[6][18] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\fifo.fifo[1][52] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\fifo.fifo[4][27] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\fifo.fifo[6][19] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\fifo.rd_data[48] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\fifo.fifo[2][6] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\fifo.fifo[4][32] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\fifo.fifo[3][33] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\fifo.fifo[1][32] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\fifo.fifo[6][17] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\fifo.fifo[0][0] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\fifo.fifo[7][5] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\fifo.fifo[0][31] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\fifo.fifo[3][7] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\fifo.fifo[4][14] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\fifo.fifo[2][29] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\fifo.fifo[7][10] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\fifo.fifo[5][38] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\fifo.fifo[6][3] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\fifo.fifo[0][53] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\fifo.fifo[1][46] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\fifo.fifo[3][25] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\fifo.fifo[4][29] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\fifo.fifo[7][16] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\fifo.fifo[7][35] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\fifo.fifo[5][11] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\fifo.fifo[2][38] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\fifo.fifo[3][4] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\fifo.fifo[4][36] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\L[17] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\fifo.rd_data[18] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\fifo.rd_data[13] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\fifo.fifo[1][39] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\fifo.fifo[7][14] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\fifo.fifo[2][31] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\fifo.fifo[4][35] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\fifo.fifo[4][25] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\fifo.fifo[5][45] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\fifo.fifo[1][0] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\fifo.fifo[1][42] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\fifo.fifo[5][52] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\fifo.fifo[6][41] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\fifo.fifo[1][44] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\fifo.rd_data[42] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\fifo.fifo[4][44] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\fifo.fifo[5][25] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\fifo.rd_data[8] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\fifo.fifo[7][39] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\fifo.fifo[6][8] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\fifo.fifo[0][19] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\fifo.fifo[0][13] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\fifo.fifo[3][35] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\fifo.fifo[3][10] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\fifo.fifo[5][27] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\L[6] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\fifo.fifo[2][0] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\fifo.rd_data[35] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\fifo.fifo[5][18] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\fifo.fifo[2][1] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\fifo.fifo[6][24] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\fifo.fifo[1][20] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\fifo.fifo[3][3] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\fifo.fifo[7][42] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\fifo.fifo[2][46] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\L[30] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\fifo.fifo[1][53] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\fifo.fifo[5][14] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\fifo.fifo[1][10] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\fifo.fifo[6][40] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\fifo.fifo[7][1] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\fifo.fifo[2][19] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\fifo.fifo[7][38] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\fifo.fifo[6][31] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\fifo.fifo[1][6] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\fifo.rd_data[0] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\fifo.fifo[3][27] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\fifo.fifo[4][52] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\fifo.fifo[3][12] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\fifo.fifo[6][49] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\fifo.fifo[6][53] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\fifo.fifo[7][31] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\fifo.fifo[1][22] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\fifo.fifo[2][5] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\fifo.fifo[6][51] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\fifo.fifo[3][48] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\fifo.fifo[2][30] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\fifo.fifo[7][33] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\fifo.fifo[4][28] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\fifo.fifo[7][9] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\fifo.fifo[0][8] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\fifo.rd_data[5] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\fifo.fifo[3][30] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\fifo.fifo[7][18] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\fifo.fifo[6][52] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\fifo.fifo[4][26] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\fifo.fifo[5][1] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\fifo.fifo[5][8] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\fifo.fifo[0][28] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\fifo.fifo[0][49] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\fifo.fifo[6][23] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\fifo.fifo[7][3] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\fifo.fifo[4][22] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\fifo.fifo[4][48] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\fifo.fifo[4][43] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\fifo.fifo[2][2] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\fifo.fifo[6][37] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\fifo.fifo[6][15] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\fifo.fifo[1][26] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\fifo.fifo[4][12] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\fifo.fifo[3][5] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\fifo.fifo[7][6] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\fifo.rd_data[15] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\fifo.fifo[0][23] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\fifo.fifo[5][34] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\fifo.fifo[3][17] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\fifo.fifo[6][28] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\fifo.fifo[3][38] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\fifo.fifo[3][13] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\fifo.fifo[1][33] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\fifo.fifo[2][8] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\fifo.fifo[5][29] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\fifo.fifo[7][34] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\fifo.fifo[7][20] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\fifo.fifo[2][34] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\fifo.fifo[2][23] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\fifo.fifo[5][44] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\fifo.fifo[6][2] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\fifo.fifo[2][37] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\fifo.fifo[0][16] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\fifo.fifo[5][46] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\fifo.fifo[3][44] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\fifo.fifo[1][38] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\fifo.fifo[7][27] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\fifo.fifo[4][16] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\fifo.fifo[4][3] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\fifo.fifo[2][21] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\fifo.fifo[0][14] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\fifo.fifo[4][49] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\fifo.fifo[1][40] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\fifo.fifo[0][51] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\fifo.rd_data[19] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\fifo.fifo[1][35] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\fifo.fifo[7][36] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\fifo.fifo[6][27] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\fifo.fifo[4][0] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\fifo.fifo[3][16] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\fifo.fifo[4][41] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\fifo.fifo[0][33] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\fifo.fifo[2][17] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\fifo.fifo[5][47] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\fifo.fifo[6][34] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\fifo.fifo[2][35] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\fifo.fifo[0][3] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\fifo.fifo[6][13] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\fifo.fifo[2][14] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\fifo.fifo[3][18] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\fifo.fifo[1][4] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\fifo.fifo[3][19] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\fifo.fifo[2][16] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\fifo.rd_data[3] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\fifo.fifo[5][49] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\fifo.fifo[4][4] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\fifo.fifo[4][33] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\fifo.fifo[3][34] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\fifo.fifo[7][4] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\fifo.fifo[7][48] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\fifo.fifo[2][25] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\fifo.fifo[5][20] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\fifo.fifo[7][43] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\fifo.fifo[0][26] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\fifo.fifo[0][36] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\fifo.fifo[6][39] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\fifo.fifo[7][17] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\fifo.fifo[7][29] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\fifo.rd_data[46] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\fifo.fifo[2][10] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\fifo.fifo[4][34] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\fifo.fifo[0][11] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\fifo.fifo[3][54] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\fifo.fifo[2][53] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\fifo.fifo[6][16] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\fifo.fifo[6][14] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\fifo.fifo[6][11] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\fifo.fifo[0][43] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\fifo.fifo[2][13] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\fifo.rd_data[44] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\fifo.fifo[1][3] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\fifo.fifo[5][12] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\fifo.fifo[0][39] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\fifo.fifo[2][36] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\fifo.fifo[3][1] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\fifo.fifo[7][25] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\fifo.fifo[7][41] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\fifo.fifo[6][55] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\fifo.fifo[2][54] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\fifo.fifo[7][21] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\fifo.fifo[3][31] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\fifo.fifo[0][44] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\fifo.fifo[7][24] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\fifo.fifo[2][26] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\fifo.fifo[7][19] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\fifo.fifo[1][48] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\fifo.fifo[6][30] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\fifo.fifo[7][46] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\fifo.fifo[6][21] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\fifo.fifo[1][24] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\fifo.fifo[7][8] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\fifo.fifo[1][47] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\fifo.fifo[5][7] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\fifo.fifo[6][33] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\fifo.fifo[3][9] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\fifo.rd_data[54] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\fifo.fifo[5][13] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\counter_inst.count[4] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\fifo.fifo[7][28] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\fifo.fifo[2][7] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\fifo.fifo[6][25] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\fifo.fifo[7][11] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\fifo.fifo[5][37] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\fifo.fifo[7][44] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\fifo.fifo[1][31] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\fifo.fifo[7][26] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\fifo.rd_data[7] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\fifo.rd_data[21] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\fifo.fifo[2][32] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\fifo.fifo[7][53] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\fifo.fifo[7][23] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\fifo.rd_data[22] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\fifo.fifo[7][7] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\fifo.fifo[4][51] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\fifo.rd_data[55] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\fifo.rd_data[30] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\fifo.fifo[0][7] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\fifo.fifo[6][10] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\fifo.rd_data[28] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\L[14] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\fifo.fifo[0][45] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\fifo.rd_data[9] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\fifo.fifo[7][45] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\fifo.fifo[7][47] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\fifo.fifo[2][24] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\fifo.fifo[1][8] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\fifo.fifo[3][26] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\fifo.fifo[6][26] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\fifo.rd_data[11] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\fifo.rd_data[2] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\fifo.rd_data[31] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\fifo.rd_data[4] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\L[29] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(net131),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\fifo.rd_data[24] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0568_),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\fifo.fifo[3][46] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0573_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(net165),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(net177),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\fifo.fifo[6][38] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(net155),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\fifo.rd_data[6] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(net148),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(net154),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\fifo.rd_data[10] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\L[27] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\fifo.fifo[4][6] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\fifo.rd_data[20] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(net138),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\L[11] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\fifo.rd_data[41] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\L[5] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\L[23] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(net179),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(net151),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\fifo.rd_data[37] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(net137),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\fifo.fifo[0][6] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(net171),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\L[3] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\L[22] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\L[18] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\fifo.rd_data[25] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\R[15] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\L[1] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\L[9] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\R[30] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(net187),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\fifo.fifo[5][53] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(net174),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(net167),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\R[21] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\L[10] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\fifo.rd_data[23] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\L[19] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\fifo.rd_data[36] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(net144),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\L[2] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\L[28] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\fifo.fifo[0][46] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\R[3] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\L[13] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\R[19] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\fifo.rd_data[39] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\fifo.rd_data[24] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\fifo.rd_data[39] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\fifo.rd_data[4] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\fifo.fifo[3][28] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\fifo.fifo[0][47] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\fifo.fifo[6][47] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\fifo.fifo[1][18] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\fifo.fifo[1][13] ),
    .X(net247));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold6 (.A(\fifo.rd_data[26] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\fifo.fifo[2][52] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\fifo.fifo[3][8] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\fifo.fifo[1][37] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\fifo.fifo[6][42] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\fifo.fifo[5][51] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\fifo.fifo[6][1] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\fifo.fifo[2][42] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\fifo.fifo[0][55] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\fifo.fifo[0][4] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\L[8] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\fifo.fifo[1][27] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\fifo.fifo[0][35] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\fifo.fifo[4][11] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\fifo.fifo[3][23] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\fifo.fifo[0][20] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\fifo.fifo[0][27] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\fifo.fifo[4][18] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\fifo.fifo[4][54] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\fifo.fifo[3][22] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\fifo.fifo[5][36] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\fifo.fifo[6][0] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\fifo.fifo[2][48] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\fifo.fifo[1][29] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\fifo.fifo[3][42] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\fifo.fifo[1][12] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\fifo.fifo[2][40] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\fifo.fifo[0][38] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\fifo.fifo[1][16] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\fifo.fifo[3][37] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\fifo.rd_data[53] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\fifo.fifo[2][20] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\fifo.fifo[3][55] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\fifo.fifo[5][21] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\fifo.fifo[0][21] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\fifo.rd_data[27] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\fifo.fifo[3][49] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\fifo.fifo[0][34] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\fifo.fifo[0][9] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\fifo.fifo[3][43] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\fifo.fifo[5][48] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\fifo.fifo[6][46] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\fifo.fifo[5][17] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\fifo.fifo[3][11] ),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(decrypt),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(desIn[17]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input100 (.A(key[3]),
    .X(net100));
 sky130_fd_sc_hd__buf_4 input101 (.A(key[40]),
    .X(net101));
 sky130_fd_sc_hd__buf_4 input102 (.A(key[41]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(key[42]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 input104 (.A(key[43]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(key[44]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(key[45]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_8 input107 (.A(key[46]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 input108 (.A(key[47]),
    .X(net108));
 sky130_fd_sc_hd__buf_4 input109 (.A(key[48]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(desIn[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input110 (.A(key[49]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_8 input111 (.A(key[4]),
    .X(net111));
 sky130_fd_sc_hd__buf_4 input112 (.A(key[50]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(key[51]),
    .X(net113));
 sky130_fd_sc_hd__buf_4 input114 (.A(key[52]),
    .X(net114));
 sky130_fd_sc_hd__buf_2 input115 (.A(key[53]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_8 input116 (.A(key[54]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_8 input117 (.A(key[55]),
    .X(net117));
 sky130_fd_sc_hd__buf_4 input118 (.A(key[5]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_8 input119 (.A(key[6]),
    .X(net119));
 sky130_fd_sc_hd__buf_4 input12 (.A(desIn[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_8 input120 (.A(key[7]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(key[8]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 input122 (.A(key[9]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 input123 (.A(reset),
    .X(net123));
 sky130_fd_sc_hd__buf_2 input13 (.A(desIn[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(desIn[20]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(desIn[21]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(desIn[22]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(desIn[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(desIn[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(desIn[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(desIn[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(desIn[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(desIn[27]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(desIn[28]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(desIn[29]),
    .X(net23));
 sky130_fd_sc_hd__buf_4 input24 (.A(desIn[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(desIn[30]),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(desIn[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(desIn[32]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(desIn[33]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(desIn[34]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(desIn[10]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input30 (.A(desIn[35]),
    .X(net30));
 sky130_fd_sc_hd__buf_4 input31 (.A(desIn[36]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(desIn[37]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(desIn[38]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(desIn[39]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(desIn[3]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(desIn[40]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(desIn[41]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(desIn[42]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(desIn[43]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input4 (.A(desIn[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(desIn[44]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(desIn[45]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(desIn[46]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(desIn[47]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(desIn[48]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(desIn[49]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(desIn[4]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(desIn[50]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(desIn[51]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 input49 (.A(desIn[52]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input5 (.A(desIn[12]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input50 (.A(desIn[53]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(desIn[54]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(desIn[55]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(desIn[56]),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input54 (.A(desIn[57]),
    .X(net54));
 sky130_fd_sc_hd__buf_2 input55 (.A(desIn[58]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(desIn[59]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 input57 (.A(desIn[5]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(desIn[60]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(desIn[61]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(desIn[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(desIn[62]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(desIn[63]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 input62 (.A(desIn[6]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 input63 (.A(desIn[7]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(desIn[8]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(desIn[9]),
    .X(net65));
 sky130_fd_sc_hd__buf_4 input66 (.A(init),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 input67 (.A(key[0]),
    .X(net67));
 sky130_fd_sc_hd__buf_4 input68 (.A(key[10]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(key[11]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(desIn[14]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input70 (.A(key[12]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 input71 (.A(key[13]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 input72 (.A(key[14]),
    .X(net72));
 sky130_fd_sc_hd__buf_4 input73 (.A(key[15]),
    .X(net73));
 sky130_fd_sc_hd__buf_4 input74 (.A(key[16]),
    .X(net74));
 sky130_fd_sc_hd__buf_4 input75 (.A(key[17]),
    .X(net75));
 sky130_fd_sc_hd__buf_4 input76 (.A(key[18]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 input77 (.A(key[19]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input78 (.A(key[1]),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(key[20]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(desIn[15]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input80 (.A(key[21]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(key[22]),
    .X(net81));
 sky130_fd_sc_hd__buf_4 input82 (.A(key[23]),
    .X(net82));
 sky130_fd_sc_hd__buf_4 input83 (.A(key[24]),
    .X(net83));
 sky130_fd_sc_hd__buf_4 input84 (.A(key[25]),
    .X(net84));
 sky130_fd_sc_hd__buf_4 input85 (.A(key[26]),
    .X(net85));
 sky130_fd_sc_hd__buf_4 input86 (.A(key[27]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(key[28]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_8 input88 (.A(key[29]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 input89 (.A(key[2]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(desIn[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_6 input90 (.A(key[30]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_8 input91 (.A(key[31]),
    .X(net91));
 sky130_fd_sc_hd__buf_4 input92 (.A(key[32]),
    .X(net92));
 sky130_fd_sc_hd__buf_4 input93 (.A(key[33]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 input94 (.A(key[34]),
    .X(net94));
 sky130_fd_sc_hd__buf_2 input95 (.A(key[35]),
    .X(net95));
 sky130_fd_sc_hd__buf_4 input96 (.A(key[36]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 input97 (.A(key[37]),
    .X(net97));
 sky130_fd_sc_hd__buf_4 input98 (.A(key[38]),
    .X(net98));
 sky130_fd_sc_hd__buf_4 input99 (.A(key[39]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 output124 (.A(net124),
    .X(desOut_ff[0]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(desOut_ff[10]));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net126),
    .X(desOut_ff[11]));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net127),
    .X(desOut_ff[12]));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net128),
    .X(desOut_ff[13]));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net129),
    .X(desOut_ff[14]));
 sky130_fd_sc_hd__clkbuf_4 output130 (.A(net130),
    .X(desOut_ff[15]));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net131),
    .X(desOut_ff[16]));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net132),
    .X(desOut_ff[17]));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net133),
    .X(desOut_ff[18]));
 sky130_fd_sc_hd__clkbuf_4 output134 (.A(net134),
    .X(desOut_ff[19]));
 sky130_fd_sc_hd__clkbuf_4 output135 (.A(net135),
    .X(desOut_ff[1]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(desOut_ff[20]));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net137),
    .X(desOut_ff[21]));
 sky130_fd_sc_hd__clkbuf_4 output138 (.A(net138),
    .X(desOut_ff[22]));
 sky130_fd_sc_hd__clkbuf_4 output139 (.A(net139),
    .X(desOut_ff[23]));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net140),
    .X(desOut_ff[24]));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net141),
    .X(desOut_ff[25]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(desOut_ff[26]));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net143),
    .X(desOut_ff[27]));
 sky130_fd_sc_hd__clkbuf_4 output144 (.A(net144),
    .X(desOut_ff[28]));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net145),
    .X(desOut_ff[29]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(desOut_ff[2]));
 sky130_fd_sc_hd__clkbuf_4 output147 (.A(net147),
    .X(desOut_ff[30]));
 sky130_fd_sc_hd__clkbuf_4 output148 (.A(net148),
    .X(desOut_ff[31]));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net149),
    .X(desOut_ff[32]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(desOut_ff[33]));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net151),
    .X(desOut_ff[34]));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net152),
    .X(desOut_ff[35]));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net153),
    .X(desOut_ff[36]));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net154),
    .X(desOut_ff[37]));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net155),
    .X(desOut_ff[38]));
 sky130_fd_sc_hd__clkbuf_4 output156 (.A(net156),
    .X(desOut_ff[39]));
 sky130_fd_sc_hd__clkbuf_4 output157 (.A(net157),
    .X(desOut_ff[3]));
 sky130_fd_sc_hd__clkbuf_4 output158 (.A(net158),
    .X(desOut_ff[40]));
 sky130_fd_sc_hd__clkbuf_4 output159 (.A(net159),
    .X(desOut_ff[41]));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net160),
    .X(desOut_ff[42]));
 sky130_fd_sc_hd__clkbuf_4 output161 (.A(net161),
    .X(desOut_ff[43]));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net162),
    .X(desOut_ff[44]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(desOut_ff[45]));
 sky130_fd_sc_hd__clkbuf_4 output164 (.A(net164),
    .X(desOut_ff[46]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(desOut_ff[47]));
 sky130_fd_sc_hd__clkbuf_4 output166 (.A(net166),
    .X(desOut_ff[48]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(desOut_ff[49]));
 sky130_fd_sc_hd__clkbuf_4 output168 (.A(net168),
    .X(desOut_ff[4]));
 sky130_fd_sc_hd__clkbuf_4 output169 (.A(net169),
    .X(desOut_ff[50]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(desOut_ff[51]));
 sky130_fd_sc_hd__clkbuf_4 output171 (.A(net171),
    .X(desOut_ff[52]));
 sky130_fd_sc_hd__clkbuf_4 output172 (.A(net172),
    .X(desOut_ff[53]));
 sky130_fd_sc_hd__clkbuf_4 output173 (.A(net173),
    .X(desOut_ff[54]));
 sky130_fd_sc_hd__clkbuf_4 output174 (.A(net174),
    .X(desOut_ff[55]));
 sky130_fd_sc_hd__clkbuf_4 output175 (.A(net175),
    .X(desOut_ff[56]));
 sky130_fd_sc_hd__clkbuf_4 output176 (.A(net176),
    .X(desOut_ff[57]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(desOut_ff[58]));
 sky130_fd_sc_hd__clkbuf_4 output178 (.A(net178),
    .X(desOut_ff[59]));
 sky130_fd_sc_hd__clkbuf_4 output179 (.A(net179),
    .X(desOut_ff[5]));
 sky130_fd_sc_hd__clkbuf_4 output180 (.A(net180),
    .X(desOut_ff[60]));
 sky130_fd_sc_hd__clkbuf_4 output181 (.A(net181),
    .X(desOut_ff[61]));
 sky130_fd_sc_hd__clkbuf_4 output182 (.A(net182),
    .X(desOut_ff[62]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(desOut_ff[63]));
 sky130_fd_sc_hd__clkbuf_4 output184 (.A(net184),
    .X(desOut_ff[6]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(desOut_ff[7]));
 sky130_fd_sc_hd__clkbuf_4 output186 (.A(net186),
    .X(desOut_ff[8]));
 sky130_fd_sc_hd__clkbuf_4 output187 (.A(net187),
    .X(desOut_ff[9]));
 sky130_fd_sc_hd__clkbuf_4 output188 (.A(net188),
    .X(finish));
endmodule

