// This is the unpowered netlist.
module aes (clk,
    decrypt_i,
    load_i,
    ready_o,
    reset,
    data_i,
    data_o,
    key_i);
 input clk;
 input decrypt_i;
 input load_i;
 output ready_o;
 input reset;
 input [127:0] data_i;
 output [127:0] data_o;
 input [127:0] key_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire addroundkey_ready_o;
 wire \addroundkey_round[0] ;
 wire \addroundkey_round[1] ;
 wire \addroundkey_round[2] ;
 wire \addroundkey_round[3] ;
 wire addroundkey_start_i;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire first_round_reg;
 wire \ks1.col[0] ;
 wire \ks1.col[16] ;
 wire \ks1.col[17] ;
 wire \ks1.col[18] ;
 wire \ks1.col[19] ;
 wire \ks1.col[1] ;
 wire \ks1.col[20] ;
 wire \ks1.col[21] ;
 wire \ks1.col[22] ;
 wire \ks1.col[23] ;
 wire \ks1.col[24] ;
 wire \ks1.col[25] ;
 wire \ks1.col[26] ;
 wire \ks1.col[27] ;
 wire \ks1.col[28] ;
 wire \ks1.col[29] ;
 wire \ks1.col[2] ;
 wire \ks1.col[30] ;
 wire \ks1.col[31] ;
 wire \ks1.col[3] ;
 wire \ks1.col[4] ;
 wire \ks1.col[5] ;
 wire \ks1.col[6] ;
 wire \ks1.col[7] ;
 wire \ks1.key_reg[0] ;
 wire \ks1.key_reg[100] ;
 wire \ks1.key_reg[101] ;
 wire \ks1.key_reg[102] ;
 wire \ks1.key_reg[103] ;
 wire \ks1.key_reg[104] ;
 wire \ks1.key_reg[105] ;
 wire \ks1.key_reg[106] ;
 wire \ks1.key_reg[107] ;
 wire \ks1.key_reg[108] ;
 wire \ks1.key_reg[109] ;
 wire \ks1.key_reg[10] ;
 wire \ks1.key_reg[110] ;
 wire \ks1.key_reg[111] ;
 wire \ks1.key_reg[112] ;
 wire \ks1.key_reg[113] ;
 wire \ks1.key_reg[114] ;
 wire \ks1.key_reg[115] ;
 wire \ks1.key_reg[116] ;
 wire \ks1.key_reg[117] ;
 wire \ks1.key_reg[118] ;
 wire \ks1.key_reg[119] ;
 wire \ks1.key_reg[11] ;
 wire \ks1.key_reg[120] ;
 wire \ks1.key_reg[121] ;
 wire \ks1.key_reg[122] ;
 wire \ks1.key_reg[123] ;
 wire \ks1.key_reg[124] ;
 wire \ks1.key_reg[125] ;
 wire \ks1.key_reg[126] ;
 wire \ks1.key_reg[127] ;
 wire \ks1.key_reg[12] ;
 wire \ks1.key_reg[13] ;
 wire \ks1.key_reg[14] ;
 wire \ks1.key_reg[15] ;
 wire \ks1.key_reg[16] ;
 wire \ks1.key_reg[17] ;
 wire \ks1.key_reg[18] ;
 wire \ks1.key_reg[19] ;
 wire \ks1.key_reg[1] ;
 wire \ks1.key_reg[20] ;
 wire \ks1.key_reg[21] ;
 wire \ks1.key_reg[22] ;
 wire \ks1.key_reg[23] ;
 wire \ks1.key_reg[24] ;
 wire \ks1.key_reg[25] ;
 wire \ks1.key_reg[26] ;
 wire \ks1.key_reg[27] ;
 wire \ks1.key_reg[28] ;
 wire \ks1.key_reg[29] ;
 wire \ks1.key_reg[2] ;
 wire \ks1.key_reg[30] ;
 wire \ks1.key_reg[31] ;
 wire \ks1.key_reg[32] ;
 wire \ks1.key_reg[33] ;
 wire \ks1.key_reg[34] ;
 wire \ks1.key_reg[35] ;
 wire \ks1.key_reg[36] ;
 wire \ks1.key_reg[37] ;
 wire \ks1.key_reg[38] ;
 wire \ks1.key_reg[39] ;
 wire \ks1.key_reg[3] ;
 wire \ks1.key_reg[40] ;
 wire \ks1.key_reg[41] ;
 wire \ks1.key_reg[42] ;
 wire \ks1.key_reg[43] ;
 wire \ks1.key_reg[44] ;
 wire \ks1.key_reg[45] ;
 wire \ks1.key_reg[46] ;
 wire \ks1.key_reg[47] ;
 wire \ks1.key_reg[48] ;
 wire \ks1.key_reg[49] ;
 wire \ks1.key_reg[4] ;
 wire \ks1.key_reg[50] ;
 wire \ks1.key_reg[51] ;
 wire \ks1.key_reg[52] ;
 wire \ks1.key_reg[53] ;
 wire \ks1.key_reg[54] ;
 wire \ks1.key_reg[55] ;
 wire \ks1.key_reg[56] ;
 wire \ks1.key_reg[57] ;
 wire \ks1.key_reg[58] ;
 wire \ks1.key_reg[59] ;
 wire \ks1.key_reg[5] ;
 wire \ks1.key_reg[60] ;
 wire \ks1.key_reg[61] ;
 wire \ks1.key_reg[62] ;
 wire \ks1.key_reg[63] ;
 wire \ks1.key_reg[64] ;
 wire \ks1.key_reg[65] ;
 wire \ks1.key_reg[66] ;
 wire \ks1.key_reg[67] ;
 wire \ks1.key_reg[68] ;
 wire \ks1.key_reg[69] ;
 wire \ks1.key_reg[6] ;
 wire \ks1.key_reg[70] ;
 wire \ks1.key_reg[71] ;
 wire \ks1.key_reg[72] ;
 wire \ks1.key_reg[73] ;
 wire \ks1.key_reg[74] ;
 wire \ks1.key_reg[75] ;
 wire \ks1.key_reg[76] ;
 wire \ks1.key_reg[77] ;
 wire \ks1.key_reg[78] ;
 wire \ks1.key_reg[79] ;
 wire \ks1.key_reg[7] ;
 wire \ks1.key_reg[80] ;
 wire \ks1.key_reg[81] ;
 wire \ks1.key_reg[82] ;
 wire \ks1.key_reg[83] ;
 wire \ks1.key_reg[84] ;
 wire \ks1.key_reg[85] ;
 wire \ks1.key_reg[86] ;
 wire \ks1.key_reg[87] ;
 wire \ks1.key_reg[88] ;
 wire \ks1.key_reg[89] ;
 wire \ks1.key_reg[8] ;
 wire \ks1.key_reg[90] ;
 wire \ks1.key_reg[91] ;
 wire \ks1.key_reg[92] ;
 wire \ks1.key_reg[93] ;
 wire \ks1.key_reg[94] ;
 wire \ks1.key_reg[95] ;
 wire \ks1.key_reg[96] ;
 wire \ks1.key_reg[97] ;
 wire \ks1.key_reg[98] ;
 wire \ks1.key_reg[99] ;
 wire \ks1.key_reg[9] ;
 wire \ks1.next_ready_o ;
 wire \ks1.ready_o ;
 wire \ks1.state[0] ;
 wire \ks1.state[1] ;
 wire \ks1.state[2] ;
 wire \mix1.data_o[0] ;
 wire \mix1.data_o[100] ;
 wire \mix1.data_o[101] ;
 wire \mix1.data_o[102] ;
 wire \mix1.data_o[103] ;
 wire \mix1.data_o[104] ;
 wire \mix1.data_o[105] ;
 wire \mix1.data_o[106] ;
 wire \mix1.data_o[107] ;
 wire \mix1.data_o[108] ;
 wire \mix1.data_o[109] ;
 wire \mix1.data_o[10] ;
 wire \mix1.data_o[110] ;
 wire \mix1.data_o[111] ;
 wire \mix1.data_o[112] ;
 wire \mix1.data_o[113] ;
 wire \mix1.data_o[114] ;
 wire \mix1.data_o[115] ;
 wire \mix1.data_o[116] ;
 wire \mix1.data_o[117] ;
 wire \mix1.data_o[118] ;
 wire \mix1.data_o[119] ;
 wire \mix1.data_o[11] ;
 wire \mix1.data_o[120] ;
 wire \mix1.data_o[121] ;
 wire \mix1.data_o[122] ;
 wire \mix1.data_o[123] ;
 wire \mix1.data_o[124] ;
 wire \mix1.data_o[125] ;
 wire \mix1.data_o[126] ;
 wire \mix1.data_o[127] ;
 wire \mix1.data_o[12] ;
 wire \mix1.data_o[13] ;
 wire \mix1.data_o[14] ;
 wire \mix1.data_o[15] ;
 wire \mix1.data_o[16] ;
 wire \mix1.data_o[17] ;
 wire \mix1.data_o[18] ;
 wire \mix1.data_o[19] ;
 wire \mix1.data_o[1] ;
 wire \mix1.data_o[20] ;
 wire \mix1.data_o[21] ;
 wire \mix1.data_o[22] ;
 wire \mix1.data_o[23] ;
 wire \mix1.data_o[24] ;
 wire \mix1.data_o[25] ;
 wire \mix1.data_o[26] ;
 wire \mix1.data_o[27] ;
 wire \mix1.data_o[28] ;
 wire \mix1.data_o[29] ;
 wire \mix1.data_o[2] ;
 wire \mix1.data_o[30] ;
 wire \mix1.data_o[31] ;
 wire \mix1.data_o[32] ;
 wire \mix1.data_o[33] ;
 wire \mix1.data_o[34] ;
 wire \mix1.data_o[35] ;
 wire \mix1.data_o[36] ;
 wire \mix1.data_o[37] ;
 wire \mix1.data_o[38] ;
 wire \mix1.data_o[39] ;
 wire \mix1.data_o[3] ;
 wire \mix1.data_o[40] ;
 wire \mix1.data_o[41] ;
 wire \mix1.data_o[42] ;
 wire \mix1.data_o[43] ;
 wire \mix1.data_o[44] ;
 wire \mix1.data_o[45] ;
 wire \mix1.data_o[46] ;
 wire \mix1.data_o[47] ;
 wire \mix1.data_o[48] ;
 wire \mix1.data_o[49] ;
 wire \mix1.data_o[4] ;
 wire \mix1.data_o[50] ;
 wire \mix1.data_o[51] ;
 wire \mix1.data_o[52] ;
 wire \mix1.data_o[53] ;
 wire \mix1.data_o[54] ;
 wire \mix1.data_o[55] ;
 wire \mix1.data_o[56] ;
 wire \mix1.data_o[57] ;
 wire \mix1.data_o[58] ;
 wire \mix1.data_o[59] ;
 wire \mix1.data_o[5] ;
 wire \mix1.data_o[60] ;
 wire \mix1.data_o[61] ;
 wire \mix1.data_o[62] ;
 wire \mix1.data_o[63] ;
 wire \mix1.data_o[64] ;
 wire \mix1.data_o[65] ;
 wire \mix1.data_o[66] ;
 wire \mix1.data_o[67] ;
 wire \mix1.data_o[68] ;
 wire \mix1.data_o[69] ;
 wire \mix1.data_o[6] ;
 wire \mix1.data_o[70] ;
 wire \mix1.data_o[71] ;
 wire \mix1.data_o[72] ;
 wire \mix1.data_o[73] ;
 wire \mix1.data_o[74] ;
 wire \mix1.data_o[75] ;
 wire \mix1.data_o[76] ;
 wire \mix1.data_o[77] ;
 wire \mix1.data_o[78] ;
 wire \mix1.data_o[79] ;
 wire \mix1.data_o[7] ;
 wire \mix1.data_o[80] ;
 wire \mix1.data_o[81] ;
 wire \mix1.data_o[82] ;
 wire \mix1.data_o[83] ;
 wire \mix1.data_o[84] ;
 wire \mix1.data_o[85] ;
 wire \mix1.data_o[86] ;
 wire \mix1.data_o[87] ;
 wire \mix1.data_o[88] ;
 wire \mix1.data_o[89] ;
 wire \mix1.data_o[8] ;
 wire \mix1.data_o[90] ;
 wire \mix1.data_o[91] ;
 wire \mix1.data_o[92] ;
 wire \mix1.data_o[93] ;
 wire \mix1.data_o[94] ;
 wire \mix1.data_o[95] ;
 wire \mix1.data_o[96] ;
 wire \mix1.data_o[97] ;
 wire \mix1.data_o[98] ;
 wire \mix1.data_o[99] ;
 wire \mix1.data_o[9] ;
 wire \mix1.data_reg[100] ;
 wire \mix1.data_reg[101] ;
 wire \mix1.data_reg[102] ;
 wire \mix1.data_reg[103] ;
 wire \mix1.data_reg[104] ;
 wire \mix1.data_reg[105] ;
 wire \mix1.data_reg[106] ;
 wire \mix1.data_reg[107] ;
 wire \mix1.data_reg[108] ;
 wire \mix1.data_reg[109] ;
 wire \mix1.data_reg[110] ;
 wire \mix1.data_reg[111] ;
 wire \mix1.data_reg[112] ;
 wire \mix1.data_reg[113] ;
 wire \mix1.data_reg[114] ;
 wire \mix1.data_reg[115] ;
 wire \mix1.data_reg[116] ;
 wire \mix1.data_reg[117] ;
 wire \mix1.data_reg[118] ;
 wire \mix1.data_reg[119] ;
 wire \mix1.data_reg[120] ;
 wire \mix1.data_reg[121] ;
 wire \mix1.data_reg[122] ;
 wire \mix1.data_reg[123] ;
 wire \mix1.data_reg[124] ;
 wire \mix1.data_reg[125] ;
 wire \mix1.data_reg[126] ;
 wire \mix1.data_reg[127] ;
 wire \mix1.data_reg[32] ;
 wire \mix1.data_reg[33] ;
 wire \mix1.data_reg[34] ;
 wire \mix1.data_reg[35] ;
 wire \mix1.data_reg[36] ;
 wire \mix1.data_reg[37] ;
 wire \mix1.data_reg[38] ;
 wire \mix1.data_reg[39] ;
 wire \mix1.data_reg[40] ;
 wire \mix1.data_reg[41] ;
 wire \mix1.data_reg[42] ;
 wire \mix1.data_reg[43] ;
 wire \mix1.data_reg[44] ;
 wire \mix1.data_reg[45] ;
 wire \mix1.data_reg[46] ;
 wire \mix1.data_reg[47] ;
 wire \mix1.data_reg[48] ;
 wire \mix1.data_reg[49] ;
 wire \mix1.data_reg[50] ;
 wire \mix1.data_reg[51] ;
 wire \mix1.data_reg[52] ;
 wire \mix1.data_reg[53] ;
 wire \mix1.data_reg[54] ;
 wire \mix1.data_reg[55] ;
 wire \mix1.data_reg[56] ;
 wire \mix1.data_reg[57] ;
 wire \mix1.data_reg[58] ;
 wire \mix1.data_reg[59] ;
 wire \mix1.data_reg[60] ;
 wire \mix1.data_reg[61] ;
 wire \mix1.data_reg[62] ;
 wire \mix1.data_reg[63] ;
 wire \mix1.data_reg[64] ;
 wire \mix1.data_reg[65] ;
 wire \mix1.data_reg[66] ;
 wire \mix1.data_reg[67] ;
 wire \mix1.data_reg[68] ;
 wire \mix1.data_reg[69] ;
 wire \mix1.data_reg[70] ;
 wire \mix1.data_reg[71] ;
 wire \mix1.data_reg[72] ;
 wire \mix1.data_reg[73] ;
 wire \mix1.data_reg[74] ;
 wire \mix1.data_reg[75] ;
 wire \mix1.data_reg[76] ;
 wire \mix1.data_reg[77] ;
 wire \mix1.data_reg[78] ;
 wire \mix1.data_reg[79] ;
 wire \mix1.data_reg[80] ;
 wire \mix1.data_reg[81] ;
 wire \mix1.data_reg[82] ;
 wire \mix1.data_reg[83] ;
 wire \mix1.data_reg[84] ;
 wire \mix1.data_reg[85] ;
 wire \mix1.data_reg[86] ;
 wire \mix1.data_reg[87] ;
 wire \mix1.data_reg[88] ;
 wire \mix1.data_reg[89] ;
 wire \mix1.data_reg[90] ;
 wire \mix1.data_reg[91] ;
 wire \mix1.data_reg[92] ;
 wire \mix1.data_reg[93] ;
 wire \mix1.data_reg[94] ;
 wire \mix1.data_reg[95] ;
 wire \mix1.data_reg[96] ;
 wire \mix1.data_reg[97] ;
 wire \mix1.data_reg[98] ;
 wire \mix1.data_reg[99] ;
 wire \mix1.next_ready_o ;
 wire \mix1.ready_o ;
 wire \mix1.state[0] ;
 wire \mix1.state[1] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire next_addroundkey_ready_o;
 wire next_addroundkey_start_i;
 wire next_first_round_reg;
 wire next_ready_o;
 wire next_state;
 wire \round[0] ;
 wire \round[1] ;
 wire \round[2] ;
 wire \round[3] ;
 wire \sbox1.ah[0] ;
 wire \sbox1.ah[1] ;
 wire \sbox1.ah[2] ;
 wire \sbox1.ah[3] ;
 wire \sbox1.ah_reg[0] ;
 wire \sbox1.ah_reg[1] ;
 wire \sbox1.ah_reg[2] ;
 wire \sbox1.ah_reg[3] ;
 wire \sbox1.alph[0] ;
 wire \sbox1.alph[1] ;
 wire \sbox1.alph[2] ;
 wire \sbox1.alph[3] ;
 wire \sbox1.intermediate_to_invert_var[0] ;
 wire \sbox1.intermediate_to_invert_var[1] ;
 wire \sbox1.intermediate_to_invert_var[2] ;
 wire \sbox1.intermediate_to_invert_var[3] ;
 wire \sbox1.inversion_to_invert_var[0] ;
 wire \sbox1.inversion_to_invert_var[1] ;
 wire \sbox1.inversion_to_invert_var[2] ;
 wire \sbox1.inversion_to_invert_var[3] ;
 wire \sbox1.next_alph[0] ;
 wire \sbox1.next_alph[1] ;
 wire \sbox1.next_alph[2] ;
 wire \sbox1.next_alph[3] ;
 wire state;
 wire \sub1.data_o[0] ;
 wire \sub1.data_o[100] ;
 wire \sub1.data_o[101] ;
 wire \sub1.data_o[102] ;
 wire \sub1.data_o[103] ;
 wire \sub1.data_o[104] ;
 wire \sub1.data_o[105] ;
 wire \sub1.data_o[106] ;
 wire \sub1.data_o[107] ;
 wire \sub1.data_o[108] ;
 wire \sub1.data_o[109] ;
 wire \sub1.data_o[10] ;
 wire \sub1.data_o[110] ;
 wire \sub1.data_o[111] ;
 wire \sub1.data_o[112] ;
 wire \sub1.data_o[113] ;
 wire \sub1.data_o[114] ;
 wire \sub1.data_o[115] ;
 wire \sub1.data_o[116] ;
 wire \sub1.data_o[117] ;
 wire \sub1.data_o[118] ;
 wire \sub1.data_o[119] ;
 wire \sub1.data_o[11] ;
 wire \sub1.data_o[120] ;
 wire \sub1.data_o[121] ;
 wire \sub1.data_o[122] ;
 wire \sub1.data_o[123] ;
 wire \sub1.data_o[124] ;
 wire \sub1.data_o[125] ;
 wire \sub1.data_o[126] ;
 wire \sub1.data_o[127] ;
 wire \sub1.data_o[12] ;
 wire \sub1.data_o[13] ;
 wire \sub1.data_o[14] ;
 wire \sub1.data_o[15] ;
 wire \sub1.data_o[16] ;
 wire \sub1.data_o[17] ;
 wire \sub1.data_o[18] ;
 wire \sub1.data_o[19] ;
 wire \sub1.data_o[1] ;
 wire \sub1.data_o[20] ;
 wire \sub1.data_o[21] ;
 wire \sub1.data_o[22] ;
 wire \sub1.data_o[23] ;
 wire \sub1.data_o[24] ;
 wire \sub1.data_o[25] ;
 wire \sub1.data_o[26] ;
 wire \sub1.data_o[27] ;
 wire \sub1.data_o[28] ;
 wire \sub1.data_o[29] ;
 wire \sub1.data_o[2] ;
 wire \sub1.data_o[30] ;
 wire \sub1.data_o[31] ;
 wire \sub1.data_o[32] ;
 wire \sub1.data_o[33] ;
 wire \sub1.data_o[34] ;
 wire \sub1.data_o[35] ;
 wire \sub1.data_o[36] ;
 wire \sub1.data_o[37] ;
 wire \sub1.data_o[38] ;
 wire \sub1.data_o[39] ;
 wire \sub1.data_o[3] ;
 wire \sub1.data_o[40] ;
 wire \sub1.data_o[41] ;
 wire \sub1.data_o[42] ;
 wire \sub1.data_o[43] ;
 wire \sub1.data_o[44] ;
 wire \sub1.data_o[45] ;
 wire \sub1.data_o[46] ;
 wire \sub1.data_o[47] ;
 wire \sub1.data_o[48] ;
 wire \sub1.data_o[49] ;
 wire \sub1.data_o[4] ;
 wire \sub1.data_o[50] ;
 wire \sub1.data_o[51] ;
 wire \sub1.data_o[52] ;
 wire \sub1.data_o[53] ;
 wire \sub1.data_o[54] ;
 wire \sub1.data_o[55] ;
 wire \sub1.data_o[56] ;
 wire \sub1.data_o[57] ;
 wire \sub1.data_o[58] ;
 wire \sub1.data_o[59] ;
 wire \sub1.data_o[5] ;
 wire \sub1.data_o[60] ;
 wire \sub1.data_o[61] ;
 wire \sub1.data_o[62] ;
 wire \sub1.data_o[63] ;
 wire \sub1.data_o[64] ;
 wire \sub1.data_o[65] ;
 wire \sub1.data_o[66] ;
 wire \sub1.data_o[67] ;
 wire \sub1.data_o[68] ;
 wire \sub1.data_o[69] ;
 wire \sub1.data_o[6] ;
 wire \sub1.data_o[70] ;
 wire \sub1.data_o[71] ;
 wire \sub1.data_o[72] ;
 wire \sub1.data_o[73] ;
 wire \sub1.data_o[74] ;
 wire \sub1.data_o[75] ;
 wire \sub1.data_o[76] ;
 wire \sub1.data_o[77] ;
 wire \sub1.data_o[78] ;
 wire \sub1.data_o[79] ;
 wire \sub1.data_o[7] ;
 wire \sub1.data_o[80] ;
 wire \sub1.data_o[81] ;
 wire \sub1.data_o[82] ;
 wire \sub1.data_o[83] ;
 wire \sub1.data_o[84] ;
 wire \sub1.data_o[85] ;
 wire \sub1.data_o[86] ;
 wire \sub1.data_o[87] ;
 wire \sub1.data_o[88] ;
 wire \sub1.data_o[89] ;
 wire \sub1.data_o[8] ;
 wire \sub1.data_o[90] ;
 wire \sub1.data_o[91] ;
 wire \sub1.data_o[92] ;
 wire \sub1.data_o[93] ;
 wire \sub1.data_o[94] ;
 wire \sub1.data_o[95] ;
 wire \sub1.data_o[96] ;
 wire \sub1.data_o[97] ;
 wire \sub1.data_o[98] ;
 wire \sub1.data_o[99] ;
 wire \sub1.data_o[9] ;
 wire \sub1.next_ready_o ;
 wire \sub1.ready_o ;
 wire \sub1.state[0] ;
 wire \sub1.state[1] ;
 wire \sub1.state[2] ;
 wire \sub1.state[3] ;
 wire \sub1.state[4] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1219_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(\mix1.data_o[84] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(\mix1.data_o[85] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(\mix1.data_o[85] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(\mix1.data_o[98] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_1516_));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_1683_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\mix1.data_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\mix1.data_o[99] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\sub1.data_o[52] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\sub1.data_o[71] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_1270_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net30));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__and2_1 _3844_ (.A(\mix1.state[1] ),
    .B(\mix1.state[0] ),
    .X(_0650_));
 sky130_fd_sc_hd__buf_4 _3845_ (.A(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__clkbuf_4 _3846_ (.A(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__clkbuf_4 _3847_ (.A(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__buf_4 _3848_ (.A(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__buf_4 _3849_ (.A(_0654_),
    .X(\mix1.next_ready_o ));
 sky130_fd_sc_hd__clkbuf_4 _3850_ (.A(\sub1.state[0] ),
    .X(_0655_));
 sky130_fd_sc_hd__clkbuf_4 _3851_ (.A(\sub1.state[1] ),
    .X(_0656_));
 sky130_fd_sc_hd__buf_4 _3852_ (.A(\sub1.state[3] ),
    .X(_0657_));
 sky130_fd_sc_hd__or4_4 _3853_ (.A(_0655_),
    .B(_0656_),
    .C(_0657_),
    .D(\sub1.state[2] ),
    .X(_0658_));
 sky130_fd_sc_hd__inv_2 _3854_ (.A(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__nand2_1 _3855_ (.A(\sub1.state[4] ),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__inv_2 _3856_ (.A(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__clkbuf_4 _3857_ (.A(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__buf_4 _3858_ (.A(_0662_),
    .X(\sub1.next_ready_o ));
 sky130_fd_sc_hd__xor2_2 _3859_ (.A(\addroundkey_round[3] ),
    .B(\round[3] ),
    .X(_0663_));
 sky130_fd_sc_hd__xor2_2 _3860_ (.A(\addroundkey_round[2] ),
    .B(\round[2] ),
    .X(_0664_));
 sky130_fd_sc_hd__clkbuf_4 _3861_ (.A(\round[1] ),
    .X(_0665_));
 sky130_fd_sc_hd__xor2_2 _3862_ (.A(\addroundkey_round[1] ),
    .B(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__buf_2 _3863_ (.A(\round[0] ),
    .X(_0667_));
 sky130_fd_sc_hd__xor2_2 _3864_ (.A(\addroundkey_round[0] ),
    .B(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__or4_1 _3865_ (.A(_0663_),
    .B(_0664_),
    .C(_0666_),
    .D(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__nand2b_2 _3866_ (.A_N(addroundkey_start_i),
    .B(\ks1.ready_o ),
    .Y(_0670_));
 sky130_fd_sc_hd__or3_1 _3867_ (.A(_0667_),
    .B(_0665_),
    .C(\round[2] ),
    .X(_0671_));
 sky130_fd_sc_hd__nor2_1 _3868_ (.A(\round[3] ),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__and2_1 _3869_ (.A(addroundkey_start_i),
    .B(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__buf_2 _3870_ (.A(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_8 _3871_ (.A(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__o21bai_2 _3872_ (.A1(_0669_),
    .A2(_0670_),
    .B1_N(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__clkbuf_8 _3873_ (.A(_0676_),
    .X(next_addroundkey_ready_o));
 sky130_fd_sc_hd__buf_4 _3874_ (.A(state),
    .X(_0677_));
 sky130_fd_sc_hd__buf_6 _3875_ (.A(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_4 _3876_ (.A(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__or4bb_2 _3877_ (.A(\round[0] ),
    .B(\round[2] ),
    .C_N(\round[3] ),
    .D_N(\round[1] ),
    .X(_0680_));
 sky130_fd_sc_hd__inv_2 _3878_ (.A(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__inv_4 _3879_ (.A(net129),
    .Y(_0682_));
 sky130_fd_sc_hd__mux2_4 _3880_ (.A0(_0672_),
    .A1(_0681_),
    .S(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__and3_2 _3881_ (.A(_0679_),
    .B(addroundkey_ready_o),
    .C(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_1 _3882_ (.A(_0684_),
    .X(next_ready_o));
 sky130_fd_sc_hd__or2_4 _3883_ (.A(\sub1.state[3] ),
    .B(\sub1.state[2] ),
    .X(_0685_));
 sky130_fd_sc_hd__nand2_2 _3884_ (.A(_0655_),
    .B(_0656_),
    .Y(_0686_));
 sky130_fd_sc_hd__nor2_4 _3885_ (.A(_0685_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__and2_1 _3886_ (.A(net129),
    .B(_0680_),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_4 _3887_ (.A(_0688_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _3888_ (.A0(net384),
    .A1(\mix1.data_o[97] ),
    .S(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__nand2b_2 _3889_ (.A_N(_0655_),
    .B(_0656_),
    .Y(_0691_));
 sky130_fd_sc_hd__nor2_4 _3890_ (.A(_0685_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__clkbuf_4 _3891_ (.A(_0689_),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _3892_ (.A0(net266),
    .A1(\mix1.data_o[105] ),
    .S(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__a22o_1 _3893_ (.A1(_0687_),
    .A2(_0690_),
    .B1(_0692_),
    .B2(_0694_),
    .X(_0695_));
 sky130_fd_sc_hd__or3b_2 _3894_ (.A(\sub1.state[0] ),
    .B(\sub1.state[1] ),
    .C_N(\sub1.state[3] ),
    .X(_0696_));
 sky130_fd_sc_hd__nor2_4 _3895_ (.A(\sub1.state[2] ),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__mux2_1 _3896_ (.A0(net340),
    .A1(\mix1.data_o[57] ),
    .S(_0689_),
    .X(_0698_));
 sky130_fd_sc_hd__inv_4 _3897_ (.A(\sub1.state[2] ),
    .Y(_0699_));
 sky130_fd_sc_hd__and4b_1 _3898_ (.A_N(_0656_),
    .B(_0657_),
    .C(_0699_),
    .D(_0655_),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _3899_ (.A0(net331),
    .A1(\mix1.data_o[49] ),
    .S(_0693_),
    .X(_0701_));
 sky130_fd_sc_hd__a22o_1 _3900_ (.A1(_0697_),
    .A2(_0698_),
    .B1(_0700_),
    .B2(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__and4b_2 _3901_ (.A_N(_0655_),
    .B(_0656_),
    .C(_0657_),
    .D(_0699_),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _3902_ (.A0(net323),
    .A1(\mix1.data_o[41] ),
    .S(_0689_),
    .X(_0704_));
 sky130_fd_sc_hd__or2b_2 _3903_ (.A(_0656_),
    .B_N(_0655_),
    .X(_0705_));
 sky130_fd_sc_hd__nor2_2 _3904_ (.A(_0685_),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__mux2_1 _3905_ (.A0(net275),
    .A1(\mix1.data_o[113] ),
    .S(_0689_),
    .X(_0707_));
 sky130_fd_sc_hd__a22o_1 _3906_ (.A1(_0703_),
    .A2(_0704_),
    .B1(_0706_),
    .B2(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__nor3_4 _3907_ (.A(_0657_),
    .B(_0699_),
    .C(_0686_),
    .Y(_0709_));
 sky130_fd_sc_hd__mux2_1 _3908_ (.A0(net349),
    .A1(\mix1.data_o[65] ),
    .S(_0689_),
    .X(_0710_));
 sky130_fd_sc_hd__and4_1 _3909_ (.A(\sub1.state[0] ),
    .B(\sub1.state[1] ),
    .C(\sub1.state[3] ),
    .D(\sub1.state[2] ),
    .X(_0711_));
 sky130_fd_sc_hd__buf_4 _3910_ (.A(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__nor2_4 _3911_ (.A(_0699_),
    .B(_0696_),
    .Y(_0713_));
 sky130_fd_sc_hd__a22o_1 _3912_ (.A1(net299),
    .A2(_0712_),
    .B1(_0713_),
    .B2(net305),
    .X(_0714_));
 sky130_fd_sc_hd__nand2_2 _3913_ (.A(net129),
    .B(_0680_),
    .Y(_0715_));
 sky130_fd_sc_hd__a22o_1 _3914_ (.A1(_0709_),
    .A2(_0710_),
    .B1(_0714_),
    .B2(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__or4_1 _3915_ (.A(_0695_),
    .B(_0702_),
    .C(_0708_),
    .D(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__a22oi_2 _3916_ (.A1(net129),
    .A2(\mix1.ready_o ),
    .B1(_0715_),
    .B2(addroundkey_ready_o),
    .Y(_0718_));
 sky130_fd_sc_hd__a21oi_4 _3917_ (.A1(state),
    .A2(_0683_),
    .B1(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__nor2_4 _3918_ (.A(\sub1.state[4] ),
    .B(_0658_),
    .Y(_0720_));
 sky130_fd_sc_hd__buf_4 _3919_ (.A(_0693_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _3920_ (.A0(net284),
    .A1(\mix1.data_o[121] ),
    .S(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__and3_1 _3921_ (.A(_0719_),
    .B(_0720_),
    .C(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__nor3_4 _3922_ (.A(_0657_),
    .B(_0699_),
    .C(_0705_),
    .Y(_0724_));
 sky130_fd_sc_hd__or2_1 _3923_ (.A(net367),
    .B(_0693_),
    .X(_0725_));
 sky130_fd_sc_hd__o211a_1 _3924_ (.A1(\mix1.data_o[81] ),
    .A2(_0715_),
    .B1(_0724_),
    .C1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__nor4_4 _3925_ (.A(_0655_),
    .B(_0656_),
    .C(_0657_),
    .D(_0699_),
    .Y(_0727_));
 sky130_fd_sc_hd__mux2_1 _3926_ (.A0(net375),
    .A1(\mix1.data_o[89] ),
    .S(_0689_),
    .X(_0728_));
 sky130_fd_sc_hd__and4_1 _3927_ (.A(_0655_),
    .B(_0656_),
    .C(_0657_),
    .D(_0699_),
    .X(_0729_));
 sky130_fd_sc_hd__clkbuf_4 _3928_ (.A(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _3929_ (.A0(net314),
    .A1(\mix1.data_o[33] ),
    .S(_0693_),
    .X(_0731_));
 sky130_fd_sc_hd__a22o_1 _3930_ (.A1(_0727_),
    .A2(_0728_),
    .B1(_0730_),
    .B2(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__and4b_1 _3931_ (.A_N(_0656_),
    .B(\sub1.state[3] ),
    .C(\sub1.state[2] ),
    .D(\sub1.state[0] ),
    .X(_0733_));
 sky130_fd_sc_hd__buf_2 _3932_ (.A(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__mux2_1 _3933_ (.A0(net296),
    .A1(\mix1.data_o[17] ),
    .S(_0689_),
    .X(_0735_));
 sky130_fd_sc_hd__a22o_1 _3934_ (.A1(\mix1.data_o[1] ),
    .A2(_0711_),
    .B1(_0713_),
    .B2(\mix1.data_o[25] ),
    .X(_0736_));
 sky130_fd_sc_hd__clkbuf_4 _3935_ (.A(_0689_),
    .X(_0737_));
 sky130_fd_sc_hd__buf_4 _3936_ (.A(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__a22o_1 _3937_ (.A1(_0734_),
    .A2(_0735_),
    .B1(_0736_),
    .B2(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__nor3_4 _3938_ (.A(_0657_),
    .B(_0699_),
    .C(_0691_),
    .Y(_0740_));
 sky130_fd_sc_hd__mux2_1 _3939_ (.A0(net358),
    .A1(\mix1.data_o[73] ),
    .S(_0693_),
    .X(_0741_));
 sky130_fd_sc_hd__and4b_1 _3940_ (.A_N(_0655_),
    .B(_0656_),
    .C(_0657_),
    .D(\sub1.state[2] ),
    .X(_0742_));
 sky130_fd_sc_hd__clkbuf_4 _3941_ (.A(_0742_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _3942_ (.A0(net387),
    .A1(\mix1.data_o[9] ),
    .S(_0693_),
    .X(_0744_));
 sky130_fd_sc_hd__a22o_1 _3943_ (.A1(_0740_),
    .A2(_0741_),
    .B1(_0743_),
    .B2(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__or4_1 _3944_ (.A(_0726_),
    .B(_0732_),
    .C(_0739_),
    .D(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__or4_4 _3945_ (.A(\round[0] ),
    .B(_0665_),
    .C(\round[2] ),
    .D(\round[3] ),
    .X(_0747_));
 sky130_fd_sc_hd__nand2_8 _3946_ (.A(addroundkey_start_i),
    .B(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__and2b_1 _3947_ (.A_N(addroundkey_start_i),
    .B(\ks1.ready_o ),
    .X(_0749_));
 sky130_fd_sc_hd__o41ai_4 _3948_ (.A1(_0663_),
    .A2(_0664_),
    .A3(_0666_),
    .A4(_0668_),
    .B1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__nand2_1 _3949_ (.A(_0748_),
    .B(net389),
    .Y(_0751_));
 sky130_fd_sc_hd__or3_2 _3950_ (.A(\ks1.state[2] ),
    .B(\ks1.state[1] ),
    .C(\ks1.state[0] ),
    .X(_0752_));
 sky130_fd_sc_hd__or3b_1 _3951_ (.A(\ks1.state[1] ),
    .B(\ks1.state[0] ),
    .C_N(\ks1.state[2] ),
    .X(_0753_));
 sky130_fd_sc_hd__buf_2 _3952_ (.A(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__a2bb2o_4 _3953_ (.A1_N(_0751_),
    .A2_N(_0752_),
    .B1(_0754_),
    .B2(\ks1.state[2] ),
    .X(_0755_));
 sky130_fd_sc_hd__o31a_1 _3954_ (.A1(_0717_),
    .A2(_0723_),
    .A3(_0746_),
    .B1(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__nor3b_4 _3955_ (.A(\ks1.state[2] ),
    .B(\ks1.state[0] ),
    .C_N(\ks1.state[1] ),
    .Y(_0757_));
 sky130_fd_sc_hd__nor3_1 _3956_ (.A(\addroundkey_round[1] ),
    .B(\addroundkey_round[3] ),
    .C(\addroundkey_round[2] ),
    .Y(_0758_));
 sky130_fd_sc_hd__and2_1 _3957_ (.A(addroundkey_start_i),
    .B(_0747_),
    .X(_0759_));
 sky130_fd_sc_hd__a21o_2 _3958_ (.A1(net389),
    .A2(_0758_),
    .B1(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__buf_4 _3959_ (.A(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _3960_ (.A0(\ks1.key_reg[9] ),
    .A1(net257),
    .S(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__nor3b_4 _3961_ (.A(\ks1.state[2] ),
    .B(\ks1.state[1] ),
    .C_N(\ks1.state[0] ),
    .Y(_0763_));
 sky130_fd_sc_hd__mux2_2 _3962_ (.A0(\ks1.key_reg[17] ),
    .A1(net166),
    .S(_0761_),
    .X(_0764_));
 sky130_fd_sc_hd__and3b_1 _3963_ (.A_N(\ks1.state[2] ),
    .B(\ks1.state[1] ),
    .C(\ks1.state[0] ),
    .X(_0765_));
 sky130_fd_sc_hd__buf_2 _3964_ (.A(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__buf_4 _3965_ (.A(_0760_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _3966_ (.A0(\ks1.key_reg[1] ),
    .A1(net169),
    .S(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__a21oi_4 _3967_ (.A1(_0748_),
    .A2(net389),
    .B1(_0752_),
    .Y(_0769_));
 sky130_fd_sc_hd__mux2_1 _3968_ (.A0(\ks1.key_reg[25] ),
    .A1(net175),
    .S(_0767_),
    .X(_0770_));
 sky130_fd_sc_hd__a22o_1 _3969_ (.A1(_0766_),
    .A2(_0768_),
    .B1(_0769_),
    .B2(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__a221o_1 _3970_ (.A1(_0757_),
    .A2(_0762_),
    .B1(_0763_),
    .B2(_0764_),
    .C1(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__or2_2 _3971_ (.A(_0756_),
    .B(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__clkbuf_4 _3972_ (.A(_0689_),
    .X(_0774_));
 sky130_fd_sc_hd__buf_4 _3973_ (.A(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _3974_ (.A0(net355),
    .A1(\mix1.data_o[70] ),
    .S(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__buf_4 _3975_ (.A(_0774_),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _3976_ (.A0(net372),
    .A1(\mix1.data_o[86] ),
    .S(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__a22o_1 _3977_ (.A1(_0709_),
    .A2(_0776_),
    .B1(_0778_),
    .B2(_0724_),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_1 _3978_ (.A0(net354),
    .A1(\mix1.data_o[6] ),
    .S(_0775_),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_1 _3979_ (.A0(net381),
    .A1(\mix1.data_o[94] ),
    .S(_0777_),
    .X(_0781_));
 sky130_fd_sc_hd__a22o_1 _3980_ (.A1(_0712_),
    .A2(_0780_),
    .B1(_0781_),
    .B2(_0727_),
    .X(_0782_));
 sky130_fd_sc_hd__mux2_1 _3981_ (.A0(net363),
    .A1(\mix1.data_o[78] ),
    .S(_0738_),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _3982_ (.A0(net311),
    .A1(\mix1.data_o[30] ),
    .S(_0777_),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_1 _3983_ (.A1(_0740_),
    .A2(_0783_),
    .B1(_0784_),
    .B2(_0713_),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _3984_ (.A0(net280),
    .A1(\mix1.data_o[118] ),
    .S(_0775_),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _3985_ (.A0(net293),
    .A1(\mix1.data_o[14] ),
    .S(_0777_),
    .X(_0787_));
 sky130_fd_sc_hd__a22o_1 _3986_ (.A1(_0706_),
    .A2(_0786_),
    .B1(_0787_),
    .B2(_0743_),
    .X(_0788_));
 sky130_fd_sc_hd__or4_2 _3987_ (.A(_0779_),
    .B(_0782_),
    .C(_0785_),
    .D(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _3988_ (.A0(net289),
    .A1(\mix1.data_o[126] ),
    .S(_0775_),
    .X(_0790_));
 sky130_fd_sc_hd__o2bb2a_2 _3989_ (.A1_N(\ks1.state[2] ),
    .A2_N(_0754_),
    .B1(_0752_),
    .B2(_0751_),
    .X(_0791_));
 sky130_fd_sc_hd__a31o_1 _3990_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0790_),
    .B1(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _3991_ (.A0(net263),
    .A1(\mix1.data_o[102] ),
    .S(_0738_),
    .X(_0793_));
 sky130_fd_sc_hd__clkbuf_4 _3992_ (.A(_0700_),
    .X(_0794_));
 sky130_fd_sc_hd__clkbuf_4 _3993_ (.A(_0703_),
    .X(_0795_));
 sky130_fd_sc_hd__a22o_1 _3994_ (.A1(net337),
    .A2(_0794_),
    .B1(_0795_),
    .B2(net328),
    .X(_0796_));
 sky130_fd_sc_hd__clkbuf_4 _3995_ (.A(_0715_),
    .X(_0797_));
 sky130_fd_sc_hd__buf_4 _3996_ (.A(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__or2_1 _3997_ (.A(net346),
    .B(_0721_),
    .X(_0799_));
 sky130_fd_sc_hd__o211a_1 _3998_ (.A1(\mix1.data_o[62] ),
    .A2(_0797_),
    .B1(_0697_),
    .C1(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__a221o_1 _3999_ (.A1(_0687_),
    .A2(_0793_),
    .B1(_0796_),
    .B2(_0798_),
    .C1(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__mux2_1 _4000_ (.A0(net272),
    .A1(\mix1.data_o[110] ),
    .S(_0775_),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_1 _4001_ (.A0(net319),
    .A1(\mix1.data_o[38] ),
    .S(_0777_),
    .X(_0803_));
 sky130_fd_sc_hd__a22o_1 _4002_ (.A1(_0692_),
    .A2(_0802_),
    .B1(_0803_),
    .B2(_0730_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _4003_ (.A0(net302),
    .A1(\mix1.data_o[22] ),
    .S(_0775_),
    .X(_0805_));
 sky130_fd_sc_hd__a22o_1 _4004_ (.A1(\mix1.data_o[54] ),
    .A2(_0794_),
    .B1(_0795_),
    .B2(\mix1.data_o[46] ),
    .X(_0806_));
 sky130_fd_sc_hd__clkbuf_4 _4005_ (.A(_0738_),
    .X(_0807_));
 sky130_fd_sc_hd__a22o_1 _4006_ (.A1(_0734_),
    .A2(_0805_),
    .B1(_0806_),
    .B2(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__or4_2 _4007_ (.A(_0792_),
    .B(_0801_),
    .C(_0804_),
    .D(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__clkbuf_8 _4008_ (.A(_0761_),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _4009_ (.A0(\ks1.key_reg[22] ),
    .A1(net172),
    .S(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _4010_ (.A0(\ks1.key_reg[6] ),
    .A1(net224),
    .S(_0761_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _4011_ (.A0(\ks1.key_reg[14] ),
    .A1(net163),
    .S(_0761_),
    .X(_0813_));
 sky130_fd_sc_hd__a22o_1 _4012_ (.A1(_0766_),
    .A2(_0812_),
    .B1(_0813_),
    .B2(_0757_),
    .X(_0814_));
 sky130_fd_sc_hd__buf_4 _4013_ (.A(_0767_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(\ks1.key_reg[30] ),
    .A1(net181),
    .S(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__a21o_1 _4015_ (.A1(_0769_),
    .A2(_0816_),
    .B1(_0755_),
    .X(_0817_));
 sky130_fd_sc_hd__a211o_2 _4016_ (.A1(_0763_),
    .A2(_0811_),
    .B1(_0814_),
    .C1(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__o21ai_4 _4017_ (.A1(_0789_),
    .A2(_0809_),
    .B1(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__mux2_1 _4018_ (.A0(net360),
    .A1(\mix1.data_o[75] ),
    .S(_0737_),
    .X(_0820_));
 sky130_fd_sc_hd__mux2_1 _4019_ (.A0(net378),
    .A1(\mix1.data_o[91] ),
    .S(_0774_),
    .X(_0821_));
 sky130_fd_sc_hd__a22o_1 _4020_ (.A1(_0740_),
    .A2(_0820_),
    .B1(_0821_),
    .B2(_0727_),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _4021_ (.A0(net316),
    .A1(\mix1.data_o[35] ),
    .S(_0737_),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _4022_ (.A0(net325),
    .A1(\mix1.data_o[43] ),
    .S(_0774_),
    .X(_0824_));
 sky130_fd_sc_hd__a22o_1 _4023_ (.A1(_0730_),
    .A2(_0823_),
    .B1(_0824_),
    .B2(_0795_),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_1 _4024_ (.A0(net342),
    .A1(\mix1.data_o[59] ),
    .S(_0737_),
    .X(_0826_));
 sky130_fd_sc_hd__mux2_1 _4025_ (.A0(net277),
    .A1(\mix1.data_o[115] ),
    .S(_0774_),
    .X(_0827_));
 sky130_fd_sc_hd__a22o_1 _4026_ (.A1(_0697_),
    .A2(_0826_),
    .B1(_0827_),
    .B2(_0706_),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(net351),
    .A1(\mix1.data_o[67] ),
    .S(_0737_),
    .X(_0829_));
 sky130_fd_sc_hd__a22o_1 _4028_ (.A1(net369),
    .A2(_0724_),
    .B1(_0734_),
    .B2(net298),
    .X(_0830_));
 sky130_fd_sc_hd__a22o_1 _4029_ (.A1(_0709_),
    .A2(_0829_),
    .B1(_0830_),
    .B2(_0797_),
    .X(_0831_));
 sky130_fd_sc_hd__or4_1 _4030_ (.A(_0822_),
    .B(_0825_),
    .C(_0828_),
    .D(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__buf_4 _4031_ (.A(_0693_),
    .X(_0833_));
 sky130_fd_sc_hd__buf_4 _4032_ (.A(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__mux2_1 _4033_ (.A0(net286),
    .A1(\mix1.data_o[123] ),
    .S(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__and3_1 _4034_ (.A(_0719_),
    .B(_0720_),
    .C(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__or2_1 _4035_ (.A(net334),
    .B(_0833_),
    .X(_0837_));
 sky130_fd_sc_hd__o211a_1 _4036_ (.A1(\mix1.data_o[51] ),
    .A2(_0797_),
    .B1(_0794_),
    .C1(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__mux2_1 _4037_ (.A0(net282),
    .A1(\mix1.data_o[11] ),
    .S(_0737_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _4038_ (.A0(net307),
    .A1(\mix1.data_o[27] ),
    .S(_0774_),
    .X(_0840_));
 sky130_fd_sc_hd__a22o_1 _4039_ (.A1(_0743_),
    .A2(_0839_),
    .B1(_0840_),
    .B2(_0713_),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _4040_ (.A0(net386),
    .A1(\mix1.data_o[99] ),
    .S(_0737_),
    .X(_0842_));
 sky130_fd_sc_hd__a22o_1 _4041_ (.A1(\mix1.data_o[83] ),
    .A2(_0724_),
    .B1(_0734_),
    .B2(\mix1.data_o[19] ),
    .X(_0843_));
 sky130_fd_sc_hd__a22o_1 _4042_ (.A1(_0687_),
    .A2(_0842_),
    .B1(_0843_),
    .B2(_0834_),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_1 _4043_ (.A0(net268),
    .A1(\mix1.data_o[107] ),
    .S(_0774_),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _4044_ (.A0(net321),
    .A1(\mix1.data_o[3] ),
    .S(_0774_),
    .X(_0846_));
 sky130_fd_sc_hd__a22o_1 _4045_ (.A1(_0692_),
    .A2(_0845_),
    .B1(_0846_),
    .B2(_0712_),
    .X(_0847_));
 sky130_fd_sc_hd__or4_1 _4046_ (.A(_0838_),
    .B(_0841_),
    .C(_0844_),
    .D(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__o31a_1 _4047_ (.A1(_0832_),
    .A2(_0836_),
    .A3(_0848_),
    .B1(_0755_),
    .X(_0849_));
 sky130_fd_sc_hd__buf_4 _4048_ (.A(_0757_),
    .X(_0850_));
 sky130_fd_sc_hd__mux2_1 _4049_ (.A0(\ks1.key_reg[11] ),
    .A1(net152),
    .S(_0815_),
    .X(_0851_));
 sky130_fd_sc_hd__mux2_1 _4050_ (.A0(\ks1.key_reg[19] ),
    .A1(net168),
    .S(_0810_),
    .X(_0852_));
 sky130_fd_sc_hd__mux2_1 _4051_ (.A0(\ks1.key_reg[3] ),
    .A1(net191),
    .S(_0761_),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _4052_ (.A0(\ks1.key_reg[27] ),
    .A1(net177),
    .S(_0761_),
    .X(_0854_));
 sky130_fd_sc_hd__a22o_1 _4053_ (.A1(_0766_),
    .A2(_0853_),
    .B1(_0854_),
    .B2(_0769_),
    .X(_0855_));
 sky130_fd_sc_hd__a221o_2 _4054_ (.A1(_0850_),
    .A2(_0851_),
    .B1(_0852_),
    .B2(_0763_),
    .C1(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__or2_4 _4055_ (.A(_0849_),
    .B(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__xor2_2 _4056_ (.A(_0819_),
    .B(_0857_),
    .X(_0858_));
 sky130_fd_sc_hd__xor2_1 _4057_ (.A(_0773_),
    .B(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__buf_4 _4058_ (.A(_0693_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _4059_ (.A0(net352),
    .A1(\mix1.data_o[68] ),
    .S(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__buf_4 _4060_ (.A(_0693_),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _4061_ (.A0(net370),
    .A1(\mix1.data_o[84] ),
    .S(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__a22o_1 _4062_ (.A1(_0709_),
    .A2(_0861_),
    .B1(_0863_),
    .B2(_0724_),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _4063_ (.A0(net332),
    .A1(\mix1.data_o[4] ),
    .S(_0860_),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _4064_ (.A0(net379),
    .A1(\mix1.data_o[92] ),
    .S(_0862_),
    .X(_0866_));
 sky130_fd_sc_hd__a22o_1 _4065_ (.A1(_0712_),
    .A2(_0865_),
    .B1(_0866_),
    .B2(_0727_),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _4066_ (.A0(net361),
    .A1(\mix1.data_o[76] ),
    .S(_0860_),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _4067_ (.A0(net308),
    .A1(\mix1.data_o[28] ),
    .S(_0862_),
    .X(_0869_));
 sky130_fd_sc_hd__a22o_1 _4068_ (.A1(_0740_),
    .A2(_0868_),
    .B1(_0869_),
    .B2(_0713_),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(net278),
    .A1(\mix1.data_o[116] ),
    .S(_0860_),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _4070_ (.A0(net291),
    .A1(\mix1.data_o[12] ),
    .S(_0862_),
    .X(_0872_));
 sky130_fd_sc_hd__a22o_1 _4071_ (.A1(_0706_),
    .A2(_0871_),
    .B1(_0872_),
    .B2(_0743_),
    .X(_0873_));
 sky130_fd_sc_hd__or4_1 _4072_ (.A(_0864_),
    .B(_0867_),
    .C(_0870_),
    .D(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _4073_ (.A0(net287),
    .A1(\mix1.data_o[124] ),
    .S(_0721_),
    .X(_0875_));
 sky130_fd_sc_hd__a31o_1 _4074_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0875_),
    .B1(_0791_),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(net261),
    .A1(\mix1.data_o[100] ),
    .S(_0774_),
    .X(_0877_));
 sky130_fd_sc_hd__a22o_1 _4076_ (.A1(net335),
    .A2(_0700_),
    .B1(_0703_),
    .B2(net326),
    .X(_0878_));
 sky130_fd_sc_hd__buf_4 _4077_ (.A(_0715_),
    .X(_0879_));
 sky130_fd_sc_hd__or2_1 _4078_ (.A(net344),
    .B(_0737_),
    .X(_0880_));
 sky130_fd_sc_hd__o211a_1 _4079_ (.A1(\mix1.data_o[60] ),
    .A2(_0879_),
    .B1(_0697_),
    .C1(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__a221o_1 _4080_ (.A1(_0687_),
    .A2(_0877_),
    .B1(_0878_),
    .B2(_0797_),
    .C1(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(net269),
    .A1(\mix1.data_o[108] ),
    .S(_0833_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _4082_ (.A0(net317),
    .A1(\mix1.data_o[36] ),
    .S(_0862_),
    .X(_0884_));
 sky130_fd_sc_hd__a22o_1 _4083_ (.A1(_0692_),
    .A2(_0883_),
    .B1(_0884_),
    .B2(_0730_),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _4084_ (.A0(net300),
    .A1(\mix1.data_o[20] ),
    .S(_0860_),
    .X(_0886_));
 sky130_fd_sc_hd__a22o_1 _4085_ (.A1(\mix1.data_o[52] ),
    .A2(_0794_),
    .B1(_0795_),
    .B2(\mix1.data_o[44] ),
    .X(_0887_));
 sky130_fd_sc_hd__a22o_1 _4086_ (.A1(_0734_),
    .A2(_0886_),
    .B1(_0887_),
    .B2(_0807_),
    .X(_0888_));
 sky130_fd_sc_hd__or4_1 _4087_ (.A(_0876_),
    .B(_0882_),
    .C(_0885_),
    .D(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__mux2_1 _4088_ (.A0(\ks1.key_reg[4] ),
    .A1(net202),
    .S(_0815_),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_2 _4089_ (.A0(\ks1.key_reg[20] ),
    .A1(net170),
    .S(_0767_),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _4090_ (.A0(\ks1.key_reg[12] ),
    .A1(net161),
    .S(_0767_),
    .X(_0892_));
 sky130_fd_sc_hd__a22o_1 _4091_ (.A1(_0763_),
    .A2(_0891_),
    .B1(_0892_),
    .B2(_0757_),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _4092_ (.A0(\ks1.key_reg[28] ),
    .A1(net178),
    .S(_0761_),
    .X(_0894_));
 sky130_fd_sc_hd__a21o_1 _4093_ (.A1(_0769_),
    .A2(_0894_),
    .B1(_0755_),
    .X(_0895_));
 sky130_fd_sc_hd__a211o_1 _4094_ (.A1(_0766_),
    .A2(_0890_),
    .B1(_0893_),
    .C1(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__o21a_1 _4095_ (.A1(_0874_),
    .A2(_0889_),
    .B1(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__inv_2 _4096_ (.A(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_4 _4097_ (.A(net129),
    .B(_0755_),
    .Y(_0899_));
 sky130_fd_sc_hd__mux2_4 _4098_ (.A0(_0859_),
    .A1(_0898_),
    .S(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _4099_ (.A0(net348),
    .A1(\mix1.data_o[64] ),
    .S(_0775_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _4100_ (.A0(\mix1.data_o[80] ),
    .A1(net366),
    .S(_0879_),
    .X(_0902_));
 sky130_fd_sc_hd__buf_4 _4101_ (.A(_0724_),
    .X(_0903_));
 sky130_fd_sc_hd__a22o_1 _4102_ (.A1(_0709_),
    .A2(_0901_),
    .B1(_0902_),
    .B2(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _4103_ (.A0(net260),
    .A1(\mix1.data_o[0] ),
    .S(_0775_),
    .X(_0905_));
 sky130_fd_sc_hd__mux2_1 _4104_ (.A0(\mix1.data_o[88] ),
    .A1(net374),
    .S(_0879_),
    .X(_0906_));
 sky130_fd_sc_hd__a22o_1 _4105_ (.A1(_0712_),
    .A2(_0905_),
    .B1(_0906_),
    .B2(_0727_),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _4106_ (.A0(net357),
    .A1(\mix1.data_o[72] ),
    .S(_0775_),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _4107_ (.A0(\mix1.data_o[24] ),
    .A1(net304),
    .S(_0879_),
    .X(_0909_));
 sky130_fd_sc_hd__a22o_1 _4108_ (.A1(_0740_),
    .A2(_0908_),
    .B1(_0909_),
    .B2(_0713_),
    .X(_0910_));
 sky130_fd_sc_hd__buf_4 _4109_ (.A(_0706_),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _4110_ (.A0(\mix1.data_o[112] ),
    .A1(net274),
    .S(_0879_),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _4111_ (.A0(\mix1.data_o[8] ),
    .A1(net376),
    .S(_0797_),
    .X(_0913_));
 sky130_fd_sc_hd__a22o_1 _4112_ (.A1(_0911_),
    .A2(_0912_),
    .B1(_0913_),
    .B2(_0743_),
    .X(_0914_));
 sky130_fd_sc_hd__or4_2 _4113_ (.A(_0904_),
    .B(_0907_),
    .C(_0910_),
    .D(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(\mix1.data_o[120] ),
    .A1(net283),
    .S(_0879_),
    .X(_0916_));
 sky130_fd_sc_hd__a31o_1 _4115_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0916_),
    .B1(_0791_),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _4116_ (.A0(net383),
    .A1(\mix1.data_o[96] ),
    .S(_0738_),
    .X(_0918_));
 sky130_fd_sc_hd__a22o_1 _4117_ (.A1(net330),
    .A2(_0794_),
    .B1(_0795_),
    .B2(net322),
    .X(_0919_));
 sky130_fd_sc_hd__or2_1 _4118_ (.A(net339),
    .B(_0862_),
    .X(_0920_));
 sky130_fd_sc_hd__o211a_1 _4119_ (.A1(\mix1.data_o[56] ),
    .A2(_0797_),
    .B1(_0697_),
    .C1(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__a221o_1 _4120_ (.A1(_0687_),
    .A2(_0918_),
    .B1(_0919_),
    .B2(_0798_),
    .C1(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__clkbuf_8 _4121_ (.A(_0692_),
    .X(_0923_));
 sky130_fd_sc_hd__mux2_1 _4122_ (.A0(\mix1.data_o[104] ),
    .A1(net265),
    .S(_0879_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _4123_ (.A0(net313),
    .A1(\mix1.data_o[32] ),
    .S(_0834_),
    .X(_0925_));
 sky130_fd_sc_hd__a22o_1 _4124_ (.A1(_0923_),
    .A2(_0924_),
    .B1(_0925_),
    .B2(_0730_),
    .X(_0926_));
 sky130_fd_sc_hd__buf_4 _4125_ (.A(_0734_),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _4126_ (.A0(\mix1.data_o[16] ),
    .A1(net295),
    .S(_0879_),
    .X(_0928_));
 sky130_fd_sc_hd__buf_4 _4127_ (.A(_0794_),
    .X(_0929_));
 sky130_fd_sc_hd__a22o_1 _4128_ (.A1(\mix1.data_o[48] ),
    .A2(_0929_),
    .B1(_0795_),
    .B2(\mix1.data_o[40] ),
    .X(_0930_));
 sky130_fd_sc_hd__a22o_1 _4129_ (.A1(_0927_),
    .A2(_0928_),
    .B1(_0930_),
    .B2(_0807_),
    .X(_0931_));
 sky130_fd_sc_hd__or4_1 _4130_ (.A(_0917_),
    .B(_0922_),
    .C(_0926_),
    .D(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_1 _4131_ (.A0(\ks1.key_reg[16] ),
    .A1(net165),
    .S(_0810_),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _4132_ (.A0(\ks1.key_reg[0] ),
    .A1(net130),
    .S(_0761_),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _4133_ (.A0(\ks1.key_reg[8] ),
    .A1(net246),
    .S(_0815_),
    .X(_0935_));
 sky130_fd_sc_hd__a22o_1 _4134_ (.A1(_0766_),
    .A2(_0934_),
    .B1(_0935_),
    .B2(_0757_),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _4135_ (.A0(\ks1.key_reg[24] ),
    .A1(net174),
    .S(_0815_),
    .X(_0937_));
 sky130_fd_sc_hd__a21o_1 _4136_ (.A1(_0769_),
    .A2(_0937_),
    .B1(_0755_),
    .X(_0938_));
 sky130_fd_sc_hd__a211o_2 _4137_ (.A1(_0763_),
    .A2(_0933_),
    .B1(_0936_),
    .C1(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__o21ai_4 _4138_ (.A1(_0915_),
    .A2(_0932_),
    .B1(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__mux2_1 _4139_ (.A0(net353),
    .A1(\mix1.data_o[69] ),
    .S(_0777_),
    .X(_0941_));
 sky130_fd_sc_hd__mux2_1 _4140_ (.A0(net371),
    .A1(\mix1.data_o[85] ),
    .S(_0834_),
    .X(_0942_));
 sky130_fd_sc_hd__a22o_1 _4141_ (.A1(_0709_),
    .A2(_0941_),
    .B1(_0942_),
    .B2(_0903_),
    .X(_0943_));
 sky130_fd_sc_hd__mux2_1 _4142_ (.A0(net343),
    .A1(\mix1.data_o[5] ),
    .S(_0777_),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_1 _4143_ (.A0(net380),
    .A1(\mix1.data_o[93] ),
    .S(_0834_),
    .X(_0945_));
 sky130_fd_sc_hd__a22o_1 _4144_ (.A1(_0712_),
    .A2(_0944_),
    .B1(_0945_),
    .B2(_0727_),
    .X(_0946_));
 sky130_fd_sc_hd__clkbuf_8 _4145_ (.A(_0740_),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _4146_ (.A0(net362),
    .A1(\mix1.data_o[77] ),
    .S(_0775_),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _4147_ (.A0(net309),
    .A1(\mix1.data_o[29] ),
    .S(_0834_),
    .X(_0949_));
 sky130_fd_sc_hd__a22o_1 _4148_ (.A1(_0947_),
    .A2(_0948_),
    .B1(_0949_),
    .B2(_0713_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _4149_ (.A0(net279),
    .A1(\mix1.data_o[117] ),
    .S(_0777_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _4150_ (.A0(net292),
    .A1(\mix1.data_o[13] ),
    .S(_0834_),
    .X(_0952_));
 sky130_fd_sc_hd__clkbuf_4 _4151_ (.A(_0743_),
    .X(_0953_));
 sky130_fd_sc_hd__a22o_1 _4152_ (.A1(_0911_),
    .A2(_0951_),
    .B1(_0952_),
    .B2(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__or4_2 _4153_ (.A(_0943_),
    .B(_0946_),
    .C(_0950_),
    .D(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _4154_ (.A0(net288),
    .A1(\mix1.data_o[125] ),
    .S(_0834_),
    .X(_0956_));
 sky130_fd_sc_hd__a31o_1 _4155_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_0956_),
    .B1(_0791_),
    .X(_0957_));
 sky130_fd_sc_hd__clkbuf_4 _4156_ (.A(_0687_),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _4157_ (.A0(net262),
    .A1(\mix1.data_o[101] ),
    .S(_0738_),
    .X(_0959_));
 sky130_fd_sc_hd__a22o_1 _4158_ (.A1(net336),
    .A2(_0794_),
    .B1(_0795_),
    .B2(net327),
    .X(_0960_));
 sky130_fd_sc_hd__clkbuf_4 _4159_ (.A(_0697_),
    .X(_0961_));
 sky130_fd_sc_hd__or2_1 _4160_ (.A(net345),
    .B(_0862_),
    .X(_0962_));
 sky130_fd_sc_hd__o211a_1 _4161_ (.A1(\mix1.data_o[61] ),
    .A2(_0797_),
    .B1(_0961_),
    .C1(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__a221o_1 _4162_ (.A1(_0958_),
    .A2(_0959_),
    .B1(_0960_),
    .B2(_0798_),
    .C1(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _4163_ (.A0(net270),
    .A1(\mix1.data_o[109] ),
    .S(_0777_),
    .X(_0965_));
 sky130_fd_sc_hd__mux2_1 _4164_ (.A0(net318),
    .A1(\mix1.data_o[37] ),
    .S(_0834_),
    .X(_0966_));
 sky130_fd_sc_hd__clkbuf_4 _4165_ (.A(_0730_),
    .X(_0967_));
 sky130_fd_sc_hd__a22o_1 _4166_ (.A1(_0923_),
    .A2(_0965_),
    .B1(_0966_),
    .B2(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _4167_ (.A0(net301),
    .A1(\mix1.data_o[21] ),
    .S(_0777_),
    .X(_0969_));
 sky130_fd_sc_hd__buf_4 _4168_ (.A(_0795_),
    .X(_0970_));
 sky130_fd_sc_hd__a22o_1 _4169_ (.A1(\mix1.data_o[53] ),
    .A2(_0929_),
    .B1(_0970_),
    .B2(\mix1.data_o[45] ),
    .X(_0971_));
 sky130_fd_sc_hd__a22o_1 _4170_ (.A1(_0927_),
    .A2(_0969_),
    .B1(_0971_),
    .B2(_0807_),
    .X(_0972_));
 sky130_fd_sc_hd__or4_2 _4171_ (.A(_0957_),
    .B(_0964_),
    .C(_0968_),
    .D(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__clkbuf_8 _4172_ (.A(_0763_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _4173_ (.A0(\ks1.key_reg[21] ),
    .A1(net171),
    .S(_0810_),
    .X(_0975_));
 sky130_fd_sc_hd__mux2_1 _4174_ (.A0(\ks1.key_reg[13] ),
    .A1(net162),
    .S(_0815_),
    .X(_0976_));
 sky130_fd_sc_hd__mux2_1 _4175_ (.A0(\ks1.key_reg[5] ),
    .A1(net213),
    .S(_0815_),
    .X(_0977_));
 sky130_fd_sc_hd__a22o_1 _4176_ (.A1(_0757_),
    .A2(_0976_),
    .B1(_0977_),
    .B2(_0766_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _4177_ (.A0(\ks1.key_reg[29] ),
    .A1(net179),
    .S(_0815_),
    .X(_0979_));
 sky130_fd_sc_hd__a21o_1 _4178_ (.A1(_0769_),
    .A2(_0979_),
    .B1(_0755_),
    .X(_0980_));
 sky130_fd_sc_hd__a211o_2 _4179_ (.A1(_0974_),
    .A2(_0975_),
    .B1(_0978_),
    .C1(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__o21ai_4 _4180_ (.A1(_0955_),
    .A2(_0973_),
    .B1(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__xor2_2 _4181_ (.A(_0940_),
    .B(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__xnor2_1 _4182_ (.A(_0857_),
    .B(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__mux2_2 _4183_ (.A0(_0984_),
    .A1(_0819_),
    .S(_0899_),
    .X(_0985_));
 sky130_fd_sc_hd__xor2_4 _4184_ (.A(_0900_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__xnor2_1 _4185_ (.A(_0773_),
    .B(_0897_),
    .Y(_0987_));
 sky130_fd_sc_hd__nor2_1 _4186_ (.A(_0819_),
    .B(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__and2_1 _4187_ (.A(_0819_),
    .B(_0987_),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _4188_ (.A0(net356),
    .A1(\mix1.data_o[71] ),
    .S(_0833_),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_2 _4189_ (.A0(net373),
    .A1(\mix1.data_o[87] ),
    .S(_0721_),
    .X(_0991_));
 sky130_fd_sc_hd__a22o_1 _4190_ (.A1(_0709_),
    .A2(_0990_),
    .B1(_0991_),
    .B2(_0724_),
    .X(_0992_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(net365),
    .A1(\mix1.data_o[7] ),
    .S(_0833_),
    .X(_0993_));
 sky130_fd_sc_hd__mux2_1 _4192_ (.A0(net382),
    .A1(\mix1.data_o[95] ),
    .S(_0721_),
    .X(_0994_));
 sky130_fd_sc_hd__a22o_1 _4193_ (.A1(_0712_),
    .A2(_0993_),
    .B1(_0994_),
    .B2(_0727_),
    .X(_0995_));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(net364),
    .A1(\mix1.data_o[79] ),
    .S(_0833_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _4195_ (.A0(net312),
    .A1(\mix1.data_o[31] ),
    .S(_0860_),
    .X(_0997_));
 sky130_fd_sc_hd__a22o_1 _4196_ (.A1(_0740_),
    .A2(_0996_),
    .B1(_0997_),
    .B2(_0713_),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_1 _4197_ (.A0(net281),
    .A1(\mix1.data_o[119] ),
    .S(_0833_),
    .X(_0999_));
 sky130_fd_sc_hd__mux2_1 _4198_ (.A0(net294),
    .A1(\mix1.data_o[15] ),
    .S(_0721_),
    .X(_1000_));
 sky130_fd_sc_hd__a22o_1 _4199_ (.A1(_0706_),
    .A2(_0999_),
    .B1(_1000_),
    .B2(_0743_),
    .X(_1001_));
 sky130_fd_sc_hd__or4_1 _4200_ (.A(_0992_),
    .B(_0995_),
    .C(_0998_),
    .D(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _4201_ (.A0(net290),
    .A1(\mix1.data_o[127] ),
    .S(_0860_),
    .X(_1003_));
 sky130_fd_sc_hd__a31o_1 _4202_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_1003_),
    .B1(_0791_),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _4203_ (.A0(net264),
    .A1(\mix1.data_o[103] ),
    .S(_0774_),
    .X(_1005_));
 sky130_fd_sc_hd__a22o_1 _4204_ (.A1(net338),
    .A2(_0700_),
    .B1(_0703_),
    .B2(net329),
    .X(_1006_));
 sky130_fd_sc_hd__or2_1 _4205_ (.A(net347),
    .B(_0737_),
    .X(_1007_));
 sky130_fd_sc_hd__o211a_1 _4206_ (.A1(\mix1.data_o[63] ),
    .A2(_0879_),
    .B1(_0697_),
    .C1(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__a221o_1 _4207_ (.A1(_0687_),
    .A2(_1005_),
    .B1(_1006_),
    .B2(_0797_),
    .C1(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _4208_ (.A0(net273),
    .A1(\mix1.data_o[111] ),
    .S(_0833_),
    .X(_1010_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(net320),
    .A1(\mix1.data_o[39] ),
    .S(_0860_),
    .X(_1011_));
 sky130_fd_sc_hd__a22o_1 _4210_ (.A1(_0692_),
    .A2(_1010_),
    .B1(_1011_),
    .B2(_0730_),
    .X(_1012_));
 sky130_fd_sc_hd__mux2_1 _4211_ (.A0(net303),
    .A1(\mix1.data_o[23] ),
    .S(_0833_),
    .X(_1013_));
 sky130_fd_sc_hd__a22o_1 _4212_ (.A1(\mix1.data_o[55] ),
    .A2(_0794_),
    .B1(_0795_),
    .B2(\mix1.data_o[47] ),
    .X(_1014_));
 sky130_fd_sc_hd__a22o_1 _4213_ (.A1(_0734_),
    .A2(_1013_),
    .B1(_1014_),
    .B2(_0834_),
    .X(_1015_));
 sky130_fd_sc_hd__or4_1 _4214_ (.A(_1004_),
    .B(_1009_),
    .C(_1012_),
    .D(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__mux2_1 _4215_ (.A0(\ks1.key_reg[7] ),
    .A1(net235),
    .S(_0815_),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _4216_ (.A0(\ks1.key_reg[23] ),
    .A1(net173),
    .S(_0767_),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _4217_ (.A0(\ks1.key_reg[15] ),
    .A1(net164),
    .S(_0767_),
    .X(_1019_));
 sky130_fd_sc_hd__a22o_1 _4218_ (.A1(_0763_),
    .A2(_1018_),
    .B1(_1019_),
    .B2(_0757_),
    .X(_1020_));
 sky130_fd_sc_hd__mux2_1 _4219_ (.A0(\ks1.key_reg[31] ),
    .A1(net182),
    .S(_0767_),
    .X(_1021_));
 sky130_fd_sc_hd__a21o_1 _4220_ (.A1(_0769_),
    .A2(_1021_),
    .B1(_0755_),
    .X(_1022_));
 sky130_fd_sc_hd__a211o_2 _4221_ (.A1(_0766_),
    .A2(_1017_),
    .B1(_1020_),
    .C1(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__o21a_2 _4222_ (.A1(_1002_),
    .A2(_1016_),
    .B1(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__nand2_1 _4223_ (.A(_0899_),
    .B(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__o31a_4 _4224_ (.A1(_0899_),
    .A2(_0988_),
    .A3(_0989_),
    .B1(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__xor2_1 _4225_ (.A(_0858_),
    .B(_0940_),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_4 _4226_ (.A0(_1027_),
    .A1(_0773_),
    .S(_0899_),
    .X(_1028_));
 sky130_fd_sc_hd__xnor2_4 _4227_ (.A(_1026_),
    .B(_1028_),
    .Y(_1029_));
 sky130_fd_sc_hd__xor2_2 _4228_ (.A(_0986_),
    .B(_1029_),
    .X(\sbox1.ah[1] ));
 sky130_fd_sc_hd__mux2_1 _4229_ (.A0(net350),
    .A1(\mix1.data_o[66] ),
    .S(_0721_),
    .X(_1030_));
 sky130_fd_sc_hd__mux2_1 _4230_ (.A0(net368),
    .A1(\mix1.data_o[82] ),
    .S(_0738_),
    .X(_1031_));
 sky130_fd_sc_hd__a22o_1 _4231_ (.A1(_0709_),
    .A2(_1030_),
    .B1(_1031_),
    .B2(_0724_),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_1 _4232_ (.A0(net310),
    .A1(\mix1.data_o[2] ),
    .S(_0721_),
    .X(_1033_));
 sky130_fd_sc_hd__mux2_1 _4233_ (.A0(net377),
    .A1(\mix1.data_o[90] ),
    .S(_0738_),
    .X(_1034_));
 sky130_fd_sc_hd__a22o_1 _4234_ (.A1(_0712_),
    .A2(_1033_),
    .B1(_1034_),
    .B2(_0727_),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _4235_ (.A0(net359),
    .A1(\mix1.data_o[74] ),
    .S(_0860_),
    .X(_1036_));
 sky130_fd_sc_hd__mux2_1 _4236_ (.A0(net306),
    .A1(\mix1.data_o[26] ),
    .S(_0862_),
    .X(_1037_));
 sky130_fd_sc_hd__a22o_1 _4237_ (.A1(_0740_),
    .A2(_1036_),
    .B1(_1037_),
    .B2(_0713_),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_1 _4238_ (.A0(net276),
    .A1(\mix1.data_o[114] ),
    .S(_0721_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _4239_ (.A0(net271),
    .A1(\mix1.data_o[10] ),
    .S(_0738_),
    .X(_1040_));
 sky130_fd_sc_hd__a22o_1 _4240_ (.A1(_0706_),
    .A2(_1039_),
    .B1(_1040_),
    .B2(_0743_),
    .X(_1041_));
 sky130_fd_sc_hd__or4_1 _4241_ (.A(_1032_),
    .B(_1035_),
    .C(_1038_),
    .D(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_1 _4242_ (.A0(net285),
    .A1(\mix1.data_o[122] ),
    .S(_0862_),
    .X(_1043_));
 sky130_fd_sc_hd__a31o_1 _4243_ (.A1(_0719_),
    .A2(_0720_),
    .A3(_1043_),
    .B1(_0791_),
    .X(_1044_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(net385),
    .A1(\mix1.data_o[98] ),
    .S(_0833_),
    .X(_1045_));
 sky130_fd_sc_hd__a22o_1 _4245_ (.A1(net333),
    .A2(_0794_),
    .B1(_0703_),
    .B2(net324),
    .X(_1046_));
 sky130_fd_sc_hd__or2_1 _4246_ (.A(net341),
    .B(_0737_),
    .X(_1047_));
 sky130_fd_sc_hd__o211a_1 _4247_ (.A1(\mix1.data_o[58] ),
    .A2(_0879_),
    .B1(_0697_),
    .C1(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__a221o_1 _4248_ (.A1(_0687_),
    .A2(_1045_),
    .B1(_1046_),
    .B2(_0797_),
    .C1(_1048_),
    .X(_1049_));
 sky130_fd_sc_hd__mux2_1 _4249_ (.A0(net267),
    .A1(\mix1.data_o[106] ),
    .S(_0860_),
    .X(_1050_));
 sky130_fd_sc_hd__mux2_1 _4250_ (.A0(net315),
    .A1(\mix1.data_o[34] ),
    .S(_0862_),
    .X(_1051_));
 sky130_fd_sc_hd__a22o_1 _4251_ (.A1(_0692_),
    .A2(_1050_),
    .B1(_1051_),
    .B2(_0730_),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _4252_ (.A0(net297),
    .A1(\mix1.data_o[18] ),
    .S(_0721_),
    .X(_1053_));
 sky130_fd_sc_hd__a22o_1 _4253_ (.A1(\mix1.data_o[50] ),
    .A2(_0794_),
    .B1(_0795_),
    .B2(\mix1.data_o[42] ),
    .X(_1054_));
 sky130_fd_sc_hd__a22o_1 _4254_ (.A1(_0734_),
    .A2(_1053_),
    .B1(_1054_),
    .B2(_0807_),
    .X(_1055_));
 sky130_fd_sc_hd__or4_1 _4255_ (.A(_1044_),
    .B(_1049_),
    .C(_1052_),
    .D(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__clkbuf_8 _4256_ (.A(_0766_),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _4257_ (.A0(\ks1.key_reg[2] ),
    .A1(net180),
    .S(_0815_),
    .X(_1057_));
 sky130_fd_sc_hd__mux2_1 _4258_ (.A0(\ks1.key_reg[10] ),
    .A1(net141),
    .S(_0767_),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _4259_ (.A0(\ks1.key_reg[18] ),
    .A1(net167),
    .S(_0767_),
    .X(_1059_));
 sky130_fd_sc_hd__a22o_1 _4260_ (.A1(_0757_),
    .A2(_1058_),
    .B1(_1059_),
    .B2(_0763_),
    .X(_1060_));
 sky130_fd_sc_hd__mux2_1 _4261_ (.A0(\ks1.key_reg[26] ),
    .A1(net176),
    .S(_0761_),
    .X(_1061_));
 sky130_fd_sc_hd__a21o_1 _4262_ (.A1(_0769_),
    .A2(_1061_),
    .B1(_0755_),
    .X(_1062_));
 sky130_fd_sc_hd__a211o_1 _4263_ (.A1(_0649_),
    .A2(_1057_),
    .B1(_1060_),
    .C1(_1062_),
    .X(_1063_));
 sky130_fd_sc_hd__o21a_2 _4264_ (.A1(_1042_),
    .A2(_1056_),
    .B1(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__xnor2_2 _4265_ (.A(_1024_),
    .B(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__xnor2_1 _4266_ (.A(_0898_),
    .B(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__mux2_4 _4267_ (.A0(_1066_),
    .A1(_0982_),
    .S(_0899_),
    .X(_1067_));
 sky130_fd_sc_hd__xor2_4 _4268_ (.A(_1026_),
    .B(_1067_),
    .X(\sbox1.ah[3] ));
 sky130_fd_sc_hd__xor2_2 _4269_ (.A(_0986_),
    .B(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__inv_2 _4270_ (.A(_1068_),
    .Y(\sbox1.ah[0] ));
 sky130_fd_sc_hd__inv_2 _4271_ (.A(_1064_),
    .Y(_1069_));
 sky130_fd_sc_hd__xnor2_1 _4272_ (.A(_0983_),
    .B(_1069_),
    .Y(_1070_));
 sky130_fd_sc_hd__mux2_1 _4273_ (.A0(_1070_),
    .A1(_0857_),
    .S(_0899_),
    .X(_1071_));
 sky130_fd_sc_hd__xor2_1 _4274_ (.A(\sbox1.ah[3] ),
    .B(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__xnor2_1 _4275_ (.A(_0987_),
    .B(_1024_),
    .Y(_1073_));
 sky130_fd_sc_hd__buf_4 _4276_ (.A(_0899_),
    .X(_1074_));
 sky130_fd_sc_hd__mux2_4 _4277_ (.A0(_1073_),
    .A1(_1069_),
    .S(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__xor2_2 _4278_ (.A(_1072_),
    .B(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__inv_2 _4279_ (.A(_1076_),
    .Y(\sbox1.ah[2] ));
 sky130_fd_sc_hd__xnor2_4 _4280_ (.A(_0900_),
    .B(_1075_),
    .Y(_1077_));
 sky130_fd_sc_hd__xnor2_1 _4281_ (.A(\sbox1.ah[3] ),
    .B(_1077_),
    .Y(\sbox1.next_alph[3] ));
 sky130_fd_sc_hd__inv_2 _4282_ (.A(_1029_),
    .Y(_1078_));
 sky130_fd_sc_hd__nand2_1 _4283_ (.A(_1078_),
    .B(\sbox1.ah[2] ),
    .Y(_1079_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_1029_),
    .B(_1076_),
    .Y(_1080_));
 sky130_fd_sc_hd__nand2_1 _4285_ (.A(_1079_),
    .B(_1080_),
    .Y(\sbox1.next_alph[2] ));
 sky130_fd_sc_hd__xnor2_4 _4286_ (.A(_1028_),
    .B(_1075_),
    .Y(_1081_));
 sky130_fd_sc_hd__xor2_1 _4287_ (.A(\sbox1.ah[1] ),
    .B(_1081_),
    .X(\sbox1.next_alph[1] ));
 sky130_fd_sc_hd__xor2_1 _4288_ (.A(_0982_),
    .B(_1065_),
    .X(_1082_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(_1082_),
    .A1(_0940_),
    .S(_1074_),
    .X(_1083_));
 sky130_fd_sc_hd__inv_2 _4290_ (.A(_1083_),
    .Y(\sbox1.next_alph[0] ));
 sky130_fd_sc_hd__xnor2_1 _4291_ (.A(_1068_),
    .B(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(_1077_),
    .A1(_1084_),
    .S(\sbox1.ah[3] ),
    .X(_1085_));
 sky130_fd_sc_hd__and2_1 _4293_ (.A(\sbox1.ah[0] ),
    .B(_1077_),
    .X(_1086_));
 sky130_fd_sc_hd__nand2_1 _4294_ (.A(_0986_),
    .B(_1078_),
    .Y(_1087_));
 sky130_fd_sc_hd__nand2_1 _4295_ (.A(\sbox1.ah[2] ),
    .B(_1081_),
    .Y(_1088_));
 sky130_fd_sc_hd__xnor2_1 _4296_ (.A(_1087_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__xnor2_1 _4297_ (.A(_1086_),
    .B(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__xnor2_1 _4298_ (.A(_1085_),
    .B(_1090_),
    .Y(\sbox1.intermediate_to_invert_var[3] ));
 sky130_fd_sc_hd__xnor2_1 _4299_ (.A(_1029_),
    .B(_1077_),
    .Y(_1091_));
 sky130_fd_sc_hd__xnor2_1 _4300_ (.A(_1077_),
    .B(_1084_),
    .Y(_1092_));
 sky130_fd_sc_hd__a211o_1 _4301_ (.A1(\sbox1.ah[3] ),
    .A2(_1091_),
    .B1(_1092_),
    .C1(_1076_),
    .X(_1093_));
 sky130_fd_sc_hd__o211ai_1 _4302_ (.A1(_1076_),
    .A2(_1092_),
    .B1(_1091_),
    .C1(\sbox1.ah[3] ),
    .Y(_1094_));
 sky130_fd_sc_hd__nand2_1 _4303_ (.A(_1093_),
    .B(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__nor2_1 _4304_ (.A(_0986_),
    .B(_1067_),
    .Y(_1096_));
 sky130_fd_sc_hd__o2bb2a_1 _4305_ (.A1_N(\sbox1.ah[1] ),
    .A2_N(_1081_),
    .B1(_1068_),
    .B2(_1078_),
    .X(_1097_));
 sky130_fd_sc_hd__a31o_1 _4306_ (.A1(_1029_),
    .A2(_1096_),
    .A3(_1081_),
    .B1(_1097_),
    .X(_1098_));
 sky130_fd_sc_hd__xnor2_1 _4307_ (.A(_0900_),
    .B(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__xnor2_1 _4308_ (.A(_1095_),
    .B(_1099_),
    .Y(\sbox1.intermediate_to_invert_var[2] ));
 sky130_fd_sc_hd__nand2_1 _4309_ (.A(\sbox1.ah[2] ),
    .B(_1091_),
    .Y(_1100_));
 sky130_fd_sc_hd__nand2_1 _4310_ (.A(\sbox1.ah[3] ),
    .B(_1081_),
    .Y(_1101_));
 sky130_fd_sc_hd__o21ai_1 _4311_ (.A1(_1078_),
    .A2(\sbox1.ah[3] ),
    .B1(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__xnor2_1 _4312_ (.A(_1100_),
    .B(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__nor2_1 _4313_ (.A(_1068_),
    .B(_1081_),
    .Y(_1104_));
 sky130_fd_sc_hd__inv_2 _4314_ (.A(\sbox1.ah[1] ),
    .Y(_1105_));
 sky130_fd_sc_hd__nor2_1 _4315_ (.A(_1105_),
    .B(_1092_),
    .Y(_1106_));
 sky130_fd_sc_hd__xnor2_1 _4316_ (.A(_1104_),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__xnor2_1 _4317_ (.A(_1103_),
    .B(_1107_),
    .Y(\sbox1.intermediate_to_invert_var[1] ));
 sky130_fd_sc_hd__or2_1 _4318_ (.A(_1105_),
    .B(_1077_),
    .X(_1108_));
 sky130_fd_sc_hd__xnor2_1 _4319_ (.A(_1101_),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__xnor2_1 _4320_ (.A(_1079_),
    .B(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(_0986_),
    .A1(_1067_),
    .S(\sbox1.next_alph[0] ),
    .X(_1111_));
 sky130_fd_sc_hd__xnor2_1 _4322_ (.A(_1110_),
    .B(_1111_),
    .Y(\sbox1.intermediate_to_invert_var[0] ));
 sky130_fd_sc_hd__inv_2 _4323_ (.A(_0754_),
    .Y(_1112_));
 sky130_fd_sc_hd__buf_4 _4324_ (.A(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__buf_4 _4325_ (.A(_1113_),
    .X(\ks1.next_ready_o ));
 sky130_fd_sc_hd__clkinv_4 _4326_ (.A(state),
    .Y(_1114_));
 sky130_fd_sc_hd__buf_4 _4327_ (.A(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__and2_1 _4328_ (.A(_1115_),
    .B(net258),
    .X(_1116_));
 sky130_fd_sc_hd__clkbuf_1 _4329_ (.A(_1116_),
    .X(next_first_round_reg));
 sky130_fd_sc_hd__a21oi_2 _4330_ (.A1(addroundkey_ready_o),
    .A2(_0683_),
    .B1(_1115_),
    .Y(_1117_));
 sky130_fd_sc_hd__or2_1 _4331_ (.A(next_first_round_reg),
    .B(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__clkbuf_1 _4332_ (.A(_1118_),
    .X(next_state));
 sky130_fd_sc_hd__buf_6 _4333_ (.A(\sub1.ready_o ),
    .X(_1119_));
 sky130_fd_sc_hd__buf_4 _4334_ (.A(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__buf_6 _4335_ (.A(net129),
    .X(_1121_));
 sky130_fd_sc_hd__nand2_8 _4336_ (.A(_1121_),
    .B(_1119_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand2_4 _4337_ (.A(_0682_),
    .B(\mix1.ready_o ),
    .Y(_1123_));
 sky130_fd_sc_hd__nand2_2 _4338_ (.A(_1122_),
    .B(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__or2_1 _4339_ (.A(first_round_reg),
    .B(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__and4bb_1 _4340_ (.A_N(_0665_),
    .B_N(\round[2] ),
    .C(\round[3] ),
    .D(_0667_),
    .X(_1126_));
 sky130_fd_sc_hd__mux2_4 _4341_ (.A0(_0672_),
    .A1(_1126_),
    .S(_0682_),
    .X(_1127_));
 sky130_fd_sc_hd__inv_2 _4342_ (.A(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(_1120_),
    .A1(_1125_),
    .S(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__a22o_1 _4344_ (.A1(_1115_),
    .A2(net483),
    .B1(_1117_),
    .B2(_1129_),
    .X(next_addroundkey_start_i));
 sky130_fd_sc_hd__nor2_1 _4345_ (.A(\addroundkey_round[0] ),
    .B(_0750_),
    .Y(_1130_));
 sky130_fd_sc_hd__a211o_1 _4346_ (.A1(\addroundkey_round[0] ),
    .A2(_0670_),
    .B1(_0759_),
    .C1(_1130_),
    .X(_0000_));
 sky130_fd_sc_hd__inv_2 _4347_ (.A(_0750_),
    .Y(_1131_));
 sky130_fd_sc_hd__xor2_2 _4348_ (.A(\addroundkey_round[0] ),
    .B(\addroundkey_round[1] ),
    .X(_1132_));
 sky130_fd_sc_hd__a32o_1 _4349_ (.A1(\addroundkey_round[1] ),
    .A2(_0670_),
    .A3(_0748_),
    .B1(_1131_),
    .B2(_1132_),
    .X(_0001_));
 sky130_fd_sc_hd__and3_1 _4350_ (.A(\addroundkey_round[0] ),
    .B(\addroundkey_round[1] ),
    .C(\addroundkey_round[2] ),
    .X(_1133_));
 sky130_fd_sc_hd__a21oi_1 _4351_ (.A1(\addroundkey_round[0] ),
    .A2(\addroundkey_round[1] ),
    .B1(\addroundkey_round[2] ),
    .Y(_1134_));
 sky130_fd_sc_hd__nor3_2 _4352_ (.A(_0750_),
    .B(_1133_),
    .C(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hd__a31o_1 _4353_ (.A1(\addroundkey_round[2] ),
    .A2(_0670_),
    .A3(_0748_),
    .B1(_1135_),
    .X(_0002_));
 sky130_fd_sc_hd__xnor2_1 _4354_ (.A(\addroundkey_round[3] ),
    .B(_1133_),
    .Y(_1136_));
 sky130_fd_sc_hd__nor2_1 _4355_ (.A(_0750_),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__a31o_1 _4356_ (.A1(\addroundkey_round[3] ),
    .A2(_0670_),
    .A3(_0748_),
    .B1(_1137_),
    .X(_0003_));
 sky130_fd_sc_hd__clkbuf_4 _4357_ (.A(_0660_),
    .X(_1138_));
 sky130_fd_sc_hd__clkbuf_4 _4358_ (.A(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__clkbuf_4 _4359_ (.A(_1139_),
    .X(_1140_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B(\sbox1.inversion_to_invert_var[0] ),
    .Y(_1141_));
 sky130_fd_sc_hd__or3_1 _4361_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B(\sbox1.inversion_to_invert_var[2] ),
    .C(\sbox1.inversion_to_invert_var[0] ),
    .X(_1142_));
 sky130_fd_sc_hd__a21boi_4 _4362_ (.A1(\sbox1.inversion_to_invert_var[1] ),
    .A2(\sbox1.inversion_to_invert_var[2] ),
    .B1_N(\sbox1.inversion_to_invert_var[3] ),
    .Y(_1143_));
 sky130_fd_sc_hd__a21oi_1 _4363_ (.A1(_1141_),
    .A2(_1142_),
    .B1(_1143_),
    .Y(_1144_));
 sky130_fd_sc_hd__and3_1 _4364_ (.A(_1143_),
    .B(_1141_),
    .C(_1142_),
    .X(_1145_));
 sky130_fd_sc_hd__nor2_2 _4365_ (.A(_1144_),
    .B(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__nand2_1 _4366_ (.A(\sbox1.alph[0] ),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__and2_1 _4367_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B(\sbox1.inversion_to_invert_var[0] ),
    .X(_1148_));
 sky130_fd_sc_hd__a21oi_1 _4368_ (.A1(\sbox1.inversion_to_invert_var[2] ),
    .A2(\sbox1.inversion_to_invert_var[0] ),
    .B1(\sbox1.inversion_to_invert_var[3] ),
    .Y(_1149_));
 sky130_fd_sc_hd__and3_1 _4369_ (.A(\sbox1.inversion_to_invert_var[2] ),
    .B(\sbox1.inversion_to_invert_var[3] ),
    .C(\sbox1.inversion_to_invert_var[0] ),
    .X(_1150_));
 sky130_fd_sc_hd__nand2_1 _4370_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B(\sbox1.inversion_to_invert_var[2] ),
    .Y(_1151_));
 sky130_fd_sc_hd__o311a_1 _4371_ (.A1(\sbox1.inversion_to_invert_var[1] ),
    .A2(_1149_),
    .A3(_1150_),
    .B1(_1151_),
    .C1(_1141_),
    .X(_1152_));
 sky130_fd_sc_hd__a21oi_4 _4372_ (.A1(\sbox1.inversion_to_invert_var[3] ),
    .A2(_1148_),
    .B1(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2_1 _4373_ (.A(\sbox1.alph[3] ),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__xnor2_2 _4374_ (.A(_1147_),
    .B(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hd__xnor2_2 _4375_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B(\sbox1.inversion_to_invert_var[2] ),
    .Y(_1156_));
 sky130_fd_sc_hd__inv_2 _4376_ (.A(\sbox1.inversion_to_invert_var[3] ),
    .Y(_1157_));
 sky130_fd_sc_hd__and3b_1 _4377_ (.A_N(\sbox1.inversion_to_invert_var[0] ),
    .B(\sbox1.inversion_to_invert_var[2] ),
    .C(\sbox1.inversion_to_invert_var[1] ),
    .X(_1158_));
 sky130_fd_sc_hd__a221oi_4 _4378_ (.A1(\sbox1.inversion_to_invert_var[0] ),
    .A2(_1143_),
    .B1(_1156_),
    .B2(_1157_),
    .C1(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__nand2_1 _4379_ (.A(\sbox1.alph[1] ),
    .B(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__and2_1 _4380_ (.A(_1148_),
    .B(_1150_),
    .X(_1161_));
 sky130_fd_sc_hd__nand2_1 _4381_ (.A(\sbox1.inversion_to_invert_var[2] ),
    .B(\sbox1.inversion_to_invert_var[3] ),
    .Y(_1162_));
 sky130_fd_sc_hd__o21ba_1 _4382_ (.A1(\sbox1.inversion_to_invert_var[2] ),
    .A2(\sbox1.inversion_to_invert_var[3] ),
    .B1_N(\sbox1.inversion_to_invert_var[0] ),
    .X(_1163_));
 sky130_fd_sc_hd__a211oi_2 _4383_ (.A1(_1162_),
    .A2(_1163_),
    .B1(_1148_),
    .C1(_1150_),
    .Y(_1164_));
 sky130_fd_sc_hd__nor2_2 _4384_ (.A(_1161_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__nand2_1 _4385_ (.A(\sbox1.alph[2] ),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__xnor2_2 _4386_ (.A(_1160_),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__xnor2_4 _4387_ (.A(_1155_),
    .B(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__nand2_1 _4388_ (.A(\sbox1.ah_reg[0] ),
    .B(_1146_),
    .Y(_1169_));
 sky130_fd_sc_hd__nand2_1 _4389_ (.A(\sbox1.ah_reg[1] ),
    .B(_1159_),
    .Y(_1170_));
 sky130_fd_sc_hd__xnor2_2 _4390_ (.A(_1169_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__nand2_1 _4391_ (.A(\sbox1.ah_reg[3] ),
    .B(_1153_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_1 _4392_ (.A(\sbox1.ah_reg[2] ),
    .B(_1165_),
    .Y(_1173_));
 sky130_fd_sc_hd__xnor2_2 _4393_ (.A(_1172_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__xnor2_4 _4394_ (.A(_1171_),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__xor2_4 _4395_ (.A(_1168_),
    .B(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__o21ai_1 _4396_ (.A1(_1161_),
    .A2(_1164_),
    .B1(_1159_),
    .Y(_1177_));
 sky130_fd_sc_hd__or3_1 _4397_ (.A(_1159_),
    .B(_1161_),
    .C(_1164_),
    .X(_1178_));
 sky130_fd_sc_hd__inv_2 _4398_ (.A(\sbox1.alph[3] ),
    .Y(_1179_));
 sky130_fd_sc_hd__a21oi_1 _4399_ (.A1(_1177_),
    .A2(_1178_),
    .B1(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__a221o_1 _4400_ (.A1(\sbox1.inversion_to_invert_var[0] ),
    .A2(_1143_),
    .B1(_1156_),
    .B2(_1157_),
    .C1(_1158_),
    .X(_1181_));
 sky130_fd_sc_hd__or3_1 _4401_ (.A(_1144_),
    .B(_1145_),
    .C(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__o21ai_1 _4402_ (.A1(_1144_),
    .A2(_1145_),
    .B1(_1181_),
    .Y(_1183_));
 sky130_fd_sc_hd__and3_1 _4403_ (.A(\sbox1.alph[2] ),
    .B(_1182_),
    .C(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__xnor2_2 _4404_ (.A(_1180_),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__nand2_1 _4405_ (.A(\sbox1.alph[0] ),
    .B(_1165_),
    .Y(_1186_));
 sky130_fd_sc_hd__nand2_1 _4406_ (.A(\sbox1.alph[1] ),
    .B(_1153_),
    .Y(_1187_));
 sky130_fd_sc_hd__xnor2_2 _4407_ (.A(_1186_),
    .B(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__xnor2_4 _4408_ (.A(_1185_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__nand2_1 _4409_ (.A(\sbox1.ah_reg[1] ),
    .B(_1146_),
    .Y(_1190_));
 sky130_fd_sc_hd__xor2_1 _4410_ (.A(\sbox1.ah_reg[0] ),
    .B(\sbox1.ah_reg[3] ),
    .X(_1191_));
 sky130_fd_sc_hd__nand2_1 _4411_ (.A(_1153_),
    .B(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__xnor2_1 _4412_ (.A(_1190_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__xor2_1 _4413_ (.A(\sbox1.ah_reg[2] ),
    .B(\sbox1.ah_reg[1] ),
    .X(_1194_));
 sky130_fd_sc_hd__nand2_1 _4414_ (.A(_1159_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__xor2_1 _4415_ (.A(\sbox1.ah_reg[3] ),
    .B(\sbox1.ah_reg[2] ),
    .X(_1196_));
 sky130_fd_sc_hd__nand2_1 _4416_ (.A(_1165_),
    .B(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__xnor2_1 _4417_ (.A(_1195_),
    .B(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hd__xnor2_2 _4418_ (.A(_1193_),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__xnor2_4 _4419_ (.A(_1175_),
    .B(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nand2_1 _4420_ (.A(\sbox1.ah_reg[3] ),
    .B(_1146_),
    .Y(_1201_));
 sky130_fd_sc_hd__nand2_1 _4421_ (.A(_1159_),
    .B(_1191_),
    .Y(_1202_));
 sky130_fd_sc_hd__xnor2_2 _4422_ (.A(_1201_),
    .B(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__nand2_1 _4423_ (.A(\sbox1.ah_reg[2] ),
    .B(_1153_),
    .Y(_1204_));
 sky130_fd_sc_hd__nand2_1 _4424_ (.A(\sbox1.ah_reg[1] ),
    .B(_1165_),
    .Y(_1205_));
 sky130_fd_sc_hd__xnor2_2 _4425_ (.A(_1204_),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__xnor2_4 _4426_ (.A(_1203_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__xor2_4 _4427_ (.A(_1200_),
    .B(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__xnor2_4 _4428_ (.A(_1189_),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__xor2_1 _4429_ (.A(_1168_),
    .B(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__mux2_1 _4430_ (.A0(_1176_),
    .A1(_1210_),
    .S(_0899_),
    .X(_1211_));
 sky130_fd_sc_hd__buf_6 _4431_ (.A(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__buf_4 _4432_ (.A(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__clkbuf_8 _4433_ (.A(_0682_),
    .X(_1214_));
 sky130_fd_sc_hd__nor2_2 _4434_ (.A(_1214_),
    .B(_1138_),
    .Y(_1215_));
 sky130_fd_sc_hd__clkbuf_4 _4435_ (.A(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__buf_4 _4436_ (.A(_1121_),
    .X(_1217_));
 sky130_fd_sc_hd__buf_4 _4437_ (.A(_1217_),
    .X(_1218_));
 sky130_fd_sc_hd__buf_6 _4438_ (.A(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__nor2_2 _4439_ (.A(_1219_),
    .B(_1139_),
    .Y(_1220_));
 sky130_fd_sc_hd__or2_4 _4440_ (.A(_0685_),
    .B(_0691_),
    .X(_1221_));
 sky130_fd_sc_hd__and3_1 _4441_ (.A(\sub1.data_o[112] ),
    .B(_1138_),
    .C(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__a221o_1 _4442_ (.A1(\sub1.data_o[16] ),
    .A2(_1216_),
    .B1(_1220_),
    .B2(\sub1.data_o[80] ),
    .C1(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__a31o_1 _4443_ (.A1(_1140_),
    .A2(_0923_),
    .A3(_1213_),
    .B1(_1223_),
    .X(_0004_));
 sky130_fd_sc_hd__xnor2_2 _4444_ (.A(_1189_),
    .B(_1207_),
    .Y(_1224_));
 sky130_fd_sc_hd__nand2_1 _4445_ (.A(\sbox1.alph[0] ),
    .B(_1159_),
    .Y(_1225_));
 sky130_fd_sc_hd__and3_1 _4446_ (.A(\sbox1.alph[3] ),
    .B(_1182_),
    .C(_1183_),
    .X(_1226_));
 sky130_fd_sc_hd__xnor2_2 _4447_ (.A(_1225_),
    .B(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__nand2_1 _4448_ (.A(\sbox1.alph[1] ),
    .B(_1165_),
    .Y(_1228_));
 sky130_fd_sc_hd__nand2_1 _4449_ (.A(\sbox1.alph[2] ),
    .B(_1153_),
    .Y(_1229_));
 sky130_fd_sc_hd__xnor2_2 _4450_ (.A(_1228_),
    .B(_1229_),
    .Y(_1230_));
 sky130_fd_sc_hd__xnor2_4 _4451_ (.A(_1227_),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__o21ai_1 _4452_ (.A1(_1179_),
    .A2(_1165_),
    .B1(_1153_),
    .Y(_1232_));
 sky130_fd_sc_hd__inv_2 _4453_ (.A(\sbox1.alph[0] ),
    .Y(_1233_));
 sky130_fd_sc_hd__a211o_1 _4454_ (.A1(_1233_),
    .A2(_1153_),
    .B1(_1165_),
    .C1(_1179_),
    .X(_1234_));
 sky130_fd_sc_hd__o221a_2 _4455_ (.A1(\sbox1.alph[3] ),
    .A2(_1153_),
    .B1(_1232_),
    .B2(\sbox1.alph[0] ),
    .C1(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__a21bo_1 _4456_ (.A1(_1177_),
    .A2(_1178_),
    .B1_N(\sbox1.alph[2] ),
    .X(_1236_));
 sky130_fd_sc_hd__and3_1 _4457_ (.A(\sbox1.alph[1] ),
    .B(_1182_),
    .C(_1183_),
    .X(_1237_));
 sky130_fd_sc_hd__xnor2_2 _4458_ (.A(_1236_),
    .B(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hd__xnor2_4 _4459_ (.A(_1235_),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__xnor2_4 _4460_ (.A(_1231_),
    .B(_1239_),
    .Y(_1240_));
 sky130_fd_sc_hd__xnor2_4 _4461_ (.A(_1224_),
    .B(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__xnor2_4 _4462_ (.A(_1175_),
    .B(_1241_),
    .Y(_1242_));
 sky130_fd_sc_hd__xnor2_1 _4463_ (.A(_1200_),
    .B(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__xnor2_1 _4464_ (.A(_1176_),
    .B(_1243_),
    .Y(_1244_));
 sky130_fd_sc_hd__mux2_1 _4465_ (.A0(_1208_),
    .A1(_1244_),
    .S(_0899_),
    .X(_1245_));
 sky130_fd_sc_hd__buf_6 _4466_ (.A(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__buf_4 _4467_ (.A(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__and3_1 _4468_ (.A(\sub1.data_o[113] ),
    .B(_1138_),
    .C(_1221_),
    .X(_1248_));
 sky130_fd_sc_hd__a221o_1 _4469_ (.A1(\sub1.data_o[17] ),
    .A2(_1216_),
    .B1(_1220_),
    .B2(\sub1.data_o[81] ),
    .C1(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__a31o_1 _4470_ (.A1(_1140_),
    .A2(_0923_),
    .A3(_1247_),
    .B1(_1249_),
    .X(_0005_));
 sky130_fd_sc_hd__xnor2_4 _4471_ (.A(_1209_),
    .B(_1242_),
    .Y(_1250_));
 sky130_fd_sc_hd__xnor2_1 _4472_ (.A(_1176_),
    .B(_1239_),
    .Y(_1251_));
 sky130_fd_sc_hd__nor2_1 _4473_ (.A(_1250_),
    .B(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__a21bo_1 _4474_ (.A1(_1250_),
    .A2(_1251_),
    .B1_N(_1074_),
    .X(_1253_));
 sky130_fd_sc_hd__xnor2_2 _4475_ (.A(_1200_),
    .B(_1239_),
    .Y(_1254_));
 sky130_fd_sc_hd__xor2_2 _4476_ (.A(_1207_),
    .B(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__o22a_4 _4477_ (.A1(_1252_),
    .A2(_1253_),
    .B1(_1255_),
    .B2(_1074_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_4 _4478_ (.A(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__and3_1 _4479_ (.A(\sub1.data_o[114] ),
    .B(_1138_),
    .C(_1221_),
    .X(_1258_));
 sky130_fd_sc_hd__a221o_1 _4480_ (.A1(\sub1.data_o[18] ),
    .A2(_1216_),
    .B1(_1220_),
    .B2(\sub1.data_o[82] ),
    .C1(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__a31o_1 _4481_ (.A1(_1140_),
    .A2(_0923_),
    .A3(_1257_),
    .B1(_1259_),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _4482_ (.A(\sbox1.ah_reg[2] ),
    .B(_1146_),
    .Y(_1260_));
 sky130_fd_sc_hd__nand2_1 _4483_ (.A(_1159_),
    .B(_1196_),
    .Y(_1261_));
 sky130_fd_sc_hd__xnor2_2 _4484_ (.A(_1260_),
    .B(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__nand2_1 _4485_ (.A(\sbox1.ah_reg[1] ),
    .B(_1153_),
    .Y(_1263_));
 sky130_fd_sc_hd__nand2_1 _4486_ (.A(_1165_),
    .B(_1191_),
    .Y(_1264_));
 sky130_fd_sc_hd__xnor2_2 _4487_ (.A(_1263_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__xnor2_4 _4488_ (.A(_1262_),
    .B(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__xor2_1 _4489_ (.A(_1254_),
    .B(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__xor2_4 _4490_ (.A(_1207_),
    .B(_1266_),
    .X(_1268_));
 sky130_fd_sc_hd__xnor2_4 _4491_ (.A(_1176_),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__xor2_4 _4492_ (.A(_1189_),
    .B(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_8 _4493_ (.A0(_1267_),
    .A1(_1270_),
    .S(_1074_),
    .X(_1271_));
 sky130_fd_sc_hd__buf_6 _4494_ (.A(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__and3_1 _4495_ (.A(\sub1.data_o[115] ),
    .B(_1138_),
    .C(_1221_),
    .X(_1273_));
 sky130_fd_sc_hd__a221o_1 _4496_ (.A1(\sub1.data_o[19] ),
    .A2(_1216_),
    .B1(_1220_),
    .B2(\sub1.data_o[83] ),
    .C1(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__a31o_1 _4497_ (.A1(_1140_),
    .A2(_0923_),
    .A3(_1272_),
    .B1(_1274_),
    .X(_0007_));
 sky130_fd_sc_hd__xor2_1 _4498_ (.A(_1231_),
    .B(_1255_),
    .X(_1275_));
 sky130_fd_sc_hd__xnor2_1 _4499_ (.A(_1240_),
    .B(_1269_),
    .Y(_1276_));
 sky130_fd_sc_hd__mux2_8 _4500_ (.A0(_1275_),
    .A1(_1276_),
    .S(_1074_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_8 _4501_ (.A(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__and3_1 _4502_ (.A(\sub1.data_o[116] ),
    .B(_1138_),
    .C(_1221_),
    .X(_1279_));
 sky130_fd_sc_hd__a221o_1 _4503_ (.A1(\sub1.data_o[20] ),
    .A2(_1216_),
    .B1(_1220_),
    .B2(\sub1.data_o[84] ),
    .C1(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__a31o_1 _4504_ (.A1(_1140_),
    .A2(_0923_),
    .A3(_1278_),
    .B1(_1280_),
    .X(_0008_));
 sky130_fd_sc_hd__xor2_1 _4505_ (.A(_1200_),
    .B(_1266_),
    .X(_1281_));
 sky130_fd_sc_hd__xnor2_2 _4506_ (.A(_1241_),
    .B(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__o21ba_1 _4507_ (.A1(_1189_),
    .A2(_1200_),
    .B1_N(_1074_),
    .X(_1283_));
 sky130_fd_sc_hd__nand2_1 _4508_ (.A(_1189_),
    .B(_1200_),
    .Y(_1284_));
 sky130_fd_sc_hd__a22o_4 _4509_ (.A1(_1074_),
    .A2(_1282_),
    .B1(_1283_),
    .B2(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__buf_6 _4510_ (.A(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__and3_1 _4511_ (.A(\sub1.data_o[117] ),
    .B(_1138_),
    .C(_1221_),
    .X(_1287_));
 sky130_fd_sc_hd__a221o_1 _4512_ (.A1(\sub1.data_o[21] ),
    .A2(_1216_),
    .B1(_1220_),
    .B2(\sub1.data_o[85] ),
    .C1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__a31o_1 _4513_ (.A1(_1140_),
    .A2(_0923_),
    .A3(_1286_),
    .B1(_1288_),
    .X(_0009_));
 sky130_fd_sc_hd__nand2_1 _4514_ (.A(_1175_),
    .B(_1268_),
    .Y(_1289_));
 sky130_fd_sc_hd__or2_1 _4515_ (.A(_1175_),
    .B(_1268_),
    .X(_1290_));
 sky130_fd_sc_hd__and3_1 _4516_ (.A(net129),
    .B(_0755_),
    .C(_1242_),
    .X(_1291_));
 sky130_fd_sc_hd__a31o_4 _4517_ (.A1(_1074_),
    .A2(_1289_),
    .A3(_1290_),
    .B1(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_4 _4518_ (.A(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__and3_1 _4519_ (.A(\sub1.data_o[118] ),
    .B(_1138_),
    .C(_1221_),
    .X(_1294_));
 sky130_fd_sc_hd__a221o_1 _4520_ (.A1(\sub1.data_o[22] ),
    .A2(_1216_),
    .B1(_1220_),
    .B2(\sub1.data_o[86] ),
    .C1(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__a31o_1 _4521_ (.A1(_1140_),
    .A2(_0923_),
    .A3(_1293_),
    .B1(_1295_),
    .X(_0010_));
 sky130_fd_sc_hd__or2_1 _4522_ (.A(_1239_),
    .B(_1282_),
    .X(_1296_));
 sky130_fd_sc_hd__nand2_1 _4523_ (.A(_1239_),
    .B(_1282_),
    .Y(_1297_));
 sky130_fd_sc_hd__a31o_1 _4524_ (.A1(_1074_),
    .A2(_1296_),
    .A3(_1297_),
    .B1(_1291_),
    .X(_1298_));
 sky130_fd_sc_hd__xnor2_4 _4525_ (.A(_1250_),
    .B(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__clkbuf_4 _4526_ (.A(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__and3_1 _4527_ (.A(\sub1.data_o[119] ),
    .B(_1138_),
    .C(_1221_),
    .X(_1301_));
 sky130_fd_sc_hd__a221o_1 _4528_ (.A1(\sub1.data_o[23] ),
    .A2(_1216_),
    .B1(_1220_),
    .B2(\sub1.data_o[87] ),
    .C1(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__a31o_1 _4529_ (.A1(_1140_),
    .A2(_0923_),
    .A3(_1300_),
    .B1(_1302_),
    .X(_0011_));
 sky130_fd_sc_hd__nor2_1 _4530_ (.A(_0679_),
    .B(net258),
    .Y(_1303_));
 sky130_fd_sc_hd__and2_1 _4531_ (.A(_0682_),
    .B(\mix1.ready_o ),
    .X(_1304_));
 sky130_fd_sc_hd__buf_2 _4532_ (.A(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__clkbuf_4 _4533_ (.A(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_4 _4534_ (.A(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__or2_1 _4535_ (.A(_0667_),
    .B(_0665_),
    .X(_1308_));
 sky130_fd_sc_hd__nand2_1 _4536_ (.A(_0667_),
    .B(_0665_),
    .Y(_1309_));
 sky130_fd_sc_hd__nand2_1 _4537_ (.A(_1308_),
    .B(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__o2bb2a_1 _4538_ (.A1_N(_1307_),
    .A2_N(_1310_),
    .B1(_1124_),
    .B2(_0665_),
    .X(_1311_));
 sky130_fd_sc_hd__nand2_1 _4539_ (.A(_1120_),
    .B(_1310_),
    .Y(_1312_));
 sky130_fd_sc_hd__o211a_1 _4540_ (.A1(_1120_),
    .A2(_1311_),
    .B1(_1312_),
    .C1(_1127_),
    .X(_1313_));
 sky130_fd_sc_hd__nand2_1 _4541_ (.A(_0667_),
    .B(_1124_),
    .Y(_1314_));
 sky130_fd_sc_hd__or2_1 _4542_ (.A(_0667_),
    .B(_1124_),
    .X(_1315_));
 sky130_fd_sc_hd__and4b_1 _4543_ (.A_N(_1313_),
    .B(_1314_),
    .C(_1315_),
    .D(_1117_),
    .X(_1316_));
 sky130_fd_sc_hd__a21o_1 _4544_ (.A1(_0667_),
    .A2(_1303_),
    .B1(_1316_),
    .X(_0012_));
 sky130_fd_sc_hd__a21oi_1 _4545_ (.A1(_1214_),
    .A2(net258),
    .B1(_0679_),
    .Y(_1317_));
 sky130_fd_sc_hd__buf_4 _4546_ (.A(_1122_),
    .X(_1318_));
 sky130_fd_sc_hd__o211a_1 _4547_ (.A1(_1318_),
    .A2(_1310_),
    .B1(_1311_),
    .C1(_1128_),
    .X(_1319_));
 sky130_fd_sc_hd__o21a_1 _4548_ (.A1(_1313_),
    .A2(_1319_),
    .B1(_1117_),
    .X(_1320_));
 sky130_fd_sc_hd__o32a_1 _4549_ (.A1(_0679_),
    .A2(_0665_),
    .A3(net258),
    .B1(_1317_),
    .B2(_1320_),
    .X(_0013_));
 sky130_fd_sc_hd__nor2_1 _4550_ (.A(_0671_),
    .B(_1318_),
    .Y(_1321_));
 sky130_fd_sc_hd__o21a_1 _4551_ (.A1(_1308_),
    .A2(_1318_),
    .B1(\round[2] ),
    .X(_1322_));
 sky130_fd_sc_hd__or3_1 _4552_ (.A(_1307_),
    .B(_1321_),
    .C(_1322_),
    .X(_1323_));
 sky130_fd_sc_hd__a21oi_1 _4553_ (.A1(_0667_),
    .A2(_0665_),
    .B1(\round[2] ),
    .Y(_1324_));
 sky130_fd_sc_hd__and3_1 _4554_ (.A(_0667_),
    .B(_0665_),
    .C(\round[2] ),
    .X(_1325_));
 sky130_fd_sc_hd__o21a_1 _4555_ (.A1(_1324_),
    .A2(_1325_),
    .B1(_1307_),
    .X(_1326_));
 sky130_fd_sc_hd__nor2_1 _4556_ (.A(_1127_),
    .B(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__a32o_1 _4557_ (.A1(_0679_),
    .A2(_1323_),
    .A3(_1327_),
    .B1(\round[2] ),
    .B2(_1303_),
    .X(_0014_));
 sky130_fd_sc_hd__o21ai_1 _4558_ (.A1(_1219_),
    .A2(addroundkey_ready_o),
    .B1(_0683_),
    .Y(_1328_));
 sky130_fd_sc_hd__buf_4 _4559_ (.A(_1123_),
    .X(_1329_));
 sky130_fd_sc_hd__or2b_1 _4560_ (.A(\round[2] ),
    .B_N(\round[3] ),
    .X(_1330_));
 sky130_fd_sc_hd__o32a_1 _4561_ (.A1(_1308_),
    .A2(_1330_),
    .A3(_1318_),
    .B1(_1321_),
    .B2(\round[3] ),
    .X(_1331_));
 sky130_fd_sc_hd__nand2_1 _4562_ (.A(\round[3] ),
    .B(_1325_),
    .Y(_1332_));
 sky130_fd_sc_hd__o21a_1 _4563_ (.A1(\round[3] ),
    .A2(_1325_),
    .B1(_1307_),
    .X(_1333_));
 sky130_fd_sc_hd__a22o_1 _4564_ (.A1(_1329_),
    .A2(_1331_),
    .B1(_1332_),
    .B2(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__a31o_1 _4565_ (.A1(_0679_),
    .A2(_1328_),
    .A3(_1334_),
    .B1(_1317_),
    .X(_1335_));
 sky130_fd_sc_hd__o31a_1 _4566_ (.A1(_0679_),
    .A2(\round[3] ),
    .A3(net258),
    .B1(_1335_),
    .X(_0015_));
 sky130_fd_sc_hd__nor2_1 _4567_ (.A(net129),
    .B(_0672_),
    .Y(_1336_));
 sky130_fd_sc_hd__clkbuf_8 _4568_ (.A(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__clkbuf_8 _4569_ (.A(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__clkbuf_4 _4570_ (.A(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__mux2_1 _4571_ (.A0(net1),
    .A1(\mix1.data_o[0] ),
    .S(_1339_),
    .X(_1340_));
 sky130_fd_sc_hd__clkbuf_4 _4572_ (.A(_0798_),
    .X(_1341_));
 sky130_fd_sc_hd__clkbuf_4 _4573_ (.A(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__clkbuf_4 _4574_ (.A(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__clkbuf_4 _4575_ (.A(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__buf_4 _4576_ (.A(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__clkbuf_4 _4577_ (.A(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__mux2_1 _4578_ (.A0(\sub1.data_o[0] ),
    .A1(_1340_),
    .S(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__a21o_4 _4579_ (.A1(_1119_),
    .A2(_1127_),
    .B1(_0683_),
    .X(_1348_));
 sky130_fd_sc_hd__o21ai_4 _4580_ (.A1(_1124_),
    .A2(_1348_),
    .B1(state),
    .Y(_1349_));
 sky130_fd_sc_hd__buf_4 _4581_ (.A(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__a21oi_2 _4582_ (.A1(_1119_),
    .A2(_1127_),
    .B1(_0683_),
    .Y(_1351_));
 sky130_fd_sc_hd__buf_4 _4583_ (.A(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__clkbuf_4 _4584_ (.A(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__nand2_4 _4585_ (.A(_1122_),
    .B(_1351_),
    .Y(_1354_));
 sky130_fd_sc_hd__buf_4 _4586_ (.A(_1354_),
    .X(_1355_));
 sky130_fd_sc_hd__clkbuf_4 _4587_ (.A(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__a32o_1 _4588_ (.A1(\mix1.data_o[0] ),
    .A2(_1307_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[0] ),
    .X(_1357_));
 sky130_fd_sc_hd__clkbuf_8 _4589_ (.A(_0677_),
    .X(_1358_));
 sky130_fd_sc_hd__a22o_2 _4590_ (.A1(_1347_),
    .A2(_1350_),
    .B1(_1357_),
    .B2(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__buf_4 _4591_ (.A(_0675_),
    .X(_1360_));
 sky130_fd_sc_hd__mux2_1 _4592_ (.A0(\ks1.key_reg[0] ),
    .A1(net130),
    .S(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__xor2_1 _4593_ (.A(_1359_),
    .B(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__mux2_1 _4594_ (.A0(net260),
    .A1(_1362_),
    .S(next_addroundkey_ready_o),
    .X(_1363_));
 sky130_fd_sc_hd__clkbuf_1 _4595_ (.A(_1363_),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_4 _4596_ (.A(_1350_),
    .X(_1364_));
 sky130_fd_sc_hd__mux2_1 _4597_ (.A0(net40),
    .A1(\mix1.data_o[1] ),
    .S(_1339_),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_1 _4598_ (.A0(\sub1.data_o[1] ),
    .A1(_1365_),
    .S(_1346_),
    .X(_1366_));
 sky130_fd_sc_hd__a32o_1 _4599_ (.A1(\mix1.data_o[1] ),
    .A2(_1307_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[1] ),
    .X(_1367_));
 sky130_fd_sc_hd__a22o_1 _4600_ (.A1(_1364_),
    .A2(_1366_),
    .B1(_1367_),
    .B2(_1358_),
    .X(_1368_));
 sky130_fd_sc_hd__mux2_1 _4601_ (.A0(\ks1.key_reg[1] ),
    .A1(net169),
    .S(_1360_),
    .X(_1369_));
 sky130_fd_sc_hd__xor2_1 _4602_ (.A(_1368_),
    .B(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_1 _4603_ (.A0(net299),
    .A1(_1370_),
    .S(next_addroundkey_ready_o),
    .X(_1371_));
 sky130_fd_sc_hd__clkbuf_1 _4604_ (.A(_1371_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _4605_ (.A0(net51),
    .A1(\mix1.data_o[2] ),
    .S(_1339_),
    .X(_1372_));
 sky130_fd_sc_hd__mux2_1 _4606_ (.A0(\sub1.data_o[2] ),
    .A1(_1372_),
    .S(_1346_),
    .X(_1373_));
 sky130_fd_sc_hd__a32o_1 _4607_ (.A1(\mix1.data_o[2] ),
    .A2(_1307_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[2] ),
    .X(_1374_));
 sky130_fd_sc_hd__clkbuf_4 _4608_ (.A(_0677_),
    .X(_1375_));
 sky130_fd_sc_hd__a22o_1 _4609_ (.A1(_1364_),
    .A2(_1373_),
    .B1(_1374_),
    .B2(_1375_),
    .X(_1376_));
 sky130_fd_sc_hd__mux2_2 _4610_ (.A0(\ks1.key_reg[2] ),
    .A1(net180),
    .S(_1360_),
    .X(_1377_));
 sky130_fd_sc_hd__xor2_1 _4611_ (.A(_1376_),
    .B(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_1 _4612_ (.A0(net310),
    .A1(_1378_),
    .S(next_addroundkey_ready_o),
    .X(_1379_));
 sky130_fd_sc_hd__clkbuf_1 _4613_ (.A(_1379_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _4614_ (.A0(net62),
    .A1(\mix1.data_o[3] ),
    .S(_1339_),
    .X(_1380_));
 sky130_fd_sc_hd__mux2_1 _4615_ (.A0(\sub1.data_o[3] ),
    .A1(_1380_),
    .S(_1346_),
    .X(_1381_));
 sky130_fd_sc_hd__a32o_1 _4616_ (.A1(\mix1.data_o[3] ),
    .A2(_1307_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[3] ),
    .X(_1382_));
 sky130_fd_sc_hd__a22o_1 _4617_ (.A1(_1364_),
    .A2(_1381_),
    .B1(_1382_),
    .B2(_1375_),
    .X(_1383_));
 sky130_fd_sc_hd__mux2_2 _4618_ (.A0(\ks1.key_reg[3] ),
    .A1(net191),
    .S(_1360_),
    .X(_1384_));
 sky130_fd_sc_hd__xor2_1 _4619_ (.A(_1383_),
    .B(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__mux2_1 _4620_ (.A0(net321),
    .A1(_1385_),
    .S(next_addroundkey_ready_o),
    .X(_1386_));
 sky130_fd_sc_hd__clkbuf_1 _4621_ (.A(_1386_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _4622_ (.A0(net73),
    .A1(\mix1.data_o[4] ),
    .S(_1339_),
    .X(_1387_));
 sky130_fd_sc_hd__mux2_1 _4623_ (.A0(\sub1.data_o[4] ),
    .A1(_1387_),
    .S(_1346_),
    .X(_1388_));
 sky130_fd_sc_hd__a32o_1 _4624_ (.A1(\mix1.data_o[4] ),
    .A2(_1307_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[4] ),
    .X(_1389_));
 sky130_fd_sc_hd__a22o_1 _4625_ (.A1(_1364_),
    .A2(_1388_),
    .B1(_1389_),
    .B2(_1375_),
    .X(_1390_));
 sky130_fd_sc_hd__mux2_2 _4626_ (.A0(\ks1.key_reg[4] ),
    .A1(net202),
    .S(_1360_),
    .X(_1391_));
 sky130_fd_sc_hd__xor2_1 _4627_ (.A(_1390_),
    .B(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__mux2_1 _4628_ (.A0(net332),
    .A1(_1392_),
    .S(next_addroundkey_ready_o),
    .X(_1393_));
 sky130_fd_sc_hd__clkbuf_1 _4629_ (.A(_1393_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _4630_ (.A0(net84),
    .A1(\mix1.data_o[5] ),
    .S(_1339_),
    .X(_1394_));
 sky130_fd_sc_hd__mux2_1 _4631_ (.A0(\sub1.data_o[5] ),
    .A1(_1394_),
    .S(_1346_),
    .X(_1395_));
 sky130_fd_sc_hd__a32o_1 _4632_ (.A1(\mix1.data_o[5] ),
    .A2(_1307_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[5] ),
    .X(_1396_));
 sky130_fd_sc_hd__a22o_2 _4633_ (.A1(_1364_),
    .A2(_1395_),
    .B1(_1396_),
    .B2(_1375_),
    .X(_1397_));
 sky130_fd_sc_hd__mux2_1 _4634_ (.A0(\ks1.key_reg[5] ),
    .A1(net213),
    .S(_1360_),
    .X(_1398_));
 sky130_fd_sc_hd__xor2_1 _4635_ (.A(_1397_),
    .B(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__mux2_1 _4636_ (.A0(net343),
    .A1(_1399_),
    .S(next_addroundkey_ready_o),
    .X(_1400_));
 sky130_fd_sc_hd__clkbuf_1 _4637_ (.A(_1400_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _4638_ (.A0(net95),
    .A1(\mix1.data_o[6] ),
    .S(_1339_),
    .X(_1401_));
 sky130_fd_sc_hd__mux2_1 _4639_ (.A0(\sub1.data_o[6] ),
    .A1(_1401_),
    .S(_1346_),
    .X(_1402_));
 sky130_fd_sc_hd__buf_4 _4640_ (.A(_1306_),
    .X(_1403_));
 sky130_fd_sc_hd__a32o_1 _4641_ (.A1(\mix1.data_o[6] ),
    .A2(_1403_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[6] ),
    .X(_1404_));
 sky130_fd_sc_hd__a22o_1 _4642_ (.A1(_1364_),
    .A2(_1402_),
    .B1(_1404_),
    .B2(_1375_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_2 _4643_ (.A0(\ks1.key_reg[6] ),
    .A1(net224),
    .S(_1360_),
    .X(_1406_));
 sky130_fd_sc_hd__xor2_1 _4644_ (.A(_1405_),
    .B(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _4645_ (.A0(net354),
    .A1(_1407_),
    .S(next_addroundkey_ready_o),
    .X(_1408_));
 sky130_fd_sc_hd__clkbuf_1 _4646_ (.A(_1408_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _4647_ (.A0(net106),
    .A1(\mix1.data_o[7] ),
    .S(_1339_),
    .X(_1409_));
 sky130_fd_sc_hd__mux2_1 _4648_ (.A0(\sub1.data_o[7] ),
    .A1(_1409_),
    .S(_1346_),
    .X(_1410_));
 sky130_fd_sc_hd__a32o_1 _4649_ (.A1(\mix1.data_o[7] ),
    .A2(_1403_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[7] ),
    .X(_1411_));
 sky130_fd_sc_hd__a22o_1 _4650_ (.A1(_1364_),
    .A2(_1410_),
    .B1(_1411_),
    .B2(_1375_),
    .X(_1412_));
 sky130_fd_sc_hd__mux2_4 _4651_ (.A0(\ks1.key_reg[7] ),
    .A1(net235),
    .S(_1360_),
    .X(_1413_));
 sky130_fd_sc_hd__xor2_1 _4652_ (.A(_1412_),
    .B(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_1 _4653_ (.A0(net365),
    .A1(_1414_),
    .S(next_addroundkey_ready_o),
    .X(_1415_));
 sky130_fd_sc_hd__clkbuf_1 _4654_ (.A(_1415_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _4655_ (.A0(net117),
    .A1(\mix1.data_o[8] ),
    .S(_1339_),
    .X(_1416_));
 sky130_fd_sc_hd__mux2_1 _4656_ (.A0(\sub1.data_o[8] ),
    .A1(_1416_),
    .S(_1346_),
    .X(_1417_));
 sky130_fd_sc_hd__a32o_1 _4657_ (.A1(\mix1.data_o[8] ),
    .A2(_1403_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[8] ),
    .X(_1418_));
 sky130_fd_sc_hd__a22o_1 _4658_ (.A1(_1364_),
    .A2(_1417_),
    .B1(_1418_),
    .B2(_1375_),
    .X(_1419_));
 sky130_fd_sc_hd__mux2_2 _4659_ (.A0(\ks1.key_reg[8] ),
    .A1(net246),
    .S(_1360_),
    .X(_1420_));
 sky130_fd_sc_hd__xor2_1 _4660_ (.A(_1419_),
    .B(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__mux2_1 _4661_ (.A0(net376),
    .A1(_1421_),
    .S(next_addroundkey_ready_o),
    .X(_1422_));
 sky130_fd_sc_hd__clkbuf_1 _4662_ (.A(_1422_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _4663_ (.A0(net128),
    .A1(\mix1.data_o[9] ),
    .S(_1339_),
    .X(_1423_));
 sky130_fd_sc_hd__mux2_1 _4664_ (.A0(\sub1.data_o[9] ),
    .A1(_1423_),
    .S(_1346_),
    .X(_1424_));
 sky130_fd_sc_hd__a32o_1 _4665_ (.A1(\mix1.data_o[9] ),
    .A2(_1403_),
    .A3(_1353_),
    .B1(_1356_),
    .B2(\sub1.data_o[9] ),
    .X(_1425_));
 sky130_fd_sc_hd__a22o_2 _4666_ (.A1(_1364_),
    .A2(_1424_),
    .B1(_1425_),
    .B2(_1375_),
    .X(_1426_));
 sky130_fd_sc_hd__mux2_1 _4667_ (.A0(\ks1.key_reg[9] ),
    .A1(net257),
    .S(_1360_),
    .X(_1427_));
 sky130_fd_sc_hd__xor2_1 _4668_ (.A(_1426_),
    .B(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__clkbuf_8 _4669_ (.A(_0676_),
    .X(_1429_));
 sky130_fd_sc_hd__buf_4 _4670_ (.A(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__mux2_1 _4671_ (.A0(net387),
    .A1(_1428_),
    .S(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__clkbuf_1 _4672_ (.A(_1431_),
    .X(_0025_));
 sky130_fd_sc_hd__clkbuf_4 _4673_ (.A(_1338_),
    .X(_1432_));
 sky130_fd_sc_hd__mux2_1 _4674_ (.A0(net12),
    .A1(\mix1.data_o[10] ),
    .S(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__clkbuf_4 _4675_ (.A(_1345_),
    .X(_1434_));
 sky130_fd_sc_hd__mux2_1 _4676_ (.A0(\sub1.data_o[10] ),
    .A1(_1433_),
    .S(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__buf_2 _4677_ (.A(_1352_),
    .X(_1436_));
 sky130_fd_sc_hd__clkbuf_4 _4678_ (.A(_1355_),
    .X(_1437_));
 sky130_fd_sc_hd__a32o_1 _4679_ (.A1(\mix1.data_o[10] ),
    .A2(_1403_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[10] ),
    .X(_1438_));
 sky130_fd_sc_hd__a22o_1 _4680_ (.A1(_1364_),
    .A2(_1435_),
    .B1(_1438_),
    .B2(_1375_),
    .X(_1439_));
 sky130_fd_sc_hd__clkbuf_4 _4681_ (.A(_0674_),
    .X(_1440_));
 sky130_fd_sc_hd__buf_4 _4682_ (.A(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__mux2_1 _4683_ (.A0(\ks1.key_reg[10] ),
    .A1(net141),
    .S(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__xor2_1 _4684_ (.A(_1439_),
    .B(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__mux2_1 _4685_ (.A0(net271),
    .A1(_1443_),
    .S(_1430_),
    .X(_1444_));
 sky130_fd_sc_hd__clkbuf_1 _4686_ (.A(_1444_),
    .X(_0026_));
 sky130_fd_sc_hd__clkbuf_4 _4687_ (.A(_1350_),
    .X(_1445_));
 sky130_fd_sc_hd__mux2_1 _4688_ (.A0(net23),
    .A1(\mix1.data_o[11] ),
    .S(_1432_),
    .X(_1446_));
 sky130_fd_sc_hd__mux2_1 _4689_ (.A0(\sub1.data_o[11] ),
    .A1(_1446_),
    .S(_1434_),
    .X(_1447_));
 sky130_fd_sc_hd__a32o_1 _4690_ (.A1(\mix1.data_o[11] ),
    .A2(_1403_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[11] ),
    .X(_1448_));
 sky130_fd_sc_hd__a22o_1 _4691_ (.A1(_1445_),
    .A2(_1447_),
    .B1(_1448_),
    .B2(_1375_),
    .X(_1449_));
 sky130_fd_sc_hd__mux2_1 _4692_ (.A0(\ks1.key_reg[11] ),
    .A1(net152),
    .S(_1441_),
    .X(_1450_));
 sky130_fd_sc_hd__xor2_1 _4693_ (.A(_1449_),
    .B(_1450_),
    .X(_1451_));
 sky130_fd_sc_hd__mux2_1 _4694_ (.A0(net282),
    .A1(_1451_),
    .S(_1430_),
    .X(_1452_));
 sky130_fd_sc_hd__clkbuf_1 _4695_ (.A(_1452_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _4696_ (.A0(net32),
    .A1(\mix1.data_o[12] ),
    .S(_1432_),
    .X(_1453_));
 sky130_fd_sc_hd__mux2_1 _4697_ (.A0(\sub1.data_o[12] ),
    .A1(_1453_),
    .S(_1434_),
    .X(_1454_));
 sky130_fd_sc_hd__a32o_1 _4698_ (.A1(\mix1.data_o[12] ),
    .A2(_1403_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[12] ),
    .X(_1455_));
 sky130_fd_sc_hd__clkbuf_4 _4699_ (.A(_0677_),
    .X(_1456_));
 sky130_fd_sc_hd__a22o_1 _4700_ (.A1(_1445_),
    .A2(_1454_),
    .B1(_1455_),
    .B2(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__mux2_1 _4701_ (.A0(\ks1.key_reg[12] ),
    .A1(net161),
    .S(_1441_),
    .X(_1458_));
 sky130_fd_sc_hd__xor2_1 _4702_ (.A(_1457_),
    .B(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__mux2_1 _4703_ (.A0(net291),
    .A1(_1459_),
    .S(_1430_),
    .X(_1460_));
 sky130_fd_sc_hd__clkbuf_1 _4704_ (.A(_1460_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _4705_ (.A0(net33),
    .A1(\mix1.data_o[13] ),
    .S(_1432_),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_1 _4706_ (.A0(\sub1.data_o[13] ),
    .A1(_1461_),
    .S(_1434_),
    .X(_1462_));
 sky130_fd_sc_hd__a32o_1 _4707_ (.A1(\mix1.data_o[13] ),
    .A2(_1403_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[13] ),
    .X(_1463_));
 sky130_fd_sc_hd__a22o_1 _4708_ (.A1(_1445_),
    .A2(_1462_),
    .B1(_1463_),
    .B2(_1456_),
    .X(_1464_));
 sky130_fd_sc_hd__mux2_1 _4709_ (.A0(\ks1.key_reg[13] ),
    .A1(net162),
    .S(_1441_),
    .X(_1465_));
 sky130_fd_sc_hd__xor2_1 _4710_ (.A(_1464_),
    .B(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _4711_ (.A0(net292),
    .A1(_1466_),
    .S(_1430_),
    .X(_1467_));
 sky130_fd_sc_hd__clkbuf_1 _4712_ (.A(_1467_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _4713_ (.A0(net34),
    .A1(\mix1.data_o[14] ),
    .S(_1432_),
    .X(_1468_));
 sky130_fd_sc_hd__mux2_1 _4714_ (.A0(\sub1.data_o[14] ),
    .A1(_1468_),
    .S(_1434_),
    .X(_1469_));
 sky130_fd_sc_hd__a32o_1 _4715_ (.A1(\mix1.data_o[14] ),
    .A2(_1403_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[14] ),
    .X(_1470_));
 sky130_fd_sc_hd__a22o_1 _4716_ (.A1(_1445_),
    .A2(_1469_),
    .B1(_1470_),
    .B2(_1456_),
    .X(_1471_));
 sky130_fd_sc_hd__mux2_1 _4717_ (.A0(\ks1.key_reg[14] ),
    .A1(net163),
    .S(_1441_),
    .X(_1472_));
 sky130_fd_sc_hd__xor2_1 _4718_ (.A(_1471_),
    .B(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__mux2_1 _4719_ (.A0(net293),
    .A1(_1473_),
    .S(_1430_),
    .X(_1474_));
 sky130_fd_sc_hd__clkbuf_1 _4720_ (.A(_1474_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _4721_ (.A0(net35),
    .A1(\mix1.data_o[15] ),
    .S(_1432_),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_1 _4722_ (.A0(\sub1.data_o[15] ),
    .A1(_1475_),
    .S(_1434_),
    .X(_1476_));
 sky130_fd_sc_hd__a32o_1 _4723_ (.A1(\mix1.data_o[15] ),
    .A2(_1403_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[15] ),
    .X(_1477_));
 sky130_fd_sc_hd__a22o_1 _4724_ (.A1(_1445_),
    .A2(_1476_),
    .B1(_1477_),
    .B2(_1456_),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _4725_ (.A0(\ks1.key_reg[15] ),
    .A1(net164),
    .S(_1441_),
    .X(_1479_));
 sky130_fd_sc_hd__xor2_1 _4726_ (.A(_1478_),
    .B(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_1 _4727_ (.A0(net294),
    .A1(_1480_),
    .S(_1430_),
    .X(_1481_));
 sky130_fd_sc_hd__clkbuf_1 _4728_ (.A(_1481_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _4729_ (.A0(net36),
    .A1(\mix1.data_o[16] ),
    .S(_1432_),
    .X(_1482_));
 sky130_fd_sc_hd__mux2_1 _4730_ (.A0(\sub1.data_o[16] ),
    .A1(_1482_),
    .S(_1434_),
    .X(_1483_));
 sky130_fd_sc_hd__clkbuf_4 _4731_ (.A(_1306_),
    .X(_1484_));
 sky130_fd_sc_hd__a32o_1 _4732_ (.A1(\mix1.data_o[16] ),
    .A2(_1484_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[16] ),
    .X(_1485_));
 sky130_fd_sc_hd__a22o_1 _4733_ (.A1(_1445_),
    .A2(_1483_),
    .B1(_1485_),
    .B2(_1456_),
    .X(_1486_));
 sky130_fd_sc_hd__mux2_1 _4734_ (.A0(\ks1.key_reg[16] ),
    .A1(net165),
    .S(_1441_),
    .X(_1487_));
 sky130_fd_sc_hd__xor2_1 _4735_ (.A(_1486_),
    .B(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__mux2_1 _4736_ (.A0(net295),
    .A1(_1488_),
    .S(_1430_),
    .X(_1489_));
 sky130_fd_sc_hd__clkbuf_1 _4737_ (.A(_1489_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _4738_ (.A0(net37),
    .A1(\mix1.data_o[17] ),
    .S(_1432_),
    .X(_1490_));
 sky130_fd_sc_hd__mux2_1 _4739_ (.A0(\sub1.data_o[17] ),
    .A1(_1490_),
    .S(_1434_),
    .X(_1491_));
 sky130_fd_sc_hd__a32o_1 _4740_ (.A1(\mix1.data_o[17] ),
    .A2(_1484_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[17] ),
    .X(_1492_));
 sky130_fd_sc_hd__a22o_1 _4741_ (.A1(_1445_),
    .A2(_1491_),
    .B1(_1492_),
    .B2(_1456_),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_1 _4742_ (.A0(\ks1.key_reg[17] ),
    .A1(net166),
    .S(_1441_),
    .X(_1494_));
 sky130_fd_sc_hd__xor2_1 _4743_ (.A(_1493_),
    .B(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_1 _4744_ (.A0(net296),
    .A1(_1495_),
    .S(_1430_),
    .X(_1496_));
 sky130_fd_sc_hd__clkbuf_1 _4745_ (.A(_1496_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _4746_ (.A0(net38),
    .A1(\mix1.data_o[18] ),
    .S(_1432_),
    .X(_1497_));
 sky130_fd_sc_hd__mux2_1 _4747_ (.A0(\sub1.data_o[18] ),
    .A1(_1497_),
    .S(_1434_),
    .X(_1498_));
 sky130_fd_sc_hd__a32o_1 _4748_ (.A1(\mix1.data_o[18] ),
    .A2(_1484_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[18] ),
    .X(_1499_));
 sky130_fd_sc_hd__a22o_1 _4749_ (.A1(_1445_),
    .A2(_1498_),
    .B1(_1499_),
    .B2(_1456_),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_1 _4750_ (.A0(\ks1.key_reg[18] ),
    .A1(net167),
    .S(_1441_),
    .X(_1501_));
 sky130_fd_sc_hd__xor2_1 _4751_ (.A(_1500_),
    .B(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__mux2_1 _4752_ (.A0(net297),
    .A1(_1502_),
    .S(_1430_),
    .X(_1503_));
 sky130_fd_sc_hd__clkbuf_1 _4753_ (.A(_1503_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _4754_ (.A0(net39),
    .A1(\mix1.data_o[19] ),
    .S(_1432_),
    .X(_1504_));
 sky130_fd_sc_hd__mux2_1 _4755_ (.A0(\sub1.data_o[19] ),
    .A1(_1504_),
    .S(_1434_),
    .X(_1505_));
 sky130_fd_sc_hd__a32o_1 _4756_ (.A1(\mix1.data_o[19] ),
    .A2(_1484_),
    .A3(_1436_),
    .B1(_1437_),
    .B2(\sub1.data_o[19] ),
    .X(_1506_));
 sky130_fd_sc_hd__a22o_1 _4757_ (.A1(_1445_),
    .A2(_1505_),
    .B1(_1506_),
    .B2(_1456_),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _4758_ (.A0(\ks1.key_reg[19] ),
    .A1(net168),
    .S(_1441_),
    .X(_1508_));
 sky130_fd_sc_hd__xor2_1 _4759_ (.A(_1507_),
    .B(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__buf_4 _4760_ (.A(_0676_),
    .X(_1510_));
 sky130_fd_sc_hd__buf_4 _4761_ (.A(_1510_),
    .X(_1511_));
 sky130_fd_sc_hd__mux2_1 _4762_ (.A0(net298),
    .A1(_1509_),
    .S(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__clkbuf_1 _4763_ (.A(_1512_),
    .X(_0035_));
 sky130_fd_sc_hd__clkbuf_8 _4764_ (.A(_1336_),
    .X(_1513_));
 sky130_fd_sc_hd__buf_4 _4765_ (.A(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__mux2_1 _4766_ (.A0(net41),
    .A1(\mix1.data_o[20] ),
    .S(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__clkbuf_8 _4767_ (.A(_1343_),
    .X(_1516_));
 sky130_fd_sc_hd__buf_4 _4768_ (.A(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _4769_ (.A0(\sub1.data_o[20] ),
    .A1(_1515_),
    .S(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__buf_4 _4770_ (.A(_1351_),
    .X(_1519_));
 sky130_fd_sc_hd__clkbuf_4 _4771_ (.A(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__clkbuf_4 _4772_ (.A(_1354_),
    .X(_1521_));
 sky130_fd_sc_hd__a32o_1 _4773_ (.A1(\mix1.data_o[20] ),
    .A2(_1484_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[20] ),
    .X(_1522_));
 sky130_fd_sc_hd__a22o_1 _4774_ (.A1(_1445_),
    .A2(_1518_),
    .B1(_1522_),
    .B2(_1456_),
    .X(_1523_));
 sky130_fd_sc_hd__buf_4 _4775_ (.A(_1440_),
    .X(_1524_));
 sky130_fd_sc_hd__mux2_1 _4776_ (.A0(\ks1.key_reg[20] ),
    .A1(net170),
    .S(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__xor2_1 _4777_ (.A(_1523_),
    .B(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__mux2_1 _4778_ (.A0(net300),
    .A1(_1526_),
    .S(_1511_),
    .X(_1527_));
 sky130_fd_sc_hd__clkbuf_1 _4779_ (.A(_1527_),
    .X(_0036_));
 sky130_fd_sc_hd__clkbuf_4 _4780_ (.A(_1349_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _4781_ (.A0(net42),
    .A1(\mix1.data_o[21] ),
    .S(_1514_),
    .X(_1529_));
 sky130_fd_sc_hd__mux2_1 _4782_ (.A0(\sub1.data_o[21] ),
    .A1(_1529_),
    .S(_1517_),
    .X(_1530_));
 sky130_fd_sc_hd__a32o_1 _4783_ (.A1(\mix1.data_o[21] ),
    .A2(_1484_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[21] ),
    .X(_1531_));
 sky130_fd_sc_hd__a22o_1 _4784_ (.A1(_1528_),
    .A2(_1530_),
    .B1(_1531_),
    .B2(_1456_),
    .X(_1532_));
 sky130_fd_sc_hd__mux2_1 _4785_ (.A0(\ks1.key_reg[21] ),
    .A1(net171),
    .S(_1524_),
    .X(_1533_));
 sky130_fd_sc_hd__xor2_1 _4786_ (.A(_1532_),
    .B(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__mux2_1 _4787_ (.A0(net301),
    .A1(_1534_),
    .S(_1511_),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _4788_ (.A(_1535_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _4789_ (.A0(net43),
    .A1(\mix1.data_o[22] ),
    .S(_1514_),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _4790_ (.A0(\sub1.data_o[22] ),
    .A1(_1536_),
    .S(_1517_),
    .X(_1537_));
 sky130_fd_sc_hd__a32o_1 _4791_ (.A1(\mix1.data_o[22] ),
    .A2(_1484_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[22] ),
    .X(_1538_));
 sky130_fd_sc_hd__clkbuf_4 _4792_ (.A(_0677_),
    .X(_1539_));
 sky130_fd_sc_hd__a22o_1 _4793_ (.A1(_1528_),
    .A2(_1537_),
    .B1(_1538_),
    .B2(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _4794_ (.A0(\ks1.key_reg[22] ),
    .A1(net172),
    .S(_1524_),
    .X(_1541_));
 sky130_fd_sc_hd__xor2_1 _4795_ (.A(_1540_),
    .B(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__mux2_1 _4796_ (.A0(net302),
    .A1(_1542_),
    .S(_1511_),
    .X(_1543_));
 sky130_fd_sc_hd__clkbuf_1 _4797_ (.A(_1543_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _4798_ (.A0(net44),
    .A1(\mix1.data_o[23] ),
    .S(_1514_),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _4799_ (.A0(\sub1.data_o[23] ),
    .A1(_1544_),
    .S(_1517_),
    .X(_1545_));
 sky130_fd_sc_hd__a32o_1 _4800_ (.A1(\mix1.data_o[23] ),
    .A2(_1484_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[23] ),
    .X(_1546_));
 sky130_fd_sc_hd__a22o_1 _4801_ (.A1(_1528_),
    .A2(_1545_),
    .B1(_1546_),
    .B2(_1539_),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_1 _4802_ (.A0(\ks1.key_reg[23] ),
    .A1(net173),
    .S(_1524_),
    .X(_1548_));
 sky130_fd_sc_hd__xor2_1 _4803_ (.A(_1547_),
    .B(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__mux2_1 _4804_ (.A0(net303),
    .A1(_1549_),
    .S(_1511_),
    .X(_1550_));
 sky130_fd_sc_hd__clkbuf_1 _4805_ (.A(_1550_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _4806_ (.A0(net45),
    .A1(\mix1.data_o[24] ),
    .S(_1514_),
    .X(_1551_));
 sky130_fd_sc_hd__mux2_1 _4807_ (.A0(\sub1.data_o[24] ),
    .A1(_1551_),
    .S(_1517_),
    .X(_1552_));
 sky130_fd_sc_hd__a32o_1 _4808_ (.A1(\mix1.data_o[24] ),
    .A2(_1484_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[24] ),
    .X(_1553_));
 sky130_fd_sc_hd__a22o_1 _4809_ (.A1(_1528_),
    .A2(_1552_),
    .B1(_1553_),
    .B2(_1539_),
    .X(_1554_));
 sky130_fd_sc_hd__mux2_1 _4810_ (.A0(\ks1.key_reg[24] ),
    .A1(net174),
    .S(_1524_),
    .X(_1555_));
 sky130_fd_sc_hd__xor2_1 _4811_ (.A(_1554_),
    .B(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__mux2_1 _4812_ (.A0(net304),
    .A1(_1556_),
    .S(_1511_),
    .X(_1557_));
 sky130_fd_sc_hd__clkbuf_1 _4813_ (.A(_1557_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _4814_ (.A0(net46),
    .A1(\mix1.data_o[25] ),
    .S(_1514_),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_1 _4815_ (.A0(\sub1.data_o[25] ),
    .A1(_1558_),
    .S(_1517_),
    .X(_1559_));
 sky130_fd_sc_hd__a32o_1 _4816_ (.A1(\mix1.data_o[25] ),
    .A2(_1484_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[25] ),
    .X(_1560_));
 sky130_fd_sc_hd__a22o_1 _4817_ (.A1(_1528_),
    .A2(_1559_),
    .B1(_1560_),
    .B2(_1539_),
    .X(_1561_));
 sky130_fd_sc_hd__mux2_1 _4818_ (.A0(\ks1.key_reg[25] ),
    .A1(net175),
    .S(_1524_),
    .X(_1562_));
 sky130_fd_sc_hd__xor2_1 _4819_ (.A(_1561_),
    .B(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__mux2_1 _4820_ (.A0(net305),
    .A1(_1563_),
    .S(_1511_),
    .X(_1564_));
 sky130_fd_sc_hd__clkbuf_1 _4821_ (.A(_1564_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(net47),
    .A1(\mix1.data_o[26] ),
    .S(_1514_),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_1 _4823_ (.A0(\sub1.data_o[26] ),
    .A1(_1565_),
    .S(_1517_),
    .X(_1566_));
 sky130_fd_sc_hd__clkbuf_4 _4824_ (.A(_1306_),
    .X(_1567_));
 sky130_fd_sc_hd__a32o_1 _4825_ (.A1(\mix1.data_o[26] ),
    .A2(_1567_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[26] ),
    .X(_1568_));
 sky130_fd_sc_hd__a22o_1 _4826_ (.A1(_1528_),
    .A2(_1566_),
    .B1(_1568_),
    .B2(_1539_),
    .X(_1569_));
 sky130_fd_sc_hd__mux2_1 _4827_ (.A0(\ks1.key_reg[26] ),
    .A1(net176),
    .S(_1524_),
    .X(_1570_));
 sky130_fd_sc_hd__xor2_1 _4828_ (.A(_1569_),
    .B(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__mux2_1 _4829_ (.A0(net306),
    .A1(_1571_),
    .S(_1511_),
    .X(_1572_));
 sky130_fd_sc_hd__clkbuf_1 _4830_ (.A(_1572_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _4831_ (.A0(net48),
    .A1(\mix1.data_o[27] ),
    .S(_1514_),
    .X(_1573_));
 sky130_fd_sc_hd__mux2_1 _4832_ (.A0(\sub1.data_o[27] ),
    .A1(_1573_),
    .S(_1517_),
    .X(_1574_));
 sky130_fd_sc_hd__a32o_1 _4833_ (.A1(\mix1.data_o[27] ),
    .A2(_1567_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[27] ),
    .X(_1575_));
 sky130_fd_sc_hd__a22o_1 _4834_ (.A1(_1528_),
    .A2(_1574_),
    .B1(_1575_),
    .B2(_1539_),
    .X(_1576_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(\ks1.key_reg[27] ),
    .A1(net177),
    .S(_1524_),
    .X(_1577_));
 sky130_fd_sc_hd__xor2_1 _4836_ (.A(_1576_),
    .B(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__mux2_1 _4837_ (.A0(net307),
    .A1(_1578_),
    .S(_1511_),
    .X(_1579_));
 sky130_fd_sc_hd__clkbuf_1 _4838_ (.A(_1579_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _4839_ (.A0(net49),
    .A1(\mix1.data_o[28] ),
    .S(_1514_),
    .X(_1580_));
 sky130_fd_sc_hd__mux2_1 _4840_ (.A0(\sub1.data_o[28] ),
    .A1(_1580_),
    .S(_1517_),
    .X(_1581_));
 sky130_fd_sc_hd__a32o_1 _4841_ (.A1(\mix1.data_o[28] ),
    .A2(_1567_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[28] ),
    .X(_1582_));
 sky130_fd_sc_hd__a22o_1 _4842_ (.A1(_1528_),
    .A2(_1581_),
    .B1(_1582_),
    .B2(_1539_),
    .X(_1583_));
 sky130_fd_sc_hd__mux2_1 _4843_ (.A0(\ks1.key_reg[28] ),
    .A1(net178),
    .S(_1524_),
    .X(_1584_));
 sky130_fd_sc_hd__xor2_1 _4844_ (.A(_1583_),
    .B(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__mux2_1 _4845_ (.A0(net308),
    .A1(_1585_),
    .S(_1511_),
    .X(_1586_));
 sky130_fd_sc_hd__clkbuf_1 _4846_ (.A(_1586_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _4847_ (.A0(net50),
    .A1(\mix1.data_o[29] ),
    .S(_1514_),
    .X(_1587_));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(\sub1.data_o[29] ),
    .A1(_1587_),
    .S(_1517_),
    .X(_1588_));
 sky130_fd_sc_hd__a32o_1 _4849_ (.A1(\mix1.data_o[29] ),
    .A2(_1567_),
    .A3(_1520_),
    .B1(_1521_),
    .B2(\sub1.data_o[29] ),
    .X(_1589_));
 sky130_fd_sc_hd__a22o_1 _4850_ (.A1(_1528_),
    .A2(_1588_),
    .B1(_1589_),
    .B2(_1539_),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_1 _4851_ (.A0(\ks1.key_reg[29] ),
    .A1(net179),
    .S(_1524_),
    .X(_1591_));
 sky130_fd_sc_hd__xor2_1 _4852_ (.A(_1590_),
    .B(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__buf_8 _4853_ (.A(_1510_),
    .X(_1593_));
 sky130_fd_sc_hd__mux2_1 _4854_ (.A0(net309),
    .A1(_1592_),
    .S(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__clkbuf_1 _4855_ (.A(_1594_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_4 _4856_ (.A(_1513_),
    .X(_1595_));
 sky130_fd_sc_hd__mux2_1 _4857_ (.A0(net52),
    .A1(\mix1.data_o[30] ),
    .S(_1595_),
    .X(_1596_));
 sky130_fd_sc_hd__clkbuf_4 _4858_ (.A(_1516_),
    .X(_1597_));
 sky130_fd_sc_hd__mux2_1 _4859_ (.A0(\sub1.data_o[30] ),
    .A1(_1596_),
    .S(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__clkbuf_4 _4860_ (.A(_1519_),
    .X(_1599_));
 sky130_fd_sc_hd__clkbuf_4 _4861_ (.A(_1354_),
    .X(_1600_));
 sky130_fd_sc_hd__a32o_1 _4862_ (.A1(\mix1.data_o[30] ),
    .A2(_1567_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[30] ),
    .X(_1601_));
 sky130_fd_sc_hd__a22o_1 _4863_ (.A1(_1528_),
    .A2(_1598_),
    .B1(_1601_),
    .B2(_1539_),
    .X(_1602_));
 sky130_fd_sc_hd__buf_4 _4864_ (.A(_1440_),
    .X(_1603_));
 sky130_fd_sc_hd__mux2_1 _4865_ (.A0(\ks1.key_reg[30] ),
    .A1(net181),
    .S(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__xor2_1 _4866_ (.A(_1602_),
    .B(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__mux2_1 _4867_ (.A0(net311),
    .A1(_1605_),
    .S(_1593_),
    .X(_1606_));
 sky130_fd_sc_hd__clkbuf_1 _4868_ (.A(_1606_),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_4 _4869_ (.A(_1349_),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_1 _4870_ (.A0(net53),
    .A1(\mix1.data_o[31] ),
    .S(_1595_),
    .X(_1608_));
 sky130_fd_sc_hd__mux2_1 _4871_ (.A0(\sub1.data_o[31] ),
    .A1(_1608_),
    .S(_1597_),
    .X(_1609_));
 sky130_fd_sc_hd__a32o_1 _4872_ (.A1(\mix1.data_o[31] ),
    .A2(_1567_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[31] ),
    .X(_1610_));
 sky130_fd_sc_hd__a22o_1 _4873_ (.A1(_1607_),
    .A2(_1609_),
    .B1(_1610_),
    .B2(_1539_),
    .X(_1611_));
 sky130_fd_sc_hd__mux2_1 _4874_ (.A0(\ks1.key_reg[31] ),
    .A1(net182),
    .S(_1603_),
    .X(_1612_));
 sky130_fd_sc_hd__xor2_1 _4875_ (.A(_1611_),
    .B(_1612_),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_1 _4876_ (.A0(net312),
    .A1(_1613_),
    .S(_1593_),
    .X(_1614_));
 sky130_fd_sc_hd__clkbuf_1 _4877_ (.A(_1614_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(net54),
    .A1(\mix1.data_o[32] ),
    .S(_1513_),
    .X(_1615_));
 sky130_fd_sc_hd__mux2_1 _4879_ (.A0(\sub1.data_o[32] ),
    .A1(_1615_),
    .S(_1516_),
    .X(_1616_));
 sky130_fd_sc_hd__buf_4 _4880_ (.A(_1348_),
    .X(_1617_));
 sky130_fd_sc_hd__clkbuf_4 _4881_ (.A(_1305_),
    .X(_1618_));
 sky130_fd_sc_hd__a31o_1 _4882_ (.A1(_1217_),
    .A2(\sub1.data_o[32] ),
    .A3(_1120_),
    .B1(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__a21o_1 _4883_ (.A1(_1318_),
    .A2(_1616_),
    .B1(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__clkbuf_4 _4884_ (.A(_1519_),
    .X(_1621_));
 sky130_fd_sc_hd__o21a_1 _4885_ (.A1(\mix1.data_o[32] ),
    .A2(_1329_),
    .B1(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__a221o_1 _4886_ (.A1(\sub1.data_o[32] ),
    .A2(_1617_),
    .B1(_1620_),
    .B2(_1622_),
    .C1(_1115_),
    .X(_1623_));
 sky130_fd_sc_hd__o21ai_1 _4887_ (.A1(_0679_),
    .A2(_1616_),
    .B1(_1623_),
    .Y(_1624_));
 sky130_fd_sc_hd__buf_4 _4888_ (.A(_1440_),
    .X(_1625_));
 sky130_fd_sc_hd__mux2_2 _4889_ (.A0(\ks1.key_reg[32] ),
    .A1(net183),
    .S(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__xnor2_1 _4890_ (.A(_1624_),
    .B(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__mux2_1 _4891_ (.A0(net313),
    .A1(_1627_),
    .S(_1593_),
    .X(_1628_));
 sky130_fd_sc_hd__clkbuf_1 _4892_ (.A(_1628_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _4893_ (.A0(net55),
    .A1(\mix1.data_o[33] ),
    .S(_1513_),
    .X(_1629_));
 sky130_fd_sc_hd__mux2_1 _4894_ (.A0(\sub1.data_o[33] ),
    .A1(_1629_),
    .S(_1516_),
    .X(_1630_));
 sky130_fd_sc_hd__a31o_1 _4895_ (.A1(_1217_),
    .A2(\sub1.data_o[33] ),
    .A3(_1120_),
    .B1(_1618_),
    .X(_1631_));
 sky130_fd_sc_hd__a21o_1 _4896_ (.A1(_1318_),
    .A2(_1630_),
    .B1(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__o21a_1 _4897_ (.A1(\mix1.data_o[33] ),
    .A2(_1329_),
    .B1(_1621_),
    .X(_1633_));
 sky130_fd_sc_hd__a221o_1 _4898_ (.A1(\sub1.data_o[33] ),
    .A2(_1617_),
    .B1(_1632_),
    .B2(_1633_),
    .C1(_1115_),
    .X(_1634_));
 sky130_fd_sc_hd__o21ai_4 _4899_ (.A1(_0679_),
    .A2(_1630_),
    .B1(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__mux2_1 _4900_ (.A0(\ks1.key_reg[33] ),
    .A1(net184),
    .S(_1625_),
    .X(_1636_));
 sky130_fd_sc_hd__xnor2_1 _4901_ (.A(_1635_),
    .B(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__mux2_1 _4902_ (.A0(net314),
    .A1(_1637_),
    .S(_1593_),
    .X(_1638_));
 sky130_fd_sc_hd__clkbuf_1 _4903_ (.A(_1638_),
    .X(_0049_));
 sky130_fd_sc_hd__buf_4 _4904_ (.A(_0678_),
    .X(_1639_));
 sky130_fd_sc_hd__mux2_1 _4905_ (.A0(net56),
    .A1(\mix1.data_o[34] ),
    .S(_1513_),
    .X(_1640_));
 sky130_fd_sc_hd__mux2_1 _4906_ (.A0(\sub1.data_o[34] ),
    .A1(_1640_),
    .S(_1516_),
    .X(_1641_));
 sky130_fd_sc_hd__a31o_1 _4907_ (.A1(_1217_),
    .A2(\sub1.data_o[34] ),
    .A3(_1120_),
    .B1(_1618_),
    .X(_1642_));
 sky130_fd_sc_hd__a21o_1 _4908_ (.A1(_1318_),
    .A2(_1641_),
    .B1(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__clkbuf_4 _4909_ (.A(_1519_),
    .X(_1644_));
 sky130_fd_sc_hd__o21a_1 _4910_ (.A1(\mix1.data_o[34] ),
    .A2(_1329_),
    .B1(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__a221o_1 _4911_ (.A1(\sub1.data_o[34] ),
    .A2(_1617_),
    .B1(_1643_),
    .B2(_1645_),
    .C1(_1115_),
    .X(_1646_));
 sky130_fd_sc_hd__o21ai_2 _4912_ (.A1(_1639_),
    .A2(_1641_),
    .B1(_1646_),
    .Y(_1647_));
 sky130_fd_sc_hd__buf_4 _4913_ (.A(_1440_),
    .X(_1648_));
 sky130_fd_sc_hd__mux2_2 _4914_ (.A0(\ks1.key_reg[34] ),
    .A1(net185),
    .S(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__xnor2_1 _4915_ (.A(_1647_),
    .B(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__mux2_1 _4916_ (.A0(net315),
    .A1(_1650_),
    .S(_1593_),
    .X(_1651_));
 sky130_fd_sc_hd__clkbuf_1 _4917_ (.A(_1651_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _4918_ (.A0(net57),
    .A1(\mix1.data_o[35] ),
    .S(_1513_),
    .X(_1652_));
 sky130_fd_sc_hd__mux2_1 _4919_ (.A0(\sub1.data_o[35] ),
    .A1(_1652_),
    .S(_1516_),
    .X(_1653_));
 sky130_fd_sc_hd__a31o_1 _4920_ (.A1(_1217_),
    .A2(\sub1.data_o[35] ),
    .A3(_1120_),
    .B1(_1618_),
    .X(_1654_));
 sky130_fd_sc_hd__a21o_1 _4921_ (.A1(_1318_),
    .A2(_1653_),
    .B1(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__o21a_1 _4922_ (.A1(\mix1.data_o[35] ),
    .A2(_1329_),
    .B1(_1644_),
    .X(_1656_));
 sky130_fd_sc_hd__a221o_1 _4923_ (.A1(\sub1.data_o[35] ),
    .A2(_1617_),
    .B1(_1655_),
    .B2(_1656_),
    .C1(_1115_),
    .X(_1657_));
 sky130_fd_sc_hd__o21ai_1 _4924_ (.A1(_1639_),
    .A2(_1653_),
    .B1(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hd__mux2_2 _4925_ (.A0(\ks1.key_reg[35] ),
    .A1(net186),
    .S(_1648_),
    .X(_1659_));
 sky130_fd_sc_hd__xnor2_1 _4926_ (.A(_1658_),
    .B(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__mux2_1 _4927_ (.A0(net316),
    .A1(_1660_),
    .S(_1593_),
    .X(_1661_));
 sky130_fd_sc_hd__clkbuf_1 _4928_ (.A(_1661_),
    .X(_0051_));
 sky130_fd_sc_hd__clkbuf_4 _4929_ (.A(_1337_),
    .X(_1662_));
 sky130_fd_sc_hd__mux2_1 _4930_ (.A0(net58),
    .A1(\mix1.data_o[36] ),
    .S(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__clkbuf_4 _4931_ (.A(_1344_),
    .X(_1664_));
 sky130_fd_sc_hd__mux2_1 _4932_ (.A0(\sub1.data_o[36] ),
    .A1(_1663_),
    .S(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__clkbuf_4 _4933_ (.A(_1119_),
    .X(_1666_));
 sky130_fd_sc_hd__a31o_1 _4934_ (.A1(_1217_),
    .A2(\sub1.data_o[36] ),
    .A3(_1666_),
    .B1(_1618_),
    .X(_1667_));
 sky130_fd_sc_hd__a21o_1 _4935_ (.A1(_1318_),
    .A2(_1665_),
    .B1(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__o21a_1 _4936_ (.A1(\mix1.data_o[36] ),
    .A2(_1329_),
    .B1(_1644_),
    .X(_1669_));
 sky130_fd_sc_hd__a221o_1 _4937_ (.A1(\sub1.data_o[36] ),
    .A2(_1617_),
    .B1(_1668_),
    .B2(_1669_),
    .C1(_1115_),
    .X(_1670_));
 sky130_fd_sc_hd__o21ai_4 _4938_ (.A1(_1639_),
    .A2(_1665_),
    .B1(_1670_),
    .Y(_1671_));
 sky130_fd_sc_hd__mux2_2 _4939_ (.A0(\ks1.key_reg[36] ),
    .A1(net187),
    .S(_1648_),
    .X(_1672_));
 sky130_fd_sc_hd__xnor2_1 _4940_ (.A(_1671_),
    .B(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__mux2_1 _4941_ (.A0(net317),
    .A1(_1673_),
    .S(_1593_),
    .X(_1674_));
 sky130_fd_sc_hd__clkbuf_1 _4942_ (.A(_1674_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _4943_ (.A0(net59),
    .A1(\mix1.data_o[37] ),
    .S(_1662_),
    .X(_1675_));
 sky130_fd_sc_hd__mux2_1 _4944_ (.A0(\sub1.data_o[37] ),
    .A1(_1675_),
    .S(_1664_),
    .X(_1676_));
 sky130_fd_sc_hd__clkbuf_4 _4945_ (.A(_1121_),
    .X(_1677_));
 sky130_fd_sc_hd__a31o_1 _4946_ (.A1(\sub1.data_o[37] ),
    .A2(_1677_),
    .A3(_1666_),
    .B1(_1618_),
    .X(_1678_));
 sky130_fd_sc_hd__a21o_1 _4947_ (.A1(_1318_),
    .A2(_1676_),
    .B1(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__o21a_1 _4948_ (.A1(\mix1.data_o[37] ),
    .A2(_1329_),
    .B1(_1644_),
    .X(_1680_));
 sky130_fd_sc_hd__a221o_1 _4949_ (.A1(\sub1.data_o[37] ),
    .A2(_1617_),
    .B1(_1679_),
    .B2(_1680_),
    .C1(_1115_),
    .X(_1681_));
 sky130_fd_sc_hd__o21ai_1 _4950_ (.A1(_1639_),
    .A2(_1676_),
    .B1(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__mux2_4 _4951_ (.A0(\ks1.key_reg[37] ),
    .A1(net188),
    .S(_1648_),
    .X(_1683_));
 sky130_fd_sc_hd__xnor2_1 _4952_ (.A(_1682_),
    .B(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__mux2_1 _4953_ (.A0(net318),
    .A1(_1684_),
    .S(_1593_),
    .X(_1685_));
 sky130_fd_sc_hd__clkbuf_1 _4954_ (.A(_1685_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _4955_ (.A0(net60),
    .A1(\mix1.data_o[38] ),
    .S(_1662_),
    .X(_1686_));
 sky130_fd_sc_hd__mux2_1 _4956_ (.A0(\sub1.data_o[38] ),
    .A1(_1686_),
    .S(_1664_),
    .X(_1687_));
 sky130_fd_sc_hd__clkbuf_4 _4957_ (.A(_1122_),
    .X(_1688_));
 sky130_fd_sc_hd__a31o_1 _4958_ (.A1(\sub1.data_o[38] ),
    .A2(_1677_),
    .A3(_1666_),
    .B1(_1618_),
    .X(_1689_));
 sky130_fd_sc_hd__a21o_1 _4959_ (.A1(_1688_),
    .A2(_1687_),
    .B1(_1689_),
    .X(_1690_));
 sky130_fd_sc_hd__o21a_1 _4960_ (.A1(\mix1.data_o[38] ),
    .A2(_1329_),
    .B1(_1644_),
    .X(_1691_));
 sky130_fd_sc_hd__a221o_1 _4961_ (.A1(\sub1.data_o[38] ),
    .A2(_1617_),
    .B1(_1690_),
    .B2(_1691_),
    .C1(_1115_),
    .X(_1692_));
 sky130_fd_sc_hd__o21ai_1 _4962_ (.A1(_1639_),
    .A2(_1687_),
    .B1(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__mux2_2 _4963_ (.A0(\ks1.key_reg[38] ),
    .A1(net189),
    .S(_1648_),
    .X(_1694_));
 sky130_fd_sc_hd__xnor2_1 _4964_ (.A(_1693_),
    .B(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__mux2_1 _4965_ (.A0(net319),
    .A1(_1695_),
    .S(_1593_),
    .X(_1696_));
 sky130_fd_sc_hd__clkbuf_1 _4966_ (.A(_1696_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _4967_ (.A0(net61),
    .A1(\mix1.data_o[39] ),
    .S(_1662_),
    .X(_1697_));
 sky130_fd_sc_hd__mux2_1 _4968_ (.A0(\sub1.data_o[39] ),
    .A1(_1697_),
    .S(_1664_),
    .X(_1698_));
 sky130_fd_sc_hd__a31o_1 _4969_ (.A1(\sub1.data_o[39] ),
    .A2(_1677_),
    .A3(_1666_),
    .B1(_1618_),
    .X(_1699_));
 sky130_fd_sc_hd__a21o_1 _4970_ (.A1(_1688_),
    .A2(_1698_),
    .B1(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__o21a_1 _4971_ (.A1(\mix1.data_o[39] ),
    .A2(_1329_),
    .B1(_1644_),
    .X(_1701_));
 sky130_fd_sc_hd__clkbuf_4 _4972_ (.A(_1114_),
    .X(_1702_));
 sky130_fd_sc_hd__a221o_1 _4973_ (.A1(\sub1.data_o[39] ),
    .A2(_1617_),
    .B1(_1700_),
    .B2(_1701_),
    .C1(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__o21ai_2 _4974_ (.A1(_1639_),
    .A2(_1698_),
    .B1(_1703_),
    .Y(_1704_));
 sky130_fd_sc_hd__mux2_1 _4975_ (.A0(\ks1.key_reg[39] ),
    .A1(net190),
    .S(_1648_),
    .X(_1705_));
 sky130_fd_sc_hd__xnor2_1 _4976_ (.A(_1704_),
    .B(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__buf_4 _4977_ (.A(_1510_),
    .X(_1707_));
 sky130_fd_sc_hd__mux2_1 _4978_ (.A0(net320),
    .A1(_1706_),
    .S(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__clkbuf_1 _4979_ (.A(_1708_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _4980_ (.A0(net63),
    .A1(\mix1.data_o[40] ),
    .S(_1595_),
    .X(_1709_));
 sky130_fd_sc_hd__mux2_1 _4981_ (.A0(\sub1.data_o[40] ),
    .A1(_1709_),
    .S(_1597_),
    .X(_1710_));
 sky130_fd_sc_hd__a32o_1 _4982_ (.A1(\mix1.data_o[40] ),
    .A2(_1567_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[40] ),
    .X(_1711_));
 sky130_fd_sc_hd__clkbuf_4 _4983_ (.A(_0677_),
    .X(_1712_));
 sky130_fd_sc_hd__a22o_1 _4984_ (.A1(_1607_),
    .A2(_1710_),
    .B1(_1711_),
    .B2(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__mux2_1 _4985_ (.A0(\ks1.key_reg[40] ),
    .A1(net192),
    .S(_1603_),
    .X(_1714_));
 sky130_fd_sc_hd__xor2_1 _4986_ (.A(_1713_),
    .B(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__mux2_1 _4987_ (.A0(net322),
    .A1(_1715_),
    .S(_1707_),
    .X(_1716_));
 sky130_fd_sc_hd__clkbuf_1 _4988_ (.A(_1716_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _4989_ (.A0(net64),
    .A1(\mix1.data_o[41] ),
    .S(_1595_),
    .X(_1717_));
 sky130_fd_sc_hd__mux2_1 _4990_ (.A0(\sub1.data_o[41] ),
    .A1(_1717_),
    .S(_1597_),
    .X(_1718_));
 sky130_fd_sc_hd__a32o_1 _4991_ (.A1(\mix1.data_o[41] ),
    .A2(_1567_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[41] ),
    .X(_1719_));
 sky130_fd_sc_hd__a22o_1 _4992_ (.A1(_1607_),
    .A2(_1718_),
    .B1(_1719_),
    .B2(_1712_),
    .X(_1720_));
 sky130_fd_sc_hd__mux2_2 _4993_ (.A0(\ks1.key_reg[41] ),
    .A1(net193),
    .S(_1603_),
    .X(_1721_));
 sky130_fd_sc_hd__xor2_1 _4994_ (.A(_1720_),
    .B(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__mux2_1 _4995_ (.A0(net323),
    .A1(_1722_),
    .S(_1707_),
    .X(_1723_));
 sky130_fd_sc_hd__clkbuf_1 _4996_ (.A(_1723_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _4997_ (.A0(net65),
    .A1(\mix1.data_o[42] ),
    .S(_1595_),
    .X(_1724_));
 sky130_fd_sc_hd__mux2_1 _4998_ (.A0(\sub1.data_o[42] ),
    .A1(_1724_),
    .S(_1597_),
    .X(_1725_));
 sky130_fd_sc_hd__a32o_1 _4999_ (.A1(\mix1.data_o[42] ),
    .A2(_1567_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[42] ),
    .X(_1726_));
 sky130_fd_sc_hd__a22o_1 _5000_ (.A1(_1607_),
    .A2(_1725_),
    .B1(_1726_),
    .B2(_1712_),
    .X(_1727_));
 sky130_fd_sc_hd__mux2_1 _5001_ (.A0(\ks1.key_reg[42] ),
    .A1(net194),
    .S(_1603_),
    .X(_1728_));
 sky130_fd_sc_hd__xor2_1 _5002_ (.A(_1727_),
    .B(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__mux2_1 _5003_ (.A0(net324),
    .A1(_1729_),
    .S(_1707_),
    .X(_1730_));
 sky130_fd_sc_hd__clkbuf_1 _5004_ (.A(_1730_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _5005_ (.A0(net66),
    .A1(\mix1.data_o[43] ),
    .S(_1595_),
    .X(_1731_));
 sky130_fd_sc_hd__mux2_1 _5006_ (.A0(\sub1.data_o[43] ),
    .A1(_1731_),
    .S(_1597_),
    .X(_1732_));
 sky130_fd_sc_hd__a32o_1 _5007_ (.A1(\mix1.data_o[43] ),
    .A2(_1567_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[43] ),
    .X(_1733_));
 sky130_fd_sc_hd__a22o_1 _5008_ (.A1(_1607_),
    .A2(_1732_),
    .B1(_1733_),
    .B2(_1712_),
    .X(_1734_));
 sky130_fd_sc_hd__mux2_1 _5009_ (.A0(\ks1.key_reg[43] ),
    .A1(net195),
    .S(_1603_),
    .X(_1735_));
 sky130_fd_sc_hd__xor2_1 _5010_ (.A(_1734_),
    .B(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__mux2_1 _5011_ (.A0(net325),
    .A1(_1736_),
    .S(_1707_),
    .X(_1737_));
 sky130_fd_sc_hd__clkbuf_1 _5012_ (.A(_1737_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _5013_ (.A0(net67),
    .A1(\mix1.data_o[44] ),
    .S(_1595_),
    .X(_1738_));
 sky130_fd_sc_hd__mux2_1 _5014_ (.A0(\sub1.data_o[44] ),
    .A1(_1738_),
    .S(_1597_),
    .X(_1739_));
 sky130_fd_sc_hd__clkbuf_4 _5015_ (.A(_1306_),
    .X(_1740_));
 sky130_fd_sc_hd__a32o_1 _5016_ (.A1(\mix1.data_o[44] ),
    .A2(_1740_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[44] ),
    .X(_1741_));
 sky130_fd_sc_hd__a22o_1 _5017_ (.A1(_1607_),
    .A2(_1739_),
    .B1(_1741_),
    .B2(_1712_),
    .X(_1742_));
 sky130_fd_sc_hd__mux2_1 _5018_ (.A0(\ks1.key_reg[44] ),
    .A1(net196),
    .S(_1603_),
    .X(_1743_));
 sky130_fd_sc_hd__xor2_1 _5019_ (.A(_1742_),
    .B(_1743_),
    .X(_1744_));
 sky130_fd_sc_hd__mux2_1 _5020_ (.A0(net326),
    .A1(_1744_),
    .S(_1707_),
    .X(_1745_));
 sky130_fd_sc_hd__clkbuf_1 _5021_ (.A(_1745_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _5022_ (.A0(net68),
    .A1(\mix1.data_o[45] ),
    .S(_1595_),
    .X(_1746_));
 sky130_fd_sc_hd__mux2_1 _5023_ (.A0(\sub1.data_o[45] ),
    .A1(_1746_),
    .S(_1597_),
    .X(_1747_));
 sky130_fd_sc_hd__a32o_1 _5024_ (.A1(\mix1.data_o[45] ),
    .A2(_1740_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[45] ),
    .X(_1748_));
 sky130_fd_sc_hd__a22o_1 _5025_ (.A1(_1607_),
    .A2(_1747_),
    .B1(_1748_),
    .B2(_1712_),
    .X(_1749_));
 sky130_fd_sc_hd__mux2_1 _5026_ (.A0(\ks1.key_reg[45] ),
    .A1(net197),
    .S(_1603_),
    .X(_1750_));
 sky130_fd_sc_hd__xor2_1 _5027_ (.A(_1749_),
    .B(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__mux2_1 _5028_ (.A0(net327),
    .A1(_1751_),
    .S(_1707_),
    .X(_1752_));
 sky130_fd_sc_hd__clkbuf_1 _5029_ (.A(_1752_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _5030_ (.A0(net69),
    .A1(\mix1.data_o[46] ),
    .S(_1595_),
    .X(_1753_));
 sky130_fd_sc_hd__mux2_1 _5031_ (.A0(\sub1.data_o[46] ),
    .A1(_1753_),
    .S(_1597_),
    .X(_1754_));
 sky130_fd_sc_hd__a32o_1 _5032_ (.A1(\mix1.data_o[46] ),
    .A2(_1740_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[46] ),
    .X(_1755_));
 sky130_fd_sc_hd__a22o_1 _5033_ (.A1(_1607_),
    .A2(_1754_),
    .B1(_1755_),
    .B2(_1712_),
    .X(_1756_));
 sky130_fd_sc_hd__mux2_1 _5034_ (.A0(\ks1.key_reg[46] ),
    .A1(net198),
    .S(_1603_),
    .X(_1757_));
 sky130_fd_sc_hd__xor2_1 _5035_ (.A(_1756_),
    .B(_1757_),
    .X(_1758_));
 sky130_fd_sc_hd__mux2_1 _5036_ (.A0(net328),
    .A1(_1758_),
    .S(_1707_),
    .X(_1759_));
 sky130_fd_sc_hd__clkbuf_1 _5037_ (.A(_1759_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _5038_ (.A0(net70),
    .A1(\mix1.data_o[47] ),
    .S(_1595_),
    .X(_1760_));
 sky130_fd_sc_hd__mux2_1 _5039_ (.A0(\sub1.data_o[47] ),
    .A1(_1760_),
    .S(_1597_),
    .X(_1761_));
 sky130_fd_sc_hd__a32o_1 _5040_ (.A1(\mix1.data_o[47] ),
    .A2(_1740_),
    .A3(_1599_),
    .B1(_1600_),
    .B2(\sub1.data_o[47] ),
    .X(_1762_));
 sky130_fd_sc_hd__a22o_1 _5041_ (.A1(_1607_),
    .A2(_1761_),
    .B1(_1762_),
    .B2(_1712_),
    .X(_1763_));
 sky130_fd_sc_hd__mux2_1 _5042_ (.A0(\ks1.key_reg[47] ),
    .A1(net199),
    .S(_1603_),
    .X(_1764_));
 sky130_fd_sc_hd__xor2_1 _5043_ (.A(_1763_),
    .B(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__mux2_1 _5044_ (.A0(net329),
    .A1(_1765_),
    .S(_1707_),
    .X(_1766_));
 sky130_fd_sc_hd__clkbuf_1 _5045_ (.A(_1766_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _5046_ (.A0(net71),
    .A1(\mix1.data_o[48] ),
    .S(_1662_),
    .X(_1767_));
 sky130_fd_sc_hd__mux2_1 _5047_ (.A0(\sub1.data_o[48] ),
    .A1(_1767_),
    .S(_1664_),
    .X(_1768_));
 sky130_fd_sc_hd__a31o_1 _5048_ (.A1(_1217_),
    .A2(_1120_),
    .A3(\sub1.data_o[48] ),
    .B1(_1618_),
    .X(_1769_));
 sky130_fd_sc_hd__a21o_1 _5049_ (.A1(_1688_),
    .A2(_1768_),
    .B1(_1769_),
    .X(_1770_));
 sky130_fd_sc_hd__o21a_1 _5050_ (.A1(\mix1.data_o[48] ),
    .A2(_1329_),
    .B1(_1644_),
    .X(_1771_));
 sky130_fd_sc_hd__a221o_1 _5051_ (.A1(\sub1.data_o[48] ),
    .A2(_1617_),
    .B1(_1770_),
    .B2(_1771_),
    .C1(_1702_),
    .X(_1772_));
 sky130_fd_sc_hd__o21ai_2 _5052_ (.A1(_1639_),
    .A2(_1768_),
    .B1(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__mux2_1 _5053_ (.A0(\ks1.key_reg[48] ),
    .A1(net200),
    .S(_1648_),
    .X(_1774_));
 sky130_fd_sc_hd__xnor2_1 _5054_ (.A(_1773_),
    .B(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__mux2_1 _5055_ (.A0(net330),
    .A1(_1775_),
    .S(_1707_),
    .X(_1776_));
 sky130_fd_sc_hd__clkbuf_1 _5056_ (.A(_1776_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(net72),
    .A1(\mix1.data_o[49] ),
    .S(_1662_),
    .X(_1777_));
 sky130_fd_sc_hd__mux2_1 _5058_ (.A0(\sub1.data_o[49] ),
    .A1(_1777_),
    .S(_1664_),
    .X(_1778_));
 sky130_fd_sc_hd__clkbuf_4 _5059_ (.A(_1305_),
    .X(_1779_));
 sky130_fd_sc_hd__a31o_1 _5060_ (.A1(_1217_),
    .A2(\sub1.data_o[49] ),
    .A3(_1666_),
    .B1(_1779_),
    .X(_1780_));
 sky130_fd_sc_hd__a21o_1 _5061_ (.A1(_1688_),
    .A2(_1778_),
    .B1(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__clkbuf_4 _5062_ (.A(_1123_),
    .X(_1782_));
 sky130_fd_sc_hd__o21a_1 _5063_ (.A1(\mix1.data_o[49] ),
    .A2(_1782_),
    .B1(_1644_),
    .X(_1783_));
 sky130_fd_sc_hd__a221o_1 _5064_ (.A1(\sub1.data_o[49] ),
    .A2(_1617_),
    .B1(_1781_),
    .B2(_1783_),
    .C1(_1702_),
    .X(_1784_));
 sky130_fd_sc_hd__o21ai_2 _5065_ (.A1(_1639_),
    .A2(_1778_),
    .B1(_1784_),
    .Y(_1785_));
 sky130_fd_sc_hd__mux2_1 _5066_ (.A0(\ks1.key_reg[49] ),
    .A1(net201),
    .S(_1648_),
    .X(_1786_));
 sky130_fd_sc_hd__xnor2_1 _5067_ (.A(_1785_),
    .B(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__clkbuf_8 _5068_ (.A(_1510_),
    .X(_1788_));
 sky130_fd_sc_hd__mux2_1 _5069_ (.A0(net331),
    .A1(_1787_),
    .S(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__clkbuf_1 _5070_ (.A(_1789_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _5071_ (.A0(net74),
    .A1(\mix1.data_o[50] ),
    .S(_1662_),
    .X(_1790_));
 sky130_fd_sc_hd__mux2_1 _5072_ (.A0(\sub1.data_o[50] ),
    .A1(_1790_),
    .S(_1664_),
    .X(_1791_));
 sky130_fd_sc_hd__clkbuf_4 _5073_ (.A(_1348_),
    .X(_1792_));
 sky130_fd_sc_hd__clkbuf_4 _5074_ (.A(_1121_),
    .X(_1793_));
 sky130_fd_sc_hd__a31o_1 _5075_ (.A1(_1793_),
    .A2(\sub1.data_o[50] ),
    .A3(_1666_),
    .B1(_1779_),
    .X(_1794_));
 sky130_fd_sc_hd__a21o_1 _5076_ (.A1(_1688_),
    .A2(_1791_),
    .B1(_1794_),
    .X(_1795_));
 sky130_fd_sc_hd__o21a_1 _5077_ (.A1(\mix1.data_o[50] ),
    .A2(_1782_),
    .B1(_1644_),
    .X(_1796_));
 sky130_fd_sc_hd__a221o_1 _5078_ (.A1(\sub1.data_o[50] ),
    .A2(_1792_),
    .B1(_1795_),
    .B2(_1796_),
    .C1(_1702_),
    .X(_1797_));
 sky130_fd_sc_hd__o21ai_2 _5079_ (.A1(_1639_),
    .A2(_1791_),
    .B1(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__mux2_1 _5080_ (.A0(\ks1.key_reg[50] ),
    .A1(net203),
    .S(_1648_),
    .X(_1799_));
 sky130_fd_sc_hd__xnor2_1 _5081_ (.A(_1798_),
    .B(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__mux2_1 _5082_ (.A0(net333),
    .A1(_1800_),
    .S(_1788_),
    .X(_1801_));
 sky130_fd_sc_hd__clkbuf_1 _5083_ (.A(_1801_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _5084_ (.A0(net75),
    .A1(\mix1.data_o[51] ),
    .S(_1662_),
    .X(_1802_));
 sky130_fd_sc_hd__mux2_1 _5085_ (.A0(\sub1.data_o[51] ),
    .A1(_1802_),
    .S(_1664_),
    .X(_1803_));
 sky130_fd_sc_hd__a31o_1 _5086_ (.A1(_1793_),
    .A2(\sub1.data_o[51] ),
    .A3(_1666_),
    .B1(_1779_),
    .X(_1804_));
 sky130_fd_sc_hd__a21o_1 _5087_ (.A1(_1688_),
    .A2(_1803_),
    .B1(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__o21a_1 _5088_ (.A1(\mix1.data_o[51] ),
    .A2(_1782_),
    .B1(_1644_),
    .X(_1806_));
 sky130_fd_sc_hd__a221o_1 _5089_ (.A1(\sub1.data_o[51] ),
    .A2(_1792_),
    .B1(_1805_),
    .B2(_1806_),
    .C1(_1702_),
    .X(_1807_));
 sky130_fd_sc_hd__o21ai_2 _5090_ (.A1(_1639_),
    .A2(_1803_),
    .B1(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__mux2_1 _5091_ (.A0(\ks1.key_reg[51] ),
    .A1(net204),
    .S(_1648_),
    .X(_1809_));
 sky130_fd_sc_hd__xnor2_1 _5092_ (.A(_1808_),
    .B(_1809_),
    .Y(_1810_));
 sky130_fd_sc_hd__mux2_1 _5093_ (.A0(net334),
    .A1(_1810_),
    .S(_1788_),
    .X(_1811_));
 sky130_fd_sc_hd__clkbuf_1 _5094_ (.A(_1811_),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_8 _5095_ (.A(_0678_),
    .X(_1812_));
 sky130_fd_sc_hd__mux2_1 _5096_ (.A0(net76),
    .A1(\mix1.data_o[52] ),
    .S(_1662_),
    .X(_1813_));
 sky130_fd_sc_hd__mux2_1 _5097_ (.A0(\sub1.data_o[52] ),
    .A1(_1813_),
    .S(_1664_),
    .X(_1814_));
 sky130_fd_sc_hd__a31o_1 _5098_ (.A1(_1793_),
    .A2(\sub1.data_o[52] ),
    .A3(_1666_),
    .B1(_1779_),
    .X(_1815_));
 sky130_fd_sc_hd__a21o_1 _5099_ (.A1(_1688_),
    .A2(_1814_),
    .B1(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__buf_2 _5100_ (.A(_1519_),
    .X(_1817_));
 sky130_fd_sc_hd__o21a_1 _5101_ (.A1(\mix1.data_o[52] ),
    .A2(_1782_),
    .B1(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__a221o_1 _5102_ (.A1(\sub1.data_o[52] ),
    .A2(_1792_),
    .B1(_1816_),
    .B2(_1818_),
    .C1(_1702_),
    .X(_1819_));
 sky130_fd_sc_hd__o21ai_2 _5103_ (.A1(_1812_),
    .A2(_1814_),
    .B1(_1819_),
    .Y(_1820_));
 sky130_fd_sc_hd__clkbuf_8 _5104_ (.A(_1440_),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _5105_ (.A0(\ks1.key_reg[52] ),
    .A1(net205),
    .S(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__xnor2_1 _5106_ (.A(_1820_),
    .B(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hd__mux2_1 _5107_ (.A0(net335),
    .A1(_1823_),
    .S(_1788_),
    .X(_1824_));
 sky130_fd_sc_hd__clkbuf_1 _5108_ (.A(_1824_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _5109_ (.A0(net77),
    .A1(\mix1.data_o[53] ),
    .S(_1662_),
    .X(_1825_));
 sky130_fd_sc_hd__mux2_1 _5110_ (.A0(\sub1.data_o[53] ),
    .A1(_1825_),
    .S(_1664_),
    .X(_1826_));
 sky130_fd_sc_hd__a31o_1 _5111_ (.A1(\sub1.data_o[53] ),
    .A2(_1677_),
    .A3(_1666_),
    .B1(_1779_),
    .X(_1827_));
 sky130_fd_sc_hd__a21o_1 _5112_ (.A1(_1688_),
    .A2(_1826_),
    .B1(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__o21a_1 _5113_ (.A1(\mix1.data_o[53] ),
    .A2(_1782_),
    .B1(_1817_),
    .X(_1829_));
 sky130_fd_sc_hd__a221o_1 _5114_ (.A1(\sub1.data_o[53] ),
    .A2(_1792_),
    .B1(_1828_),
    .B2(_1829_),
    .C1(_1702_),
    .X(_1830_));
 sky130_fd_sc_hd__o21ai_2 _5115_ (.A1(_1812_),
    .A2(_1826_),
    .B1(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__mux2_1 _5116_ (.A0(\ks1.key_reg[53] ),
    .A1(net206),
    .S(_1821_),
    .X(_1832_));
 sky130_fd_sc_hd__xnor2_1 _5117_ (.A(_1831_),
    .B(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__mux2_1 _5118_ (.A0(net336),
    .A1(_1833_),
    .S(_1788_),
    .X(_1834_));
 sky130_fd_sc_hd__clkbuf_1 _5119_ (.A(_1834_),
    .X(_0069_));
 sky130_fd_sc_hd__buf_4 _5120_ (.A(_1337_),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_1 _5121_ (.A0(net78),
    .A1(\mix1.data_o[54] ),
    .S(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__clkbuf_4 _5122_ (.A(_1344_),
    .X(_1837_));
 sky130_fd_sc_hd__mux2_1 _5123_ (.A0(\sub1.data_o[54] ),
    .A1(_1836_),
    .S(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__a31o_1 _5124_ (.A1(\sub1.data_o[54] ),
    .A2(_1677_),
    .A3(_1666_),
    .B1(_1779_),
    .X(_1839_));
 sky130_fd_sc_hd__a21o_1 _5125_ (.A1(_1688_),
    .A2(_1838_),
    .B1(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__o21a_1 _5126_ (.A1(\mix1.data_o[54] ),
    .A2(_1782_),
    .B1(_1817_),
    .X(_1841_));
 sky130_fd_sc_hd__a221o_1 _5127_ (.A1(\sub1.data_o[54] ),
    .A2(_1792_),
    .B1(_1840_),
    .B2(_1841_),
    .C1(_1702_),
    .X(_1842_));
 sky130_fd_sc_hd__o21ai_2 _5128_ (.A1(_1812_),
    .A2(_1838_),
    .B1(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__mux2_1 _5129_ (.A0(\ks1.key_reg[54] ),
    .A1(net207),
    .S(_1821_),
    .X(_1844_));
 sky130_fd_sc_hd__xnor2_1 _5130_ (.A(_1843_),
    .B(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__mux2_1 _5131_ (.A0(net337),
    .A1(_1845_),
    .S(_1788_),
    .X(_1846_));
 sky130_fd_sc_hd__clkbuf_1 _5132_ (.A(_1846_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _5133_ (.A0(net79),
    .A1(\mix1.data_o[55] ),
    .S(_1835_),
    .X(_1847_));
 sky130_fd_sc_hd__mux2_1 _5134_ (.A0(\sub1.data_o[55] ),
    .A1(_1847_),
    .S(_1837_),
    .X(_1848_));
 sky130_fd_sc_hd__clkbuf_4 _5135_ (.A(_1119_),
    .X(_1849_));
 sky130_fd_sc_hd__a31o_1 _5136_ (.A1(_1793_),
    .A2(\sub1.data_o[55] ),
    .A3(_1849_),
    .B1(_1779_),
    .X(_1850_));
 sky130_fd_sc_hd__a21o_1 _5137_ (.A1(_1688_),
    .A2(_1848_),
    .B1(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__o21a_1 _5138_ (.A1(\mix1.data_o[55] ),
    .A2(_1782_),
    .B1(_1817_),
    .X(_1852_));
 sky130_fd_sc_hd__a221o_1 _5139_ (.A1(\sub1.data_o[55] ),
    .A2(_1792_),
    .B1(_1851_),
    .B2(_1852_),
    .C1(_1702_),
    .X(_1853_));
 sky130_fd_sc_hd__o21ai_2 _5140_ (.A1(_1812_),
    .A2(_1848_),
    .B1(_1853_),
    .Y(_1854_));
 sky130_fd_sc_hd__mux2_1 _5141_ (.A0(\ks1.key_reg[55] ),
    .A1(net208),
    .S(_1821_),
    .X(_1855_));
 sky130_fd_sc_hd__xnor2_1 _5142_ (.A(_1854_),
    .B(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__mux2_1 _5143_ (.A0(net338),
    .A1(_1856_),
    .S(_1788_),
    .X(_1857_));
 sky130_fd_sc_hd__clkbuf_1 _5144_ (.A(_1857_),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_4 _5145_ (.A(_1513_),
    .X(_1858_));
 sky130_fd_sc_hd__mux2_1 _5146_ (.A0(net80),
    .A1(\mix1.data_o[56] ),
    .S(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__clkbuf_4 _5147_ (.A(_1516_),
    .X(_1860_));
 sky130_fd_sc_hd__mux2_1 _5148_ (.A0(\sub1.data_o[56] ),
    .A1(_1859_),
    .S(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__buf_2 _5149_ (.A(_1519_),
    .X(_1862_));
 sky130_fd_sc_hd__buf_2 _5150_ (.A(_1354_),
    .X(_1863_));
 sky130_fd_sc_hd__a32o_1 _5151_ (.A1(\mix1.data_o[56] ),
    .A2(_1740_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[56] ),
    .X(_1864_));
 sky130_fd_sc_hd__a22o_1 _5152_ (.A1(_1607_),
    .A2(_1861_),
    .B1(_1864_),
    .B2(_1712_),
    .X(_1865_));
 sky130_fd_sc_hd__buf_4 _5153_ (.A(_1440_),
    .X(_1866_));
 sky130_fd_sc_hd__mux2_1 _5154_ (.A0(\ks1.key_reg[56] ),
    .A1(net209),
    .S(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__xor2_1 _5155_ (.A(_1865_),
    .B(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__mux2_1 _5156_ (.A0(net339),
    .A1(_1868_),
    .S(_1788_),
    .X(_1869_));
 sky130_fd_sc_hd__clkbuf_1 _5157_ (.A(_1869_),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_4 _5158_ (.A(_1349_),
    .X(_1870_));
 sky130_fd_sc_hd__mux2_1 _5159_ (.A0(net81),
    .A1(\mix1.data_o[57] ),
    .S(_1858_),
    .X(_1871_));
 sky130_fd_sc_hd__mux2_1 _5160_ (.A0(\sub1.data_o[57] ),
    .A1(_1871_),
    .S(_1860_),
    .X(_1872_));
 sky130_fd_sc_hd__a32o_1 _5161_ (.A1(\mix1.data_o[57] ),
    .A2(_1740_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[57] ),
    .X(_1873_));
 sky130_fd_sc_hd__a22o_1 _5162_ (.A1(_1870_),
    .A2(_1872_),
    .B1(_1873_),
    .B2(_1712_),
    .X(_1874_));
 sky130_fd_sc_hd__mux2_1 _5163_ (.A0(\ks1.key_reg[57] ),
    .A1(net210),
    .S(_1866_),
    .X(_1875_));
 sky130_fd_sc_hd__xor2_1 _5164_ (.A(_1874_),
    .B(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__mux2_1 _5165_ (.A0(net340),
    .A1(_1876_),
    .S(_1788_),
    .X(_1877_));
 sky130_fd_sc_hd__clkbuf_1 _5166_ (.A(_1877_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _5167_ (.A0(net82),
    .A1(\mix1.data_o[58] ),
    .S(_1858_),
    .X(_1878_));
 sky130_fd_sc_hd__mux2_1 _5168_ (.A0(\sub1.data_o[58] ),
    .A1(_1878_),
    .S(_1860_),
    .X(_1879_));
 sky130_fd_sc_hd__a32o_1 _5169_ (.A1(\mix1.data_o[58] ),
    .A2(_1740_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[58] ),
    .X(_1880_));
 sky130_fd_sc_hd__clkbuf_4 _5170_ (.A(_0677_),
    .X(_1881_));
 sky130_fd_sc_hd__a22o_1 _5171_ (.A1(_1870_),
    .A2(_1879_),
    .B1(_1880_),
    .B2(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _5172_ (.A0(\ks1.key_reg[58] ),
    .A1(net211),
    .S(_1866_),
    .X(_1883_));
 sky130_fd_sc_hd__xor2_1 _5173_ (.A(_1882_),
    .B(_1883_),
    .X(_1884_));
 sky130_fd_sc_hd__mux2_1 _5174_ (.A0(net341),
    .A1(_1884_),
    .S(_1788_),
    .X(_1885_));
 sky130_fd_sc_hd__clkbuf_1 _5175_ (.A(_1885_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _5176_ (.A0(net83),
    .A1(\mix1.data_o[59] ),
    .S(_1858_),
    .X(_1886_));
 sky130_fd_sc_hd__mux2_1 _5177_ (.A0(\sub1.data_o[59] ),
    .A1(_1886_),
    .S(_1860_),
    .X(_1887_));
 sky130_fd_sc_hd__a32o_1 _5178_ (.A1(\mix1.data_o[59] ),
    .A2(_1740_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[59] ),
    .X(_1888_));
 sky130_fd_sc_hd__a22o_1 _5179_ (.A1(_1870_),
    .A2(_1887_),
    .B1(_1888_),
    .B2(_1881_),
    .X(_1889_));
 sky130_fd_sc_hd__mux2_1 _5180_ (.A0(\ks1.key_reg[59] ),
    .A1(net212),
    .S(_1866_),
    .X(_1890_));
 sky130_fd_sc_hd__xor2_1 _5181_ (.A(_1889_),
    .B(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__buf_4 _5182_ (.A(_1510_),
    .X(_1892_));
 sky130_fd_sc_hd__mux2_1 _5183_ (.A0(net342),
    .A1(_1891_),
    .S(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__clkbuf_1 _5184_ (.A(_1893_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _5185_ (.A0(net85),
    .A1(\mix1.data_o[60] ),
    .S(_1858_),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_1 _5186_ (.A0(\sub1.data_o[60] ),
    .A1(_1894_),
    .S(_1860_),
    .X(_1895_));
 sky130_fd_sc_hd__a32o_1 _5187_ (.A1(\mix1.data_o[60] ),
    .A2(_1740_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[60] ),
    .X(_1896_));
 sky130_fd_sc_hd__a22o_1 _5188_ (.A1(_1870_),
    .A2(_1895_),
    .B1(_1896_),
    .B2(_1881_),
    .X(_1897_));
 sky130_fd_sc_hd__mux2_1 _5189_ (.A0(\ks1.key_reg[60] ),
    .A1(net214),
    .S(_1866_),
    .X(_1898_));
 sky130_fd_sc_hd__xor2_1 _5190_ (.A(_1897_),
    .B(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__mux2_1 _5191_ (.A0(net344),
    .A1(_1899_),
    .S(_1892_),
    .X(_1900_));
 sky130_fd_sc_hd__clkbuf_1 _5192_ (.A(_1900_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _5193_ (.A0(net86),
    .A1(\mix1.data_o[61] ),
    .S(_1858_),
    .X(_1901_));
 sky130_fd_sc_hd__mux2_1 _5194_ (.A0(\sub1.data_o[61] ),
    .A1(_1901_),
    .S(_1860_),
    .X(_1902_));
 sky130_fd_sc_hd__a32o_1 _5195_ (.A1(\mix1.data_o[61] ),
    .A2(_1740_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[61] ),
    .X(_1903_));
 sky130_fd_sc_hd__a22o_1 _5196_ (.A1(_1870_),
    .A2(_1902_),
    .B1(_1903_),
    .B2(_1881_),
    .X(_1904_));
 sky130_fd_sc_hd__mux2_1 _5197_ (.A0(\ks1.key_reg[61] ),
    .A1(net215),
    .S(_1866_),
    .X(_1905_));
 sky130_fd_sc_hd__xor2_1 _5198_ (.A(_1904_),
    .B(_1905_),
    .X(_1906_));
 sky130_fd_sc_hd__mux2_1 _5199_ (.A0(net345),
    .A1(_1906_),
    .S(_1892_),
    .X(_1907_));
 sky130_fd_sc_hd__clkbuf_1 _5200_ (.A(_1907_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _5201_ (.A0(net87),
    .A1(\mix1.data_o[62] ),
    .S(_1858_),
    .X(_1908_));
 sky130_fd_sc_hd__mux2_1 _5202_ (.A0(\sub1.data_o[62] ),
    .A1(_1908_),
    .S(_1860_),
    .X(_1909_));
 sky130_fd_sc_hd__clkbuf_4 _5203_ (.A(_1306_),
    .X(_1910_));
 sky130_fd_sc_hd__a32o_1 _5204_ (.A1(\mix1.data_o[62] ),
    .A2(_1910_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[62] ),
    .X(_1911_));
 sky130_fd_sc_hd__a22o_1 _5205_ (.A1(_1870_),
    .A2(_1909_),
    .B1(_1911_),
    .B2(_1881_),
    .X(_1912_));
 sky130_fd_sc_hd__mux2_1 _5206_ (.A0(\ks1.key_reg[62] ),
    .A1(net216),
    .S(_1866_),
    .X(_1913_));
 sky130_fd_sc_hd__xor2_1 _5207_ (.A(_1912_),
    .B(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__mux2_1 _5208_ (.A0(net346),
    .A1(_1914_),
    .S(_1892_),
    .X(_1915_));
 sky130_fd_sc_hd__clkbuf_1 _5209_ (.A(_1915_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _5210_ (.A0(net88),
    .A1(\mix1.data_o[63] ),
    .S(_1858_),
    .X(_1916_));
 sky130_fd_sc_hd__mux2_1 _5211_ (.A0(\sub1.data_o[63] ),
    .A1(_1916_),
    .S(_1860_),
    .X(_1917_));
 sky130_fd_sc_hd__a32o_1 _5212_ (.A1(\mix1.data_o[63] ),
    .A2(_1910_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[63] ),
    .X(_1918_));
 sky130_fd_sc_hd__a22o_1 _5213_ (.A1(_1870_),
    .A2(_1917_),
    .B1(_1918_),
    .B2(_1881_),
    .X(_1919_));
 sky130_fd_sc_hd__mux2_1 _5214_ (.A0(\ks1.key_reg[63] ),
    .A1(net217),
    .S(_1866_),
    .X(_1920_));
 sky130_fd_sc_hd__xor2_1 _5215_ (.A(_1919_),
    .B(_1920_),
    .X(_1921_));
 sky130_fd_sc_hd__mux2_1 _5216_ (.A0(net347),
    .A1(_1921_),
    .S(_1892_),
    .X(_1922_));
 sky130_fd_sc_hd__clkbuf_1 _5217_ (.A(_1922_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _5218_ (.A0(net89),
    .A1(\mix1.data_o[64] ),
    .S(_1858_),
    .X(_1923_));
 sky130_fd_sc_hd__mux2_1 _5219_ (.A0(\sub1.data_o[64] ),
    .A1(_1923_),
    .S(_1860_),
    .X(_1924_));
 sky130_fd_sc_hd__a32o_1 _5220_ (.A1(\mix1.data_o[64] ),
    .A2(_1910_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[64] ),
    .X(_1925_));
 sky130_fd_sc_hd__a22o_1 _5221_ (.A1(_1870_),
    .A2(_1924_),
    .B1(_1925_),
    .B2(_1881_),
    .X(_1926_));
 sky130_fd_sc_hd__mux2_1 _5222_ (.A0(\ks1.key_reg[64] ),
    .A1(net218),
    .S(_1866_),
    .X(_1927_));
 sky130_fd_sc_hd__xor2_1 _5223_ (.A(_1926_),
    .B(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__mux2_1 _5224_ (.A0(net348),
    .A1(_1928_),
    .S(_1892_),
    .X(_1929_));
 sky130_fd_sc_hd__clkbuf_1 _5225_ (.A(_1929_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _5226_ (.A0(net90),
    .A1(\mix1.data_o[65] ),
    .S(_1858_),
    .X(_1930_));
 sky130_fd_sc_hd__mux2_1 _5227_ (.A0(\sub1.data_o[65] ),
    .A1(_1930_),
    .S(_1860_),
    .X(_1931_));
 sky130_fd_sc_hd__a32o_1 _5228_ (.A1(\mix1.data_o[65] ),
    .A2(_1910_),
    .A3(_1862_),
    .B1(_1863_),
    .B2(\sub1.data_o[65] ),
    .X(_1932_));
 sky130_fd_sc_hd__a22o_1 _5229_ (.A1(_1870_),
    .A2(_1931_),
    .B1(_1932_),
    .B2(_1881_),
    .X(_1933_));
 sky130_fd_sc_hd__mux2_1 _5230_ (.A0(\ks1.key_reg[65] ),
    .A1(net219),
    .S(_1866_),
    .X(_1934_));
 sky130_fd_sc_hd__xor2_1 _5231_ (.A(_1933_),
    .B(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__mux2_1 _5232_ (.A0(net349),
    .A1(_1935_),
    .S(_1892_),
    .X(_1936_));
 sky130_fd_sc_hd__clkbuf_1 _5233_ (.A(_1936_),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_4 _5234_ (.A(_1513_),
    .X(_1937_));
 sky130_fd_sc_hd__mux2_1 _5235_ (.A0(net91),
    .A1(\mix1.data_o[66] ),
    .S(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__clkbuf_4 _5236_ (.A(_1516_),
    .X(_1939_));
 sky130_fd_sc_hd__mux2_1 _5237_ (.A0(\sub1.data_o[66] ),
    .A1(_1938_),
    .S(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__buf_2 _5238_ (.A(_1519_),
    .X(_1941_));
 sky130_fd_sc_hd__clkbuf_4 _5239_ (.A(_1354_),
    .X(_1942_));
 sky130_fd_sc_hd__a32o_1 _5240_ (.A1(\mix1.data_o[66] ),
    .A2(_1910_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[66] ),
    .X(_1943_));
 sky130_fd_sc_hd__a22o_1 _5241_ (.A1(_1870_),
    .A2(_1940_),
    .B1(_1943_),
    .B2(_1881_),
    .X(_1944_));
 sky130_fd_sc_hd__buf_4 _5242_ (.A(_1440_),
    .X(_1945_));
 sky130_fd_sc_hd__mux2_2 _5243_ (.A0(\ks1.key_reg[66] ),
    .A1(net220),
    .S(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__xor2_1 _5244_ (.A(_1944_),
    .B(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__mux2_1 _5245_ (.A0(net350),
    .A1(_1947_),
    .S(_1892_),
    .X(_1948_));
 sky130_fd_sc_hd__clkbuf_1 _5246_ (.A(_1948_),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_4 _5247_ (.A(_1349_),
    .X(_1949_));
 sky130_fd_sc_hd__mux2_1 _5248_ (.A0(net92),
    .A1(\mix1.data_o[67] ),
    .S(_1937_),
    .X(_1950_));
 sky130_fd_sc_hd__mux2_1 _5249_ (.A0(\sub1.data_o[67] ),
    .A1(_1950_),
    .S(_1939_),
    .X(_1951_));
 sky130_fd_sc_hd__a32o_1 _5250_ (.A1(\mix1.data_o[67] ),
    .A2(_1910_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[67] ),
    .X(_1952_));
 sky130_fd_sc_hd__a22o_1 _5251_ (.A1(_1949_),
    .A2(_1951_),
    .B1(_1952_),
    .B2(_1881_),
    .X(_1953_));
 sky130_fd_sc_hd__mux2_2 _5252_ (.A0(\ks1.key_reg[67] ),
    .A1(net221),
    .S(_1945_),
    .X(_1954_));
 sky130_fd_sc_hd__xor2_1 _5253_ (.A(_1953_),
    .B(_1954_),
    .X(_1955_));
 sky130_fd_sc_hd__mux2_1 _5254_ (.A0(net351),
    .A1(_1955_),
    .S(_1892_),
    .X(_1956_));
 sky130_fd_sc_hd__clkbuf_1 _5255_ (.A(_1956_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(net93),
    .A1(\mix1.data_o[68] ),
    .S(_1937_),
    .X(_1957_));
 sky130_fd_sc_hd__mux2_1 _5257_ (.A0(\sub1.data_o[68] ),
    .A1(_1957_),
    .S(_1939_),
    .X(_1958_));
 sky130_fd_sc_hd__a32o_1 _5258_ (.A1(\mix1.data_o[68] ),
    .A2(_1910_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[68] ),
    .X(_1959_));
 sky130_fd_sc_hd__clkbuf_4 _5259_ (.A(_0677_),
    .X(_1960_));
 sky130_fd_sc_hd__a22o_2 _5260_ (.A1(_1949_),
    .A2(_1958_),
    .B1(_1959_),
    .B2(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__mux2_1 _5261_ (.A0(\ks1.key_reg[68] ),
    .A1(net222),
    .S(_1945_),
    .X(_1962_));
 sky130_fd_sc_hd__xor2_1 _5262_ (.A(_1961_),
    .B(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__mux2_1 _5263_ (.A0(net352),
    .A1(_1963_),
    .S(_1892_),
    .X(_1964_));
 sky130_fd_sc_hd__clkbuf_1 _5264_ (.A(_1964_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _5265_ (.A0(net94),
    .A1(\mix1.data_o[69] ),
    .S(_1937_),
    .X(_1965_));
 sky130_fd_sc_hd__mux2_1 _5266_ (.A0(\sub1.data_o[69] ),
    .A1(_1965_),
    .S(_1939_),
    .X(_1966_));
 sky130_fd_sc_hd__a32o_1 _5267_ (.A1(\mix1.data_o[69] ),
    .A2(_1910_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[69] ),
    .X(_1967_));
 sky130_fd_sc_hd__a22o_1 _5268_ (.A1(_1949_),
    .A2(_1966_),
    .B1(_1967_),
    .B2(_1960_),
    .X(_1968_));
 sky130_fd_sc_hd__mux2_1 _5269_ (.A0(\ks1.key_reg[69] ),
    .A1(net223),
    .S(_1945_),
    .X(_1969_));
 sky130_fd_sc_hd__xor2_1 _5270_ (.A(_1968_),
    .B(_1969_),
    .X(_1970_));
 sky130_fd_sc_hd__clkbuf_8 _5271_ (.A(_1510_),
    .X(_1971_));
 sky130_fd_sc_hd__mux2_1 _5272_ (.A0(net353),
    .A1(_1970_),
    .S(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__clkbuf_1 _5273_ (.A(_1972_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _5274_ (.A0(net96),
    .A1(\mix1.data_o[70] ),
    .S(_1937_),
    .X(_1973_));
 sky130_fd_sc_hd__mux2_1 _5275_ (.A0(\sub1.data_o[70] ),
    .A1(_1973_),
    .S(_1939_),
    .X(_1974_));
 sky130_fd_sc_hd__a32o_1 _5276_ (.A1(\mix1.data_o[70] ),
    .A2(_1910_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[70] ),
    .X(_1975_));
 sky130_fd_sc_hd__a22o_1 _5277_ (.A1(_1949_),
    .A2(_1974_),
    .B1(_1975_),
    .B2(_1960_),
    .X(_1976_));
 sky130_fd_sc_hd__mux2_1 _5278_ (.A0(\ks1.key_reg[70] ),
    .A1(net225),
    .S(_1945_),
    .X(_1977_));
 sky130_fd_sc_hd__xor2_1 _5279_ (.A(_1976_),
    .B(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__mux2_1 _5280_ (.A0(net355),
    .A1(_1978_),
    .S(_1971_),
    .X(_1979_));
 sky130_fd_sc_hd__clkbuf_1 _5281_ (.A(_1979_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _5282_ (.A0(net97),
    .A1(\mix1.data_o[71] ),
    .S(_1937_),
    .X(_1980_));
 sky130_fd_sc_hd__mux2_1 _5283_ (.A0(\sub1.data_o[71] ),
    .A1(_1980_),
    .S(_1939_),
    .X(_1981_));
 sky130_fd_sc_hd__a32o_1 _5284_ (.A1(\mix1.data_o[71] ),
    .A2(_1910_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[71] ),
    .X(_1982_));
 sky130_fd_sc_hd__a22o_1 _5285_ (.A1(_1949_),
    .A2(_1981_),
    .B1(_1982_),
    .B2(_1960_),
    .X(_1983_));
 sky130_fd_sc_hd__mux2_1 _5286_ (.A0(\ks1.key_reg[71] ),
    .A1(net226),
    .S(_1945_),
    .X(_1984_));
 sky130_fd_sc_hd__xor2_1 _5287_ (.A(_1983_),
    .B(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__mux2_1 _5288_ (.A0(net356),
    .A1(_1985_),
    .S(_1971_),
    .X(_1986_));
 sky130_fd_sc_hd__clkbuf_1 _5289_ (.A(_1986_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _5290_ (.A0(net98),
    .A1(\mix1.data_o[72] ),
    .S(_1937_),
    .X(_1987_));
 sky130_fd_sc_hd__mux2_1 _5291_ (.A0(\sub1.data_o[72] ),
    .A1(_1987_),
    .S(_1939_),
    .X(_1988_));
 sky130_fd_sc_hd__clkbuf_4 _5292_ (.A(_1306_),
    .X(_1989_));
 sky130_fd_sc_hd__a32o_1 _5293_ (.A1(\mix1.data_o[72] ),
    .A2(_1989_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[72] ),
    .X(_1990_));
 sky130_fd_sc_hd__a22o_1 _5294_ (.A1(_1949_),
    .A2(_1988_),
    .B1(_1990_),
    .B2(_1960_),
    .X(_1991_));
 sky130_fd_sc_hd__mux2_1 _5295_ (.A0(\ks1.key_reg[72] ),
    .A1(net227),
    .S(_1945_),
    .X(_1992_));
 sky130_fd_sc_hd__xor2_1 _5296_ (.A(_1991_),
    .B(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__mux2_1 _5297_ (.A0(net357),
    .A1(_1993_),
    .S(_1971_),
    .X(_1994_));
 sky130_fd_sc_hd__clkbuf_1 _5298_ (.A(_1994_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _5299_ (.A0(net99),
    .A1(\mix1.data_o[73] ),
    .S(_1937_),
    .X(_1995_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(\sub1.data_o[73] ),
    .A1(_1995_),
    .S(_1939_),
    .X(_1996_));
 sky130_fd_sc_hd__a32o_1 _5301_ (.A1(\mix1.data_o[73] ),
    .A2(_1989_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[73] ),
    .X(_1997_));
 sky130_fd_sc_hd__a22o_1 _5302_ (.A1(_1949_),
    .A2(_1996_),
    .B1(_1997_),
    .B2(_1960_),
    .X(_1998_));
 sky130_fd_sc_hd__mux2_1 _5303_ (.A0(\ks1.key_reg[73] ),
    .A1(net228),
    .S(_1945_),
    .X(_1999_));
 sky130_fd_sc_hd__xor2_1 _5304_ (.A(_1998_),
    .B(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__mux2_1 _5305_ (.A0(net358),
    .A1(_2000_),
    .S(_1971_),
    .X(_2001_));
 sky130_fd_sc_hd__clkbuf_1 _5306_ (.A(_2001_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _5307_ (.A0(net100),
    .A1(\mix1.data_o[74] ),
    .S(_1937_),
    .X(_2002_));
 sky130_fd_sc_hd__mux2_1 _5308_ (.A0(\sub1.data_o[74] ),
    .A1(_2002_),
    .S(_1939_),
    .X(_2003_));
 sky130_fd_sc_hd__a32o_1 _5309_ (.A1(\mix1.data_o[74] ),
    .A2(_1989_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[74] ),
    .X(_2004_));
 sky130_fd_sc_hd__a22o_1 _5310_ (.A1(_1949_),
    .A2(_2003_),
    .B1(_2004_),
    .B2(_1960_),
    .X(_2005_));
 sky130_fd_sc_hd__mux2_1 _5311_ (.A0(\ks1.key_reg[74] ),
    .A1(net229),
    .S(_1945_),
    .X(_2006_));
 sky130_fd_sc_hd__xor2_1 _5312_ (.A(_2005_),
    .B(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__mux2_1 _5313_ (.A0(net359),
    .A1(_2007_),
    .S(_1971_),
    .X(_2008_));
 sky130_fd_sc_hd__clkbuf_1 _5314_ (.A(_2008_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _5315_ (.A0(net101),
    .A1(\mix1.data_o[75] ),
    .S(_1937_),
    .X(_2009_));
 sky130_fd_sc_hd__mux2_1 _5316_ (.A0(\sub1.data_o[75] ),
    .A1(_2009_),
    .S(_1939_),
    .X(_2010_));
 sky130_fd_sc_hd__a32o_1 _5317_ (.A1(\mix1.data_o[75] ),
    .A2(_1989_),
    .A3(_1941_),
    .B1(_1942_),
    .B2(\sub1.data_o[75] ),
    .X(_2011_));
 sky130_fd_sc_hd__a22o_1 _5318_ (.A1(_1949_),
    .A2(_2010_),
    .B1(_2011_),
    .B2(_1960_),
    .X(_2012_));
 sky130_fd_sc_hd__mux2_1 _5319_ (.A0(\ks1.key_reg[75] ),
    .A1(net230),
    .S(_1945_),
    .X(_2013_));
 sky130_fd_sc_hd__xor2_1 _5320_ (.A(_2012_),
    .B(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__mux2_1 _5321_ (.A0(net360),
    .A1(_2014_),
    .S(_1971_),
    .X(_2015_));
 sky130_fd_sc_hd__clkbuf_1 _5322_ (.A(_2015_),
    .X(_0091_));
 sky130_fd_sc_hd__buf_4 _5323_ (.A(_1513_),
    .X(_2016_));
 sky130_fd_sc_hd__mux2_1 _5324_ (.A0(net102),
    .A1(\mix1.data_o[76] ),
    .S(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__buf_4 _5325_ (.A(_1516_),
    .X(_2018_));
 sky130_fd_sc_hd__mux2_1 _5326_ (.A0(\sub1.data_o[76] ),
    .A1(_2017_),
    .S(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__clkbuf_4 _5327_ (.A(_1519_),
    .X(_2020_));
 sky130_fd_sc_hd__clkbuf_4 _5328_ (.A(_1354_),
    .X(_2021_));
 sky130_fd_sc_hd__a32o_1 _5329_ (.A1(\mix1.data_o[76] ),
    .A2(_1989_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[76] ),
    .X(_2022_));
 sky130_fd_sc_hd__a22o_1 _5330_ (.A1(_1949_),
    .A2(_2019_),
    .B1(_2022_),
    .B2(_1960_),
    .X(_2023_));
 sky130_fd_sc_hd__buf_4 _5331_ (.A(_1440_),
    .X(_2024_));
 sky130_fd_sc_hd__mux2_1 _5332_ (.A0(\ks1.key_reg[76] ),
    .A1(net231),
    .S(_2024_),
    .X(_2025_));
 sky130_fd_sc_hd__xor2_1 _5333_ (.A(_2023_),
    .B(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__mux2_1 _5334_ (.A0(net361),
    .A1(_2026_),
    .S(_1971_),
    .X(_2027_));
 sky130_fd_sc_hd__clkbuf_1 _5335_ (.A(_2027_),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_4 _5336_ (.A(_1349_),
    .X(_2028_));
 sky130_fd_sc_hd__mux2_1 _5337_ (.A0(net103),
    .A1(\mix1.data_o[77] ),
    .S(_2016_),
    .X(_2029_));
 sky130_fd_sc_hd__mux2_1 _5338_ (.A0(\sub1.data_o[77] ),
    .A1(_2029_),
    .S(_2018_),
    .X(_2030_));
 sky130_fd_sc_hd__a32o_1 _5339_ (.A1(\mix1.data_o[77] ),
    .A2(_1989_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[77] ),
    .X(_2031_));
 sky130_fd_sc_hd__a22o_1 _5340_ (.A1(_2028_),
    .A2(_2030_),
    .B1(_2031_),
    .B2(_1960_),
    .X(_2032_));
 sky130_fd_sc_hd__mux2_1 _5341_ (.A0(\ks1.key_reg[77] ),
    .A1(net232),
    .S(_2024_),
    .X(_2033_));
 sky130_fd_sc_hd__xor2_1 _5342_ (.A(_2032_),
    .B(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__mux2_1 _5343_ (.A0(net362),
    .A1(_2034_),
    .S(_1971_),
    .X(_2035_));
 sky130_fd_sc_hd__clkbuf_1 _5344_ (.A(_2035_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _5345_ (.A0(net104),
    .A1(\mix1.data_o[78] ),
    .S(_2016_),
    .X(_2036_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(\sub1.data_o[78] ),
    .A1(_2036_),
    .S(_2018_),
    .X(_2037_));
 sky130_fd_sc_hd__a32o_1 _5347_ (.A1(\mix1.data_o[78] ),
    .A2(_1989_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[78] ),
    .X(_2038_));
 sky130_fd_sc_hd__clkbuf_4 _5348_ (.A(_0677_),
    .X(_2039_));
 sky130_fd_sc_hd__a22o_1 _5349_ (.A1(_2028_),
    .A2(_2037_),
    .B1(_2038_),
    .B2(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(\ks1.key_reg[78] ),
    .A1(net233),
    .S(_2024_),
    .X(_2041_));
 sky130_fd_sc_hd__xor2_1 _5351_ (.A(_2040_),
    .B(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__mux2_1 _5352_ (.A0(net363),
    .A1(_2042_),
    .S(_1971_),
    .X(_2043_));
 sky130_fd_sc_hd__clkbuf_1 _5353_ (.A(_2043_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _5354_ (.A0(net105),
    .A1(\mix1.data_o[79] ),
    .S(_2016_),
    .X(_2044_));
 sky130_fd_sc_hd__mux2_1 _5355_ (.A0(\sub1.data_o[79] ),
    .A1(_2044_),
    .S(_2018_),
    .X(_2045_));
 sky130_fd_sc_hd__a32o_1 _5356_ (.A1(\mix1.data_o[79] ),
    .A2(_1989_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[79] ),
    .X(_2046_));
 sky130_fd_sc_hd__a22o_1 _5357_ (.A1(_2028_),
    .A2(_2045_),
    .B1(_2046_),
    .B2(_2039_),
    .X(_2047_));
 sky130_fd_sc_hd__mux2_1 _5358_ (.A0(\ks1.key_reg[79] ),
    .A1(net234),
    .S(_2024_),
    .X(_2048_));
 sky130_fd_sc_hd__xor2_1 _5359_ (.A(_2047_),
    .B(_2048_),
    .X(_2049_));
 sky130_fd_sc_hd__clkbuf_8 _5360_ (.A(_1510_),
    .X(_2050_));
 sky130_fd_sc_hd__mux2_1 _5361_ (.A0(net364),
    .A1(_2049_),
    .S(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__clkbuf_1 _5362_ (.A(_2051_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _5363_ (.A0(net107),
    .A1(\mix1.data_o[80] ),
    .S(_1835_),
    .X(_2052_));
 sky130_fd_sc_hd__mux2_1 _5364_ (.A0(\sub1.data_o[80] ),
    .A1(_2052_),
    .S(_1837_),
    .X(_2053_));
 sky130_fd_sc_hd__clkbuf_4 _5365_ (.A(_1122_),
    .X(_2054_));
 sky130_fd_sc_hd__a31o_1 _5366_ (.A1(_1793_),
    .A2(_1120_),
    .A3(\sub1.data_o[80] ),
    .B1(_1779_),
    .X(_2055_));
 sky130_fd_sc_hd__a21o_1 _5367_ (.A1(_2054_),
    .A2(_2053_),
    .B1(_2055_),
    .X(_2056_));
 sky130_fd_sc_hd__o21a_1 _5368_ (.A1(\mix1.data_o[80] ),
    .A2(_1782_),
    .B1(_1817_),
    .X(_2057_));
 sky130_fd_sc_hd__a221o_1 _5369_ (.A1(\sub1.data_o[80] ),
    .A2(_1792_),
    .B1(_2056_),
    .B2(_2057_),
    .C1(_1702_),
    .X(_2058_));
 sky130_fd_sc_hd__o21ai_1 _5370_ (.A1(_1812_),
    .A2(_2053_),
    .B1(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(\ks1.key_reg[80] ),
    .A1(net236),
    .S(_1821_),
    .X(_2060_));
 sky130_fd_sc_hd__xnor2_1 _5372_ (.A(_2059_),
    .B(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(net366),
    .A1(_2061_),
    .S(_2050_),
    .X(_2062_));
 sky130_fd_sc_hd__clkbuf_1 _5374_ (.A(_2062_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _5375_ (.A0(net108),
    .A1(\mix1.data_o[81] ),
    .S(_1835_),
    .X(_2063_));
 sky130_fd_sc_hd__mux2_1 _5376_ (.A0(\sub1.data_o[81] ),
    .A1(_2063_),
    .S(_1837_),
    .X(_2064_));
 sky130_fd_sc_hd__a31o_1 _5377_ (.A1(_1793_),
    .A2(\sub1.data_o[81] ),
    .A3(_1849_),
    .B1(_1779_),
    .X(_2065_));
 sky130_fd_sc_hd__a21o_1 _5378_ (.A1(_2054_),
    .A2(_2064_),
    .B1(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__o21a_1 _5379_ (.A1(\mix1.data_o[81] ),
    .A2(_1782_),
    .B1(_1817_),
    .X(_2067_));
 sky130_fd_sc_hd__clkbuf_4 _5380_ (.A(_1114_),
    .X(_2068_));
 sky130_fd_sc_hd__a221o_1 _5381_ (.A1(\sub1.data_o[81] ),
    .A2(_1792_),
    .B1(_2066_),
    .B2(_2067_),
    .C1(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__o21ai_2 _5382_ (.A1(_1812_),
    .A2(_2064_),
    .B1(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(\ks1.key_reg[81] ),
    .A1(net237),
    .S(_1821_),
    .X(_2071_));
 sky130_fd_sc_hd__xnor2_1 _5384_ (.A(_2070_),
    .B(_2071_),
    .Y(_2072_));
 sky130_fd_sc_hd__mux2_1 _5385_ (.A0(net367),
    .A1(_2072_),
    .S(_2050_),
    .X(_2073_));
 sky130_fd_sc_hd__clkbuf_1 _5386_ (.A(_2073_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _5387_ (.A0(net109),
    .A1(\mix1.data_o[82] ),
    .S(_1835_),
    .X(_2074_));
 sky130_fd_sc_hd__mux2_1 _5388_ (.A0(\sub1.data_o[82] ),
    .A1(_2074_),
    .S(_1837_),
    .X(_2075_));
 sky130_fd_sc_hd__a31o_1 _5389_ (.A1(_1793_),
    .A2(\sub1.data_o[82] ),
    .A3(_1849_),
    .B1(_1779_),
    .X(_2076_));
 sky130_fd_sc_hd__a21o_1 _5390_ (.A1(_2054_),
    .A2(_2075_),
    .B1(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__o21a_1 _5391_ (.A1(\mix1.data_o[82] ),
    .A2(_1782_),
    .B1(_1817_),
    .X(_2078_));
 sky130_fd_sc_hd__a221o_1 _5392_ (.A1(\sub1.data_o[82] ),
    .A2(_1792_),
    .B1(_2077_),
    .B2(_2078_),
    .C1(_2068_),
    .X(_2079_));
 sky130_fd_sc_hd__o21ai_2 _5393_ (.A1(_1812_),
    .A2(_2075_),
    .B1(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__mux2_1 _5394_ (.A0(\ks1.key_reg[82] ),
    .A1(net238),
    .S(_1821_),
    .X(_2081_));
 sky130_fd_sc_hd__xnor2_1 _5395_ (.A(_2080_),
    .B(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__mux2_1 _5396_ (.A0(net368),
    .A1(_2082_),
    .S(_2050_),
    .X(_2083_));
 sky130_fd_sc_hd__clkbuf_1 _5397_ (.A(_2083_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _5398_ (.A0(net110),
    .A1(\mix1.data_o[83] ),
    .S(_1835_),
    .X(_2084_));
 sky130_fd_sc_hd__mux2_1 _5399_ (.A0(\sub1.data_o[83] ),
    .A1(_2084_),
    .S(_1837_),
    .X(_2085_));
 sky130_fd_sc_hd__clkbuf_4 _5400_ (.A(_1305_),
    .X(_2086_));
 sky130_fd_sc_hd__a31o_1 _5401_ (.A1(_1793_),
    .A2(\sub1.data_o[83] ),
    .A3(_1849_),
    .B1(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__a21o_1 _5402_ (.A1(_2054_),
    .A2(_2085_),
    .B1(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__clkbuf_4 _5403_ (.A(_1123_),
    .X(_2089_));
 sky130_fd_sc_hd__o21a_1 _5404_ (.A1(\mix1.data_o[83] ),
    .A2(_2089_),
    .B1(_1817_),
    .X(_2090_));
 sky130_fd_sc_hd__a221o_1 _5405_ (.A1(\sub1.data_o[83] ),
    .A2(_1792_),
    .B1(_2088_),
    .B2(_2090_),
    .C1(_2068_),
    .X(_2091_));
 sky130_fd_sc_hd__o21ai_2 _5406_ (.A1(_1812_),
    .A2(_2085_),
    .B1(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(\ks1.key_reg[83] ),
    .A1(net239),
    .S(_1821_),
    .X(_2093_));
 sky130_fd_sc_hd__xnor2_1 _5408_ (.A(_2092_),
    .B(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__mux2_1 _5409_ (.A0(net369),
    .A1(_2094_),
    .S(_2050_),
    .X(_2095_));
 sky130_fd_sc_hd__clkbuf_1 _5410_ (.A(_2095_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _5411_ (.A0(net111),
    .A1(\mix1.data_o[84] ),
    .S(_1835_),
    .X(_2096_));
 sky130_fd_sc_hd__mux2_1 _5412_ (.A0(\sub1.data_o[84] ),
    .A1(_2096_),
    .S(_1837_),
    .X(_2097_));
 sky130_fd_sc_hd__clkbuf_4 _5413_ (.A(_1348_),
    .X(_2098_));
 sky130_fd_sc_hd__a31o_1 _5414_ (.A1(_1793_),
    .A2(\sub1.data_o[84] ),
    .A3(_1849_),
    .B1(_2086_),
    .X(_2099_));
 sky130_fd_sc_hd__a21o_1 _5415_ (.A1(_2054_),
    .A2(_2097_),
    .B1(_2099_),
    .X(_2100_));
 sky130_fd_sc_hd__o21a_1 _5416_ (.A1(\mix1.data_o[84] ),
    .A2(_2089_),
    .B1(_1817_),
    .X(_2101_));
 sky130_fd_sc_hd__a221o_1 _5417_ (.A1(\sub1.data_o[84] ),
    .A2(_2098_),
    .B1(_2100_),
    .B2(_2101_),
    .C1(_2068_),
    .X(_2102_));
 sky130_fd_sc_hd__o21ai_4 _5418_ (.A1(_1812_),
    .A2(_2097_),
    .B1(_2102_),
    .Y(_2103_));
 sky130_fd_sc_hd__mux2_1 _5419_ (.A0(\ks1.key_reg[84] ),
    .A1(net240),
    .S(_1821_),
    .X(_2104_));
 sky130_fd_sc_hd__xnor2_1 _5420_ (.A(_2103_),
    .B(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__mux2_1 _5421_ (.A0(net370),
    .A1(_2105_),
    .S(_2050_),
    .X(_2106_));
 sky130_fd_sc_hd__clkbuf_1 _5422_ (.A(_2106_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _5423_ (.A0(net112),
    .A1(\mix1.data_o[85] ),
    .S(_1835_),
    .X(_2107_));
 sky130_fd_sc_hd__mux2_1 _5424_ (.A0(\sub1.data_o[85] ),
    .A1(_2107_),
    .S(_1837_),
    .X(_2108_));
 sky130_fd_sc_hd__a31o_1 _5425_ (.A1(\sub1.data_o[85] ),
    .A2(_1677_),
    .A3(_1849_),
    .B1(_2086_),
    .X(_2109_));
 sky130_fd_sc_hd__a21o_1 _5426_ (.A1(_2054_),
    .A2(_2108_),
    .B1(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__o21a_1 _5427_ (.A1(\mix1.data_o[85] ),
    .A2(_2089_),
    .B1(_1817_),
    .X(_2111_));
 sky130_fd_sc_hd__a221o_1 _5428_ (.A1(\sub1.data_o[85] ),
    .A2(_2098_),
    .B1(_2110_),
    .B2(_2111_),
    .C1(_2068_),
    .X(_2112_));
 sky130_fd_sc_hd__o21ai_2 _5429_ (.A1(_1812_),
    .A2(_2108_),
    .B1(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__mux2_1 _5430_ (.A0(\ks1.key_reg[85] ),
    .A1(net241),
    .S(_1821_),
    .X(_2114_));
 sky130_fd_sc_hd__xnor2_1 _5431_ (.A(_2113_),
    .B(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__mux2_1 _5432_ (.A0(net371),
    .A1(_2115_),
    .S(_2050_),
    .X(_2116_));
 sky130_fd_sc_hd__clkbuf_1 _5433_ (.A(_2116_),
    .X(_0101_));
 sky130_fd_sc_hd__buf_4 _5434_ (.A(_0678_),
    .X(_2117_));
 sky130_fd_sc_hd__mux2_1 _5435_ (.A0(net113),
    .A1(\mix1.data_o[86] ),
    .S(_1835_),
    .X(_2118_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(\sub1.data_o[86] ),
    .A1(_2118_),
    .S(_1837_),
    .X(_2119_));
 sky130_fd_sc_hd__a31o_1 _5437_ (.A1(\sub1.data_o[86] ),
    .A2(_1677_),
    .A3(_1849_),
    .B1(_2086_),
    .X(_2120_));
 sky130_fd_sc_hd__a21o_1 _5438_ (.A1(_2054_),
    .A2(_2119_),
    .B1(_2120_),
    .X(_2121_));
 sky130_fd_sc_hd__clkbuf_4 _5439_ (.A(_1519_),
    .X(_2122_));
 sky130_fd_sc_hd__o21a_1 _5440_ (.A1(\mix1.data_o[86] ),
    .A2(_2089_),
    .B1(_2122_),
    .X(_2123_));
 sky130_fd_sc_hd__a221o_1 _5441_ (.A1(\sub1.data_o[86] ),
    .A2(_2098_),
    .B1(_2121_),
    .B2(_2123_),
    .C1(_2068_),
    .X(_2124_));
 sky130_fd_sc_hd__o21ai_1 _5442_ (.A1(_2117_),
    .A2(_2119_),
    .B1(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__clkbuf_8 _5443_ (.A(_0674_),
    .X(_2126_));
 sky130_fd_sc_hd__mux2_1 _5444_ (.A0(\ks1.key_reg[86] ),
    .A1(net242),
    .S(_2126_),
    .X(_2127_));
 sky130_fd_sc_hd__xnor2_1 _5445_ (.A(_2125_),
    .B(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hd__mux2_1 _5446_ (.A0(net372),
    .A1(_2128_),
    .S(_2050_),
    .X(_2129_));
 sky130_fd_sc_hd__clkbuf_1 _5447_ (.A(_2129_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _5448_ (.A0(net114),
    .A1(\mix1.data_o[87] ),
    .S(_1835_),
    .X(_2130_));
 sky130_fd_sc_hd__mux2_1 _5449_ (.A0(\sub1.data_o[87] ),
    .A1(_2130_),
    .S(_1837_),
    .X(_2131_));
 sky130_fd_sc_hd__a31o_1 _5450_ (.A1(_1793_),
    .A2(\sub1.data_o[87] ),
    .A3(_1849_),
    .B1(_2086_),
    .X(_2132_));
 sky130_fd_sc_hd__a21o_1 _5451_ (.A1(_2054_),
    .A2(_2131_),
    .B1(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__o21a_1 _5452_ (.A1(\mix1.data_o[87] ),
    .A2(_2089_),
    .B1(_2122_),
    .X(_2134_));
 sky130_fd_sc_hd__a221o_1 _5453_ (.A1(\sub1.data_o[87] ),
    .A2(_2098_),
    .B1(_2133_),
    .B2(_2134_),
    .C1(_2068_),
    .X(_2135_));
 sky130_fd_sc_hd__o21ai_1 _5454_ (.A1(_2117_),
    .A2(_2131_),
    .B1(_2135_),
    .Y(_2136_));
 sky130_fd_sc_hd__mux2_1 _5455_ (.A0(\ks1.key_reg[87] ),
    .A1(net243),
    .S(_2126_),
    .X(_2137_));
 sky130_fd_sc_hd__xnor2_1 _5456_ (.A(_2136_),
    .B(_2137_),
    .Y(_2138_));
 sky130_fd_sc_hd__mux2_1 _5457_ (.A0(net373),
    .A1(_2138_),
    .S(_2050_),
    .X(_2139_));
 sky130_fd_sc_hd__clkbuf_1 _5458_ (.A(_2139_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _5459_ (.A0(net115),
    .A1(\mix1.data_o[88] ),
    .S(_2016_),
    .X(_2140_));
 sky130_fd_sc_hd__mux2_1 _5460_ (.A0(\sub1.data_o[88] ),
    .A1(_2140_),
    .S(_2018_),
    .X(_2141_));
 sky130_fd_sc_hd__a32o_1 _5461_ (.A1(\mix1.data_o[88] ),
    .A2(_1989_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[88] ),
    .X(_2142_));
 sky130_fd_sc_hd__a22o_1 _5462_ (.A1(_2028_),
    .A2(_2141_),
    .B1(_2142_),
    .B2(_2039_),
    .X(_2143_));
 sky130_fd_sc_hd__mux2_1 _5463_ (.A0(\ks1.key_reg[88] ),
    .A1(net244),
    .S(_2024_),
    .X(_2144_));
 sky130_fd_sc_hd__xor2_1 _5464_ (.A(_2143_),
    .B(_2144_),
    .X(_2145_));
 sky130_fd_sc_hd__mux2_1 _5465_ (.A0(net374),
    .A1(_2145_),
    .S(_2050_),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_1 _5466_ (.A(_2146_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _5467_ (.A0(net116),
    .A1(\mix1.data_o[89] ),
    .S(_2016_),
    .X(_2147_));
 sky130_fd_sc_hd__mux2_1 _5468_ (.A0(\sub1.data_o[89] ),
    .A1(_2147_),
    .S(_2018_),
    .X(_2148_));
 sky130_fd_sc_hd__a32o_1 _5469_ (.A1(\mix1.data_o[89] ),
    .A2(_1989_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[89] ),
    .X(_2149_));
 sky130_fd_sc_hd__a22o_1 _5470_ (.A1(_2028_),
    .A2(_2148_),
    .B1(_2149_),
    .B2(_2039_),
    .X(_2150_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(\ks1.key_reg[89] ),
    .A1(net245),
    .S(_2024_),
    .X(_2151_));
 sky130_fd_sc_hd__xor2_1 _5472_ (.A(_2150_),
    .B(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__buf_8 _5473_ (.A(_1510_),
    .X(_2153_));
 sky130_fd_sc_hd__mux2_1 _5474_ (.A0(net375),
    .A1(_2152_),
    .S(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__clkbuf_1 _5475_ (.A(_2154_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _5476_ (.A0(net118),
    .A1(\mix1.data_o[90] ),
    .S(_2016_),
    .X(_2155_));
 sky130_fd_sc_hd__mux2_1 _5477_ (.A0(\sub1.data_o[90] ),
    .A1(_2155_),
    .S(_2018_),
    .X(_2156_));
 sky130_fd_sc_hd__clkbuf_4 _5478_ (.A(_1306_),
    .X(_2157_));
 sky130_fd_sc_hd__a32o_1 _5479_ (.A1(\mix1.data_o[90] ),
    .A2(_2157_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[90] ),
    .X(_2158_));
 sky130_fd_sc_hd__a22o_1 _5480_ (.A1(_2028_),
    .A2(_2156_),
    .B1(_2158_),
    .B2(_2039_),
    .X(_2159_));
 sky130_fd_sc_hd__mux2_2 _5481_ (.A0(\ks1.key_reg[90] ),
    .A1(net247),
    .S(_2024_),
    .X(_2160_));
 sky130_fd_sc_hd__xor2_1 _5482_ (.A(_2159_),
    .B(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__mux2_1 _5483_ (.A0(net377),
    .A1(_2161_),
    .S(_2153_),
    .X(_2162_));
 sky130_fd_sc_hd__clkbuf_1 _5484_ (.A(_2162_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _5485_ (.A0(net119),
    .A1(\mix1.data_o[91] ),
    .S(_2016_),
    .X(_2163_));
 sky130_fd_sc_hd__mux2_1 _5486_ (.A0(\sub1.data_o[91] ),
    .A1(_2163_),
    .S(_2018_),
    .X(_2164_));
 sky130_fd_sc_hd__a32o_1 _5487_ (.A1(\mix1.data_o[91] ),
    .A2(_2157_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[91] ),
    .X(_2165_));
 sky130_fd_sc_hd__a22o_1 _5488_ (.A1(_2028_),
    .A2(_2164_),
    .B1(_2165_),
    .B2(_2039_),
    .X(_2166_));
 sky130_fd_sc_hd__mux2_1 _5489_ (.A0(\ks1.key_reg[91] ),
    .A1(net248),
    .S(_2024_),
    .X(_2167_));
 sky130_fd_sc_hd__xor2_1 _5490_ (.A(_2166_),
    .B(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__mux2_1 _5491_ (.A0(net378),
    .A1(_2168_),
    .S(_2153_),
    .X(_2169_));
 sky130_fd_sc_hd__clkbuf_1 _5492_ (.A(_2169_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _5493_ (.A0(net120),
    .A1(\mix1.data_o[92] ),
    .S(_2016_),
    .X(_2170_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(\sub1.data_o[92] ),
    .A1(_2170_),
    .S(_2018_),
    .X(_2171_));
 sky130_fd_sc_hd__a32o_1 _5495_ (.A1(\mix1.data_o[92] ),
    .A2(_2157_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[92] ),
    .X(_2172_));
 sky130_fd_sc_hd__a22o_1 _5496_ (.A1(_2028_),
    .A2(_2171_),
    .B1(_2172_),
    .B2(_2039_),
    .X(_2173_));
 sky130_fd_sc_hd__mux2_1 _5497_ (.A0(\ks1.key_reg[92] ),
    .A1(net249),
    .S(_2024_),
    .X(_2174_));
 sky130_fd_sc_hd__xor2_1 _5498_ (.A(_2173_),
    .B(_2174_),
    .X(_2175_));
 sky130_fd_sc_hd__mux2_1 _5499_ (.A0(net379),
    .A1(_2175_),
    .S(_2153_),
    .X(_2176_));
 sky130_fd_sc_hd__clkbuf_1 _5500_ (.A(_2176_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _5501_ (.A0(net121),
    .A1(\mix1.data_o[93] ),
    .S(_2016_),
    .X(_2177_));
 sky130_fd_sc_hd__mux2_1 _5502_ (.A0(\sub1.data_o[93] ),
    .A1(_2177_),
    .S(_2018_),
    .X(_2178_));
 sky130_fd_sc_hd__a32o_1 _5503_ (.A1(\mix1.data_o[93] ),
    .A2(_2157_),
    .A3(_2020_),
    .B1(_2021_),
    .B2(\sub1.data_o[93] ),
    .X(_2179_));
 sky130_fd_sc_hd__a22o_1 _5504_ (.A1(_2028_),
    .A2(_2178_),
    .B1(_2179_),
    .B2(_2039_),
    .X(_2180_));
 sky130_fd_sc_hd__mux2_1 _5505_ (.A0(\ks1.key_reg[93] ),
    .A1(net250),
    .S(_2024_),
    .X(_2181_));
 sky130_fd_sc_hd__xor2_1 _5506_ (.A(_2180_),
    .B(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__mux2_1 _5507_ (.A0(net380),
    .A1(_2182_),
    .S(_2153_),
    .X(_2183_));
 sky130_fd_sc_hd__clkbuf_1 _5508_ (.A(_2183_),
    .X(_0109_));
 sky130_fd_sc_hd__buf_4 _5509_ (.A(_1513_),
    .X(_2184_));
 sky130_fd_sc_hd__mux2_1 _5510_ (.A0(net122),
    .A1(\mix1.data_o[94] ),
    .S(_2184_),
    .X(_2185_));
 sky130_fd_sc_hd__buf_4 _5511_ (.A(_1516_),
    .X(_2186_));
 sky130_fd_sc_hd__mux2_1 _5512_ (.A0(\sub1.data_o[94] ),
    .A1(_2185_),
    .S(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__clkbuf_4 _5513_ (.A(_1519_),
    .X(_2188_));
 sky130_fd_sc_hd__clkbuf_4 _5514_ (.A(_1354_),
    .X(_2189_));
 sky130_fd_sc_hd__a32o_1 _5515_ (.A1(\mix1.data_o[94] ),
    .A2(_2157_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[94] ),
    .X(_2190_));
 sky130_fd_sc_hd__a22o_1 _5516_ (.A1(_2028_),
    .A2(_2187_),
    .B1(_2190_),
    .B2(_2039_),
    .X(_2191_));
 sky130_fd_sc_hd__buf_4 _5517_ (.A(_1440_),
    .X(_2192_));
 sky130_fd_sc_hd__mux2_2 _5518_ (.A0(\ks1.key_reg[94] ),
    .A1(net251),
    .S(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__xor2_1 _5519_ (.A(_2191_),
    .B(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__mux2_1 _5520_ (.A0(net381),
    .A1(_2194_),
    .S(_2153_),
    .X(_2195_));
 sky130_fd_sc_hd__clkbuf_1 _5521_ (.A(_2195_),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_4 _5522_ (.A(_1349_),
    .X(_2196_));
 sky130_fd_sc_hd__mux2_1 _5523_ (.A0(net123),
    .A1(\mix1.data_o[95] ),
    .S(_2184_),
    .X(_2197_));
 sky130_fd_sc_hd__mux2_1 _5524_ (.A0(\sub1.data_o[95] ),
    .A1(_2197_),
    .S(_2186_),
    .X(_2198_));
 sky130_fd_sc_hd__a32o_1 _5525_ (.A1(\mix1.data_o[95] ),
    .A2(_2157_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[95] ),
    .X(_2199_));
 sky130_fd_sc_hd__a22o_1 _5526_ (.A1(_2196_),
    .A2(_2198_),
    .B1(_2199_),
    .B2(_2039_),
    .X(_2200_));
 sky130_fd_sc_hd__mux2_1 _5527_ (.A0(\ks1.key_reg[95] ),
    .A1(net252),
    .S(_2192_),
    .X(_2201_));
 sky130_fd_sc_hd__xor2_1 _5528_ (.A(_2200_),
    .B(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__mux2_1 _5529_ (.A0(net382),
    .A1(_2202_),
    .S(_2153_),
    .X(_2203_));
 sky130_fd_sc_hd__clkbuf_1 _5530_ (.A(_2203_),
    .X(_0111_));
 sky130_fd_sc_hd__buf_4 _5531_ (.A(_1337_),
    .X(_2204_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(net124),
    .A1(\mix1.data_o[96] ),
    .S(_2204_),
    .X(_2205_));
 sky130_fd_sc_hd__clkbuf_4 _5533_ (.A(_1344_),
    .X(_2206_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(\sub1.data_o[96] ),
    .A1(_2205_),
    .S(_2206_),
    .X(_2207_));
 sky130_fd_sc_hd__clkbuf_4 _5535_ (.A(_1121_),
    .X(_2208_));
 sky130_fd_sc_hd__a31o_1 _5536_ (.A1(_2208_),
    .A2(\sub1.data_o[96] ),
    .A3(_1849_),
    .B1(_2086_),
    .X(_2209_));
 sky130_fd_sc_hd__a21o_1 _5537_ (.A1(_2054_),
    .A2(_2207_),
    .B1(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__o21a_1 _5538_ (.A1(\mix1.data_o[96] ),
    .A2(_2089_),
    .B1(_2122_),
    .X(_2211_));
 sky130_fd_sc_hd__a221o_1 _5539_ (.A1(\sub1.data_o[96] ),
    .A2(_2098_),
    .B1(_2210_),
    .B2(_2211_),
    .C1(_2068_),
    .X(_2212_));
 sky130_fd_sc_hd__o21ai_1 _5540_ (.A1(_2117_),
    .A2(_2207_),
    .B1(_2212_),
    .Y(_2213_));
 sky130_fd_sc_hd__mux2_2 _5541_ (.A0(\ks1.key_reg[96] ),
    .A1(net253),
    .S(_2126_),
    .X(_2214_));
 sky130_fd_sc_hd__xnor2_1 _5542_ (.A(_2213_),
    .B(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__mux2_1 _5543_ (.A0(net383),
    .A1(_2215_),
    .S(_2153_),
    .X(_2216_));
 sky130_fd_sc_hd__clkbuf_1 _5544_ (.A(_2216_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _5545_ (.A0(net125),
    .A1(\mix1.data_o[97] ),
    .S(_2204_),
    .X(_2217_));
 sky130_fd_sc_hd__mux2_1 _5546_ (.A0(\sub1.data_o[97] ),
    .A1(_2217_),
    .S(_2206_),
    .X(_2218_));
 sky130_fd_sc_hd__a31o_1 _5547_ (.A1(_2208_),
    .A2(\sub1.data_o[97] ),
    .A3(_1849_),
    .B1(_2086_),
    .X(_2219_));
 sky130_fd_sc_hd__a21o_1 _5548_ (.A1(_2054_),
    .A2(_2218_),
    .B1(_2219_),
    .X(_2220_));
 sky130_fd_sc_hd__o21a_1 _5549_ (.A1(\mix1.data_o[97] ),
    .A2(_2089_),
    .B1(_2122_),
    .X(_2221_));
 sky130_fd_sc_hd__a221o_1 _5550_ (.A1(\sub1.data_o[97] ),
    .A2(_2098_),
    .B1(_2220_),
    .B2(_2221_),
    .C1(_2068_),
    .X(_2222_));
 sky130_fd_sc_hd__o21ai_1 _5551_ (.A1(_2117_),
    .A2(_2218_),
    .B1(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__mux2_1 _5552_ (.A0(\ks1.key_reg[97] ),
    .A1(net254),
    .S(_2126_),
    .X(_2224_));
 sky130_fd_sc_hd__xnor2_1 _5553_ (.A(_2223_),
    .B(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__mux2_1 _5554_ (.A0(net384),
    .A1(_2225_),
    .S(_2153_),
    .X(_2226_));
 sky130_fd_sc_hd__clkbuf_1 _5555_ (.A(_2226_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _5556_ (.A0(net126),
    .A1(\mix1.data_o[98] ),
    .S(_2204_),
    .X(_2227_));
 sky130_fd_sc_hd__mux2_1 _5557_ (.A0(\sub1.data_o[98] ),
    .A1(_2227_),
    .S(_2206_),
    .X(_2228_));
 sky130_fd_sc_hd__clkbuf_4 _5558_ (.A(_1122_),
    .X(_2229_));
 sky130_fd_sc_hd__clkbuf_4 _5559_ (.A(_1119_),
    .X(_2230_));
 sky130_fd_sc_hd__a31o_1 _5560_ (.A1(_2208_),
    .A2(\sub1.data_o[98] ),
    .A3(_2230_),
    .B1(_2086_),
    .X(_2231_));
 sky130_fd_sc_hd__a21o_1 _5561_ (.A1(_2229_),
    .A2(_2228_),
    .B1(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__o21a_1 _5562_ (.A1(\mix1.data_o[98] ),
    .A2(_2089_),
    .B1(_2122_),
    .X(_2233_));
 sky130_fd_sc_hd__a221o_1 _5563_ (.A1(\sub1.data_o[98] ),
    .A2(_2098_),
    .B1(_2232_),
    .B2(_2233_),
    .C1(_2068_),
    .X(_2234_));
 sky130_fd_sc_hd__o21ai_2 _5564_ (.A1(_2117_),
    .A2(_2228_),
    .B1(_2234_),
    .Y(_2235_));
 sky130_fd_sc_hd__mux2_1 _5565_ (.A0(\ks1.key_reg[98] ),
    .A1(net255),
    .S(_2126_),
    .X(_2236_));
 sky130_fd_sc_hd__xnor2_1 _5566_ (.A(_2235_),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__mux2_1 _5567_ (.A0(net385),
    .A1(_2237_),
    .S(_2153_),
    .X(_2238_));
 sky130_fd_sc_hd__clkbuf_1 _5568_ (.A(_2238_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _5569_ (.A0(net127),
    .A1(\mix1.data_o[99] ),
    .S(_2204_),
    .X(_2239_));
 sky130_fd_sc_hd__mux2_1 _5570_ (.A0(\sub1.data_o[99] ),
    .A1(_2239_),
    .S(_2206_),
    .X(_2240_));
 sky130_fd_sc_hd__a31o_1 _5571_ (.A1(_2208_),
    .A2(\sub1.data_o[99] ),
    .A3(_2230_),
    .B1(_2086_),
    .X(_2241_));
 sky130_fd_sc_hd__a21o_1 _5572_ (.A1(_2229_),
    .A2(_2240_),
    .B1(_2241_),
    .X(_2242_));
 sky130_fd_sc_hd__o21a_1 _5573_ (.A1(\mix1.data_o[99] ),
    .A2(_2089_),
    .B1(_2122_),
    .X(_2243_));
 sky130_fd_sc_hd__clkbuf_4 _5574_ (.A(_1114_),
    .X(_2244_));
 sky130_fd_sc_hd__a221o_1 _5575_ (.A1(\sub1.data_o[99] ),
    .A2(_2098_),
    .B1(_2242_),
    .B2(_2243_),
    .C1(_2244_),
    .X(_2245_));
 sky130_fd_sc_hd__o21ai_1 _5576_ (.A1(_2117_),
    .A2(_2240_),
    .B1(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__mux2_2 _5577_ (.A0(\ks1.key_reg[99] ),
    .A1(net256),
    .S(_2126_),
    .X(_2247_));
 sky130_fd_sc_hd__xnor2_1 _5578_ (.A(_2246_),
    .B(_2247_),
    .Y(_2248_));
 sky130_fd_sc_hd__buf_6 _5579_ (.A(_1510_),
    .X(_2249_));
 sky130_fd_sc_hd__mux2_1 _5580_ (.A0(net386),
    .A1(_2248_),
    .S(_2249_),
    .X(_2250_));
 sky130_fd_sc_hd__clkbuf_1 _5581_ (.A(_2250_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _5582_ (.A0(net2),
    .A1(\mix1.data_o[100] ),
    .S(_2204_),
    .X(_2251_));
 sky130_fd_sc_hd__mux2_1 _5583_ (.A0(\sub1.data_o[100] ),
    .A1(_2251_),
    .S(_2206_),
    .X(_2252_));
 sky130_fd_sc_hd__a31o_1 _5584_ (.A1(_2208_),
    .A2(\sub1.data_o[100] ),
    .A3(_2230_),
    .B1(_2086_),
    .X(_2253_));
 sky130_fd_sc_hd__a21o_1 _5585_ (.A1(_2229_),
    .A2(_2252_),
    .B1(_2253_),
    .X(_2254_));
 sky130_fd_sc_hd__o21a_1 _5586_ (.A1(\mix1.data_o[100] ),
    .A2(_2089_),
    .B1(_2122_),
    .X(_2255_));
 sky130_fd_sc_hd__a221o_1 _5587_ (.A1(\sub1.data_o[100] ),
    .A2(_2098_),
    .B1(_2254_),
    .B2(_2255_),
    .C1(_2244_),
    .X(_2256_));
 sky130_fd_sc_hd__o21ai_4 _5588_ (.A1(_2117_),
    .A2(_2252_),
    .B1(_2256_),
    .Y(_2257_));
 sky130_fd_sc_hd__mux2_2 _5589_ (.A0(\ks1.key_reg[100] ),
    .A1(net131),
    .S(_2126_),
    .X(_2258_));
 sky130_fd_sc_hd__xnor2_1 _5590_ (.A(_2257_),
    .B(_2258_),
    .Y(_2259_));
 sky130_fd_sc_hd__mux2_1 _5591_ (.A0(net261),
    .A1(_2259_),
    .S(_2249_),
    .X(_2260_));
 sky130_fd_sc_hd__clkbuf_1 _5592_ (.A(_2260_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _5593_ (.A0(net3),
    .A1(\mix1.data_o[101] ),
    .S(_2204_),
    .X(_2261_));
 sky130_fd_sc_hd__mux2_1 _5594_ (.A0(\sub1.data_o[101] ),
    .A1(_2261_),
    .S(_2206_),
    .X(_2262_));
 sky130_fd_sc_hd__clkbuf_4 _5595_ (.A(_1305_),
    .X(_2263_));
 sky130_fd_sc_hd__a31o_1 _5596_ (.A1(\sub1.data_o[101] ),
    .A2(_1677_),
    .A3(_2230_),
    .B1(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__a21o_1 _5597_ (.A1(_2229_),
    .A2(_2262_),
    .B1(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__clkbuf_4 _5598_ (.A(_1123_),
    .X(_2266_));
 sky130_fd_sc_hd__o21a_1 _5599_ (.A1(\mix1.data_o[101] ),
    .A2(_2266_),
    .B1(_2122_),
    .X(_2267_));
 sky130_fd_sc_hd__a221o_1 _5600_ (.A1(\sub1.data_o[101] ),
    .A2(_2098_),
    .B1(_2265_),
    .B2(_2267_),
    .C1(_2244_),
    .X(_2268_));
 sky130_fd_sc_hd__o21ai_4 _5601_ (.A1(_2117_),
    .A2(_2262_),
    .B1(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__mux2_2 _5602_ (.A0(\ks1.key_reg[101] ),
    .A1(net132),
    .S(_2126_),
    .X(_2270_));
 sky130_fd_sc_hd__xnor2_1 _5603_ (.A(_2269_),
    .B(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__mux2_1 _5604_ (.A0(net262),
    .A1(_2271_),
    .S(_2249_),
    .X(_2272_));
 sky130_fd_sc_hd__clkbuf_1 _5605_ (.A(_2272_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _5606_ (.A0(net4),
    .A1(\mix1.data_o[102] ),
    .S(_2204_),
    .X(_2273_));
 sky130_fd_sc_hd__mux2_1 _5607_ (.A0(\sub1.data_o[102] ),
    .A1(_2273_),
    .S(_2206_),
    .X(_2274_));
 sky130_fd_sc_hd__clkbuf_4 _5608_ (.A(_1348_),
    .X(_2275_));
 sky130_fd_sc_hd__a31o_1 _5609_ (.A1(\sub1.data_o[102] ),
    .A2(_1677_),
    .A3(_2230_),
    .B1(_2263_),
    .X(_2276_));
 sky130_fd_sc_hd__a21o_1 _5610_ (.A1(_2229_),
    .A2(_2274_),
    .B1(_2276_),
    .X(_2277_));
 sky130_fd_sc_hd__o21a_1 _5611_ (.A1(\mix1.data_o[102] ),
    .A2(_2266_),
    .B1(_2122_),
    .X(_2278_));
 sky130_fd_sc_hd__a221o_1 _5612_ (.A1(\sub1.data_o[102] ),
    .A2(_2275_),
    .B1(_2277_),
    .B2(_2278_),
    .C1(_2244_),
    .X(_2279_));
 sky130_fd_sc_hd__o21ai_1 _5613_ (.A1(_2117_),
    .A2(_2274_),
    .B1(_2279_),
    .Y(_2280_));
 sky130_fd_sc_hd__mux2_1 _5614_ (.A0(\ks1.key_reg[102] ),
    .A1(net133),
    .S(_2126_),
    .X(_2281_));
 sky130_fd_sc_hd__xnor2_1 _5615_ (.A(_2280_),
    .B(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__mux2_1 _5616_ (.A0(net263),
    .A1(_2282_),
    .S(_2249_),
    .X(_2283_));
 sky130_fd_sc_hd__clkbuf_1 _5617_ (.A(_2283_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _5618_ (.A0(net5),
    .A1(\mix1.data_o[103] ),
    .S(_2204_),
    .X(_2284_));
 sky130_fd_sc_hd__mux2_1 _5619_ (.A0(\sub1.data_o[103] ),
    .A1(_2284_),
    .S(_2206_),
    .X(_2285_));
 sky130_fd_sc_hd__a31o_1 _5620_ (.A1(\sub1.data_o[103] ),
    .A2(_1121_),
    .A3(_2230_),
    .B1(_2263_),
    .X(_2286_));
 sky130_fd_sc_hd__a21o_1 _5621_ (.A1(_2229_),
    .A2(_2285_),
    .B1(_2286_),
    .X(_2287_));
 sky130_fd_sc_hd__o21a_1 _5622_ (.A1(\mix1.data_o[103] ),
    .A2(_2266_),
    .B1(_2122_),
    .X(_2288_));
 sky130_fd_sc_hd__a221o_1 _5623_ (.A1(\sub1.data_o[103] ),
    .A2(_2275_),
    .B1(_2287_),
    .B2(_2288_),
    .C1(_2244_),
    .X(_2289_));
 sky130_fd_sc_hd__o21ai_1 _5624_ (.A1(_2117_),
    .A2(_2285_),
    .B1(_2289_),
    .Y(_2290_));
 sky130_fd_sc_hd__mux2_2 _5625_ (.A0(\ks1.key_reg[103] ),
    .A1(net134),
    .S(_2126_),
    .X(_2291_));
 sky130_fd_sc_hd__xnor2_1 _5626_ (.A(_2290_),
    .B(_2291_),
    .Y(_2292_));
 sky130_fd_sc_hd__mux2_1 _5627_ (.A0(net264),
    .A1(_2292_),
    .S(_2249_),
    .X(_2293_));
 sky130_fd_sc_hd__clkbuf_1 _5628_ (.A(_2293_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _5629_ (.A0(net6),
    .A1(\mix1.data_o[104] ),
    .S(_2184_),
    .X(_2294_));
 sky130_fd_sc_hd__mux2_1 _5630_ (.A0(\sub1.data_o[104] ),
    .A1(_2294_),
    .S(_2186_),
    .X(_2295_));
 sky130_fd_sc_hd__a32o_1 _5631_ (.A1(\mix1.data_o[104] ),
    .A2(_2157_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[104] ),
    .X(_2296_));
 sky130_fd_sc_hd__clkbuf_4 _5632_ (.A(_0677_),
    .X(_2297_));
 sky130_fd_sc_hd__a22o_1 _5633_ (.A1(_2196_),
    .A2(_2295_),
    .B1(_2296_),
    .B2(_2297_),
    .X(_2298_));
 sky130_fd_sc_hd__mux2_1 _5634_ (.A0(\ks1.key_reg[104] ),
    .A1(net135),
    .S(_2192_),
    .X(_2299_));
 sky130_fd_sc_hd__xor2_1 _5635_ (.A(_2298_),
    .B(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__mux2_1 _5636_ (.A0(net265),
    .A1(_2300_),
    .S(_2249_),
    .X(_2301_));
 sky130_fd_sc_hd__clkbuf_1 _5637_ (.A(_2301_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _5638_ (.A0(net7),
    .A1(\mix1.data_o[105] ),
    .S(_2184_),
    .X(_2302_));
 sky130_fd_sc_hd__mux2_1 _5639_ (.A0(\sub1.data_o[105] ),
    .A1(_2302_),
    .S(_2186_),
    .X(_2303_));
 sky130_fd_sc_hd__a32o_1 _5640_ (.A1(\mix1.data_o[105] ),
    .A2(_2157_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[105] ),
    .X(_2304_));
 sky130_fd_sc_hd__a22o_1 _5641_ (.A1(_2196_),
    .A2(_2303_),
    .B1(_2304_),
    .B2(_2297_),
    .X(_2305_));
 sky130_fd_sc_hd__mux2_1 _5642_ (.A0(\ks1.key_reg[105] ),
    .A1(net136),
    .S(_2192_),
    .X(_2306_));
 sky130_fd_sc_hd__xor2_1 _5643_ (.A(_2305_),
    .B(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__mux2_1 _5644_ (.A0(net266),
    .A1(_2307_),
    .S(_2249_),
    .X(_2308_));
 sky130_fd_sc_hd__clkbuf_1 _5645_ (.A(_2308_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _5646_ (.A0(net8),
    .A1(\mix1.data_o[106] ),
    .S(_2184_),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_1 _5647_ (.A0(\sub1.data_o[106] ),
    .A1(_2309_),
    .S(_2186_),
    .X(_2310_));
 sky130_fd_sc_hd__a32o_1 _5648_ (.A1(\mix1.data_o[106] ),
    .A2(_2157_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[106] ),
    .X(_2311_));
 sky130_fd_sc_hd__a22o_1 _5649_ (.A1(_2196_),
    .A2(_2310_),
    .B1(_2311_),
    .B2(_2297_),
    .X(_2312_));
 sky130_fd_sc_hd__mux2_2 _5650_ (.A0(\ks1.key_reg[106] ),
    .A1(net137),
    .S(_2192_),
    .X(_2313_));
 sky130_fd_sc_hd__xor2_1 _5651_ (.A(_2312_),
    .B(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__mux2_1 _5652_ (.A0(net267),
    .A1(_2314_),
    .S(_2249_),
    .X(_2315_));
 sky130_fd_sc_hd__clkbuf_1 _5653_ (.A(_2315_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _5654_ (.A0(net9),
    .A1(\mix1.data_o[107] ),
    .S(_2184_),
    .X(_2316_));
 sky130_fd_sc_hd__mux2_1 _5655_ (.A0(\sub1.data_o[107] ),
    .A1(_2316_),
    .S(_2186_),
    .X(_2317_));
 sky130_fd_sc_hd__a32o_1 _5656_ (.A1(\mix1.data_o[107] ),
    .A2(_2157_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[107] ),
    .X(_2318_));
 sky130_fd_sc_hd__a22o_1 _5657_ (.A1(_2196_),
    .A2(_2317_),
    .B1(_2318_),
    .B2(_2297_),
    .X(_2319_));
 sky130_fd_sc_hd__mux2_2 _5658_ (.A0(\ks1.key_reg[107] ),
    .A1(net138),
    .S(_2192_),
    .X(_2320_));
 sky130_fd_sc_hd__xor2_1 _5659_ (.A(_2319_),
    .B(_2320_),
    .X(_2321_));
 sky130_fd_sc_hd__mux2_1 _5660_ (.A0(net268),
    .A1(_2321_),
    .S(_2249_),
    .X(_2322_));
 sky130_fd_sc_hd__clkbuf_1 _5661_ (.A(_2322_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _5662_ (.A0(net10),
    .A1(\mix1.data_o[108] ),
    .S(_2184_),
    .X(_2323_));
 sky130_fd_sc_hd__mux2_1 _5663_ (.A0(\sub1.data_o[108] ),
    .A1(_2323_),
    .S(_2186_),
    .X(_2324_));
 sky130_fd_sc_hd__clkbuf_4 _5664_ (.A(_1618_),
    .X(_2325_));
 sky130_fd_sc_hd__a32o_1 _5665_ (.A1(\mix1.data_o[108] ),
    .A2(_2325_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[108] ),
    .X(_2326_));
 sky130_fd_sc_hd__a22o_1 _5666_ (.A1(_2196_),
    .A2(_2324_),
    .B1(_2326_),
    .B2(_2297_),
    .X(_2327_));
 sky130_fd_sc_hd__mux2_2 _5667_ (.A0(\ks1.key_reg[108] ),
    .A1(net139),
    .S(_2192_),
    .X(_2328_));
 sky130_fd_sc_hd__xor2_1 _5668_ (.A(_2327_),
    .B(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__mux2_1 _5669_ (.A0(net269),
    .A1(_2329_),
    .S(_2249_),
    .X(_2330_));
 sky130_fd_sc_hd__clkbuf_1 _5670_ (.A(_2330_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _5671_ (.A0(net11),
    .A1(\mix1.data_o[109] ),
    .S(_2184_),
    .X(_2331_));
 sky130_fd_sc_hd__mux2_1 _5672_ (.A0(\sub1.data_o[109] ),
    .A1(_2331_),
    .S(_2186_),
    .X(_2332_));
 sky130_fd_sc_hd__a32o_1 _5673_ (.A1(\mix1.data_o[109] ),
    .A2(_2325_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[109] ),
    .X(_2333_));
 sky130_fd_sc_hd__a22o_1 _5674_ (.A1(_2196_),
    .A2(_2332_),
    .B1(_2333_),
    .B2(_2297_),
    .X(_2334_));
 sky130_fd_sc_hd__mux2_1 _5675_ (.A0(\ks1.key_reg[109] ),
    .A1(net140),
    .S(_2192_),
    .X(_2335_));
 sky130_fd_sc_hd__xor2_1 _5676_ (.A(_2334_),
    .B(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__buf_8 _5677_ (.A(_1510_),
    .X(_2337_));
 sky130_fd_sc_hd__mux2_1 _5678_ (.A0(net270),
    .A1(_2336_),
    .S(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__clkbuf_1 _5679_ (.A(_2338_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _5680_ (.A0(net13),
    .A1(\mix1.data_o[110] ),
    .S(_2184_),
    .X(_2339_));
 sky130_fd_sc_hd__mux2_1 _5681_ (.A0(\sub1.data_o[110] ),
    .A1(_2339_),
    .S(_2186_),
    .X(_2340_));
 sky130_fd_sc_hd__a32o_1 _5682_ (.A1(\mix1.data_o[110] ),
    .A2(_2325_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[110] ),
    .X(_2341_));
 sky130_fd_sc_hd__a22o_1 _5683_ (.A1(_2196_),
    .A2(_2340_),
    .B1(_2341_),
    .B2(_2297_),
    .X(_2342_));
 sky130_fd_sc_hd__mux2_1 _5684_ (.A0(\ks1.key_reg[110] ),
    .A1(net142),
    .S(_2192_),
    .X(_2343_));
 sky130_fd_sc_hd__xor2_1 _5685_ (.A(_2342_),
    .B(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__mux2_1 _5686_ (.A0(net272),
    .A1(_2344_),
    .S(_2337_),
    .X(_2345_));
 sky130_fd_sc_hd__clkbuf_1 _5687_ (.A(_2345_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _5688_ (.A0(net14),
    .A1(\mix1.data_o[111] ),
    .S(_2184_),
    .X(_2346_));
 sky130_fd_sc_hd__mux2_1 _5689_ (.A0(\sub1.data_o[111] ),
    .A1(_2346_),
    .S(_2186_),
    .X(_2347_));
 sky130_fd_sc_hd__a32o_1 _5690_ (.A1(\mix1.data_o[111] ),
    .A2(_2325_),
    .A3(_2188_),
    .B1(_2189_),
    .B2(\sub1.data_o[111] ),
    .X(_2348_));
 sky130_fd_sc_hd__a22o_1 _5691_ (.A1(_2196_),
    .A2(_2347_),
    .B1(_2348_),
    .B2(_2297_),
    .X(_2349_));
 sky130_fd_sc_hd__mux2_2 _5692_ (.A0(\ks1.key_reg[111] ),
    .A1(net143),
    .S(_2192_),
    .X(_2350_));
 sky130_fd_sc_hd__xor2_1 _5693_ (.A(_2349_),
    .B(_2350_),
    .X(_2351_));
 sky130_fd_sc_hd__mux2_1 _5694_ (.A0(net273),
    .A1(_2351_),
    .S(_2337_),
    .X(_2352_));
 sky130_fd_sc_hd__clkbuf_1 _5695_ (.A(_2352_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _5696_ (.A0(net15),
    .A1(\mix1.data_o[112] ),
    .S(_2204_),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _5697_ (.A0(\sub1.data_o[112] ),
    .A1(_2353_),
    .S(_2206_),
    .X(_2354_));
 sky130_fd_sc_hd__a31o_1 _5698_ (.A1(_2208_),
    .A2(_1120_),
    .A3(\sub1.data_o[112] ),
    .B1(_2263_),
    .X(_2355_));
 sky130_fd_sc_hd__a21o_1 _5699_ (.A1(_2229_),
    .A2(_2354_),
    .B1(_2355_),
    .X(_2356_));
 sky130_fd_sc_hd__o21a_1 _5700_ (.A1(\mix1.data_o[112] ),
    .A2(_2266_),
    .B1(_1352_),
    .X(_2357_));
 sky130_fd_sc_hd__a221o_1 _5701_ (.A1(\sub1.data_o[112] ),
    .A2(_2275_),
    .B1(_2356_),
    .B2(_2357_),
    .C1(_2244_),
    .X(_2358_));
 sky130_fd_sc_hd__o21ai_4 _5702_ (.A1(_1358_),
    .A2(_2354_),
    .B1(_2358_),
    .Y(_2359_));
 sky130_fd_sc_hd__mux2_2 _5703_ (.A0(\ks1.key_reg[112] ),
    .A1(net144),
    .S(_0675_),
    .X(_2360_));
 sky130_fd_sc_hd__xnor2_1 _5704_ (.A(_2359_),
    .B(_2360_),
    .Y(_2361_));
 sky130_fd_sc_hd__mux2_1 _5705_ (.A0(net274),
    .A1(_2361_),
    .S(_2337_),
    .X(_2362_));
 sky130_fd_sc_hd__clkbuf_1 _5706_ (.A(_2362_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _5707_ (.A0(net16),
    .A1(\mix1.data_o[113] ),
    .S(_2204_),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_1 _5708_ (.A0(\sub1.data_o[113] ),
    .A1(_2363_),
    .S(_2206_),
    .X(_2364_));
 sky130_fd_sc_hd__a31o_1 _5709_ (.A1(_2208_),
    .A2(\sub1.data_o[113] ),
    .A3(_2230_),
    .B1(_2263_),
    .X(_2365_));
 sky130_fd_sc_hd__a21o_1 _5710_ (.A1(_2229_),
    .A2(_2364_),
    .B1(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__o21a_1 _5711_ (.A1(\mix1.data_o[113] ),
    .A2(_2266_),
    .B1(_1352_),
    .X(_2367_));
 sky130_fd_sc_hd__a221o_1 _5712_ (.A1(\sub1.data_o[113] ),
    .A2(_2275_),
    .B1(_2366_),
    .B2(_2367_),
    .C1(_2244_),
    .X(_2368_));
 sky130_fd_sc_hd__o21ai_1 _5713_ (.A1(_1358_),
    .A2(_2364_),
    .B1(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__mux2_2 _5714_ (.A0(\ks1.key_reg[113] ),
    .A1(net145),
    .S(_0675_),
    .X(_2370_));
 sky130_fd_sc_hd__xnor2_1 _5715_ (.A(_2369_),
    .B(_2370_),
    .Y(_2371_));
 sky130_fd_sc_hd__mux2_1 _5716_ (.A0(net275),
    .A1(_2371_),
    .S(_2337_),
    .X(_2372_));
 sky130_fd_sc_hd__clkbuf_1 _5717_ (.A(_2372_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(net17),
    .A1(\mix1.data_o[114] ),
    .S(_1337_),
    .X(_2373_));
 sky130_fd_sc_hd__mux2_1 _5719_ (.A0(\sub1.data_o[114] ),
    .A1(_2373_),
    .S(_1344_),
    .X(_2374_));
 sky130_fd_sc_hd__a31o_1 _5720_ (.A1(_2208_),
    .A2(\sub1.data_o[114] ),
    .A3(_2230_),
    .B1(_2263_),
    .X(_2375_));
 sky130_fd_sc_hd__a21o_1 _5721_ (.A1(_2229_),
    .A2(_2374_),
    .B1(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__o21a_1 _5722_ (.A1(\mix1.data_o[114] ),
    .A2(_2266_),
    .B1(_1352_),
    .X(_2377_));
 sky130_fd_sc_hd__a221o_1 _5723_ (.A1(\sub1.data_o[114] ),
    .A2(_2275_),
    .B1(_2376_),
    .B2(_2377_),
    .C1(_2244_),
    .X(_2378_));
 sky130_fd_sc_hd__o21ai_1 _5724_ (.A1(_1358_),
    .A2(_2374_),
    .B1(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__mux2_2 _5725_ (.A0(\ks1.key_reg[114] ),
    .A1(net146),
    .S(_0675_),
    .X(_2380_));
 sky130_fd_sc_hd__xnor2_1 _5726_ (.A(_2379_),
    .B(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__mux2_1 _5727_ (.A0(net276),
    .A1(_2381_),
    .S(_2337_),
    .X(_2382_));
 sky130_fd_sc_hd__clkbuf_1 _5728_ (.A(_2382_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _5729_ (.A0(net18),
    .A1(\mix1.data_o[115] ),
    .S(_1337_),
    .X(_2383_));
 sky130_fd_sc_hd__mux2_1 _5730_ (.A0(\sub1.data_o[115] ),
    .A1(_2383_),
    .S(_1344_),
    .X(_2384_));
 sky130_fd_sc_hd__a31o_1 _5731_ (.A1(_2208_),
    .A2(\sub1.data_o[115] ),
    .A3(_2230_),
    .B1(_2263_),
    .X(_2385_));
 sky130_fd_sc_hd__a21o_1 _5732_ (.A1(_2229_),
    .A2(_2384_),
    .B1(_2385_),
    .X(_2386_));
 sky130_fd_sc_hd__o21a_1 _5733_ (.A1(\mix1.data_o[115] ),
    .A2(_2266_),
    .B1(_1352_),
    .X(_2387_));
 sky130_fd_sc_hd__a221o_1 _5734_ (.A1(\sub1.data_o[115] ),
    .A2(_2275_),
    .B1(_2386_),
    .B2(_2387_),
    .C1(_2244_),
    .X(_2388_));
 sky130_fd_sc_hd__o21ai_2 _5735_ (.A1(_1358_),
    .A2(_2384_),
    .B1(_2388_),
    .Y(_2389_));
 sky130_fd_sc_hd__mux2_1 _5736_ (.A0(\ks1.key_reg[115] ),
    .A1(net147),
    .S(_0675_),
    .X(_2390_));
 sky130_fd_sc_hd__xnor2_1 _5737_ (.A(_2389_),
    .B(_2390_),
    .Y(_2391_));
 sky130_fd_sc_hd__mux2_1 _5738_ (.A0(net277),
    .A1(_2391_),
    .S(_2337_),
    .X(_2392_));
 sky130_fd_sc_hd__clkbuf_1 _5739_ (.A(_2392_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _5740_ (.A0(net19),
    .A1(\mix1.data_o[116] ),
    .S(_1337_),
    .X(_2393_));
 sky130_fd_sc_hd__mux2_1 _5741_ (.A0(\sub1.data_o[116] ),
    .A1(_2393_),
    .S(_1344_),
    .X(_2394_));
 sky130_fd_sc_hd__a31o_1 _5742_ (.A1(_2208_),
    .A2(\sub1.data_o[116] ),
    .A3(_2230_),
    .B1(_2263_),
    .X(_2395_));
 sky130_fd_sc_hd__a21o_1 _5743_ (.A1(_1122_),
    .A2(_2394_),
    .B1(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__o21a_1 _5744_ (.A1(\mix1.data_o[116] ),
    .A2(_2266_),
    .B1(_1352_),
    .X(_2397_));
 sky130_fd_sc_hd__a221o_1 _5745_ (.A1(\sub1.data_o[116] ),
    .A2(_2275_),
    .B1(_2396_),
    .B2(_2397_),
    .C1(_2244_),
    .X(_2398_));
 sky130_fd_sc_hd__o21ai_1 _5746_ (.A1(_1358_),
    .A2(_2394_),
    .B1(_2398_),
    .Y(_2399_));
 sky130_fd_sc_hd__mux2_4 _5747_ (.A0(\ks1.key_reg[116] ),
    .A1(net148),
    .S(_0675_),
    .X(_2400_));
 sky130_fd_sc_hd__xnor2_1 _5748_ (.A(_2399_),
    .B(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__mux2_1 _5749_ (.A0(net278),
    .A1(_2401_),
    .S(_2337_),
    .X(_2402_));
 sky130_fd_sc_hd__clkbuf_1 _5750_ (.A(_2402_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _5751_ (.A0(net20),
    .A1(\mix1.data_o[117] ),
    .S(_1337_),
    .X(_2403_));
 sky130_fd_sc_hd__mux2_1 _5752_ (.A0(\sub1.data_o[117] ),
    .A1(_2403_),
    .S(_1344_),
    .X(_2404_));
 sky130_fd_sc_hd__a31o_1 _5753_ (.A1(\sub1.data_o[117] ),
    .A2(_1121_),
    .A3(_1119_),
    .B1(_2263_),
    .X(_2405_));
 sky130_fd_sc_hd__a21o_1 _5754_ (.A1(_1122_),
    .A2(_2404_),
    .B1(_2405_),
    .X(_2406_));
 sky130_fd_sc_hd__o21a_1 _5755_ (.A1(\mix1.data_o[117] ),
    .A2(_2266_),
    .B1(_1352_),
    .X(_2407_));
 sky130_fd_sc_hd__a221o_1 _5756_ (.A1(\sub1.data_o[117] ),
    .A2(_2275_),
    .B1(_2406_),
    .B2(_2407_),
    .C1(_1114_),
    .X(_2408_));
 sky130_fd_sc_hd__o21ai_4 _5757_ (.A1(_1358_),
    .A2(_2404_),
    .B1(_2408_),
    .Y(_2409_));
 sky130_fd_sc_hd__mux2_1 _5758_ (.A0(\ks1.key_reg[117] ),
    .A1(net149),
    .S(_0675_),
    .X(_2410_));
 sky130_fd_sc_hd__xnor2_1 _5759_ (.A(_2409_),
    .B(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__mux2_1 _5760_ (.A0(net279),
    .A1(_2411_),
    .S(_2337_),
    .X(_2412_));
 sky130_fd_sc_hd__clkbuf_1 _5761_ (.A(_2412_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _5762_ (.A0(net21),
    .A1(\mix1.data_o[118] ),
    .S(_1337_),
    .X(_2413_));
 sky130_fd_sc_hd__mux2_1 _5763_ (.A0(\sub1.data_o[118] ),
    .A1(_2413_),
    .S(_1344_),
    .X(_2414_));
 sky130_fd_sc_hd__a31o_1 _5764_ (.A1(\sub1.data_o[118] ),
    .A2(_1121_),
    .A3(_1119_),
    .B1(_2263_),
    .X(_2415_));
 sky130_fd_sc_hd__a21o_1 _5765_ (.A1(_1122_),
    .A2(_2414_),
    .B1(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__o21a_1 _5766_ (.A1(\mix1.data_o[118] ),
    .A2(_2266_),
    .B1(_1352_),
    .X(_2417_));
 sky130_fd_sc_hd__a221o_1 _5767_ (.A1(\sub1.data_o[118] ),
    .A2(_2275_),
    .B1(_2416_),
    .B2(_2417_),
    .C1(_1114_),
    .X(_2418_));
 sky130_fd_sc_hd__o21ai_1 _5768_ (.A1(_1358_),
    .A2(_2414_),
    .B1(_2418_),
    .Y(_2419_));
 sky130_fd_sc_hd__mux2_2 _5769_ (.A0(\ks1.key_reg[118] ),
    .A1(net150),
    .S(_0675_),
    .X(_2420_));
 sky130_fd_sc_hd__xnor2_1 _5770_ (.A(_2419_),
    .B(_2420_),
    .Y(_2421_));
 sky130_fd_sc_hd__mux2_1 _5771_ (.A0(net280),
    .A1(_2421_),
    .S(_2337_),
    .X(_2422_));
 sky130_fd_sc_hd__clkbuf_1 _5772_ (.A(_2422_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _5773_ (.A0(net22),
    .A1(\mix1.data_o[119] ),
    .S(_1337_),
    .X(_2423_));
 sky130_fd_sc_hd__mux2_1 _5774_ (.A0(\sub1.data_o[119] ),
    .A1(_2423_),
    .S(_1344_),
    .X(_2424_));
 sky130_fd_sc_hd__a31o_1 _5775_ (.A1(_1677_),
    .A2(\sub1.data_o[119] ),
    .A3(_1119_),
    .B1(_1305_),
    .X(_2425_));
 sky130_fd_sc_hd__a21o_1 _5776_ (.A1(_1122_),
    .A2(_2424_),
    .B1(_2425_),
    .X(_2426_));
 sky130_fd_sc_hd__o21a_1 _5777_ (.A1(\mix1.data_o[119] ),
    .A2(_1123_),
    .B1(_1352_),
    .X(_2427_));
 sky130_fd_sc_hd__a221o_1 _5778_ (.A1(\sub1.data_o[119] ),
    .A2(_2275_),
    .B1(_2426_),
    .B2(_2427_),
    .C1(_1114_),
    .X(_2428_));
 sky130_fd_sc_hd__o21ai_2 _5779_ (.A1(_1358_),
    .A2(_2424_),
    .B1(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__mux2_1 _5780_ (.A0(\ks1.key_reg[119] ),
    .A1(net151),
    .S(_0675_),
    .X(_2430_));
 sky130_fd_sc_hd__xnor2_1 _5781_ (.A(_2429_),
    .B(_2430_),
    .Y(_2431_));
 sky130_fd_sc_hd__mux2_1 _5782_ (.A0(net281),
    .A1(_2431_),
    .S(_1429_),
    .X(_2432_));
 sky130_fd_sc_hd__clkbuf_1 _5783_ (.A(_2432_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _5784_ (.A0(net24),
    .A1(\mix1.data_o[120] ),
    .S(_1338_),
    .X(_2433_));
 sky130_fd_sc_hd__mux2_1 _5785_ (.A0(\sub1.data_o[120] ),
    .A1(_2433_),
    .S(_1345_),
    .X(_2434_));
 sky130_fd_sc_hd__a32o_1 _5786_ (.A1(\mix1.data_o[120] ),
    .A2(_2325_),
    .A3(_1621_),
    .B1(_1355_),
    .B2(\sub1.data_o[120] ),
    .X(_2435_));
 sky130_fd_sc_hd__a22o_1 _5787_ (.A1(_2196_),
    .A2(_2434_),
    .B1(_2435_),
    .B2(_2297_),
    .X(_2436_));
 sky130_fd_sc_hd__mux2_2 _5788_ (.A0(\ks1.key_reg[120] ),
    .A1(net153),
    .S(_1625_),
    .X(_2437_));
 sky130_fd_sc_hd__xor2_1 _5789_ (.A(_2436_),
    .B(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__mux2_1 _5790_ (.A0(net283),
    .A1(_2438_),
    .S(_1429_),
    .X(_2439_));
 sky130_fd_sc_hd__clkbuf_1 _5791_ (.A(_2439_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _5792_ (.A0(net25),
    .A1(\mix1.data_o[121] ),
    .S(_1338_),
    .X(_2440_));
 sky130_fd_sc_hd__mux2_1 _5793_ (.A0(\sub1.data_o[121] ),
    .A1(_2440_),
    .S(_1345_),
    .X(_2441_));
 sky130_fd_sc_hd__a32o_1 _5794_ (.A1(\mix1.data_o[121] ),
    .A2(_2325_),
    .A3(_1621_),
    .B1(_1355_),
    .B2(\sub1.data_o[121] ),
    .X(_2442_));
 sky130_fd_sc_hd__a22o_1 _5795_ (.A1(_1350_),
    .A2(_2441_),
    .B1(_2442_),
    .B2(_2297_),
    .X(_2443_));
 sky130_fd_sc_hd__mux2_1 _5796_ (.A0(\ks1.key_reg[121] ),
    .A1(net154),
    .S(_1625_),
    .X(_2444_));
 sky130_fd_sc_hd__xor2_1 _5797_ (.A(_2443_),
    .B(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__mux2_1 _5798_ (.A0(net284),
    .A1(_2445_),
    .S(_1429_),
    .X(_2446_));
 sky130_fd_sc_hd__clkbuf_1 _5799_ (.A(_2446_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _5800_ (.A0(net26),
    .A1(\mix1.data_o[122] ),
    .S(_1338_),
    .X(_2447_));
 sky130_fd_sc_hd__mux2_1 _5801_ (.A0(\sub1.data_o[122] ),
    .A1(_2447_),
    .S(_1345_),
    .X(_2448_));
 sky130_fd_sc_hd__a32o_1 _5802_ (.A1(\mix1.data_o[122] ),
    .A2(_2325_),
    .A3(_1621_),
    .B1(_1355_),
    .B2(\sub1.data_o[122] ),
    .X(_2449_));
 sky130_fd_sc_hd__a22o_1 _5803_ (.A1(_1350_),
    .A2(_2448_),
    .B1(_2449_),
    .B2(_0678_),
    .X(_2450_));
 sky130_fd_sc_hd__mux2_2 _5804_ (.A0(\ks1.key_reg[122] ),
    .A1(net155),
    .S(_1625_),
    .X(_2451_));
 sky130_fd_sc_hd__xor2_1 _5805_ (.A(_2450_),
    .B(_2451_),
    .X(_2452_));
 sky130_fd_sc_hd__mux2_1 _5806_ (.A0(net285),
    .A1(_2452_),
    .S(_1429_),
    .X(_2453_));
 sky130_fd_sc_hd__clkbuf_1 _5807_ (.A(_2453_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _5808_ (.A0(net27),
    .A1(\mix1.data_o[123] ),
    .S(_1338_),
    .X(_2454_));
 sky130_fd_sc_hd__mux2_1 _5809_ (.A0(\sub1.data_o[123] ),
    .A1(_2454_),
    .S(_1345_),
    .X(_2455_));
 sky130_fd_sc_hd__a32o_1 _5810_ (.A1(\mix1.data_o[123] ),
    .A2(_2325_),
    .A3(_1621_),
    .B1(_1355_),
    .B2(\sub1.data_o[123] ),
    .X(_2456_));
 sky130_fd_sc_hd__a22o_1 _5811_ (.A1(_1350_),
    .A2(_2455_),
    .B1(_2456_),
    .B2(_0678_),
    .X(_2457_));
 sky130_fd_sc_hd__mux2_1 _5812_ (.A0(\ks1.key_reg[123] ),
    .A1(net156),
    .S(_1625_),
    .X(_2458_));
 sky130_fd_sc_hd__xor2_1 _5813_ (.A(_2457_),
    .B(_2458_),
    .X(_2459_));
 sky130_fd_sc_hd__mux2_1 _5814_ (.A0(net286),
    .A1(_2459_),
    .S(_1429_),
    .X(_2460_));
 sky130_fd_sc_hd__clkbuf_1 _5815_ (.A(_2460_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _5816_ (.A0(net28),
    .A1(\mix1.data_o[124] ),
    .S(_1338_),
    .X(_2461_));
 sky130_fd_sc_hd__mux2_1 _5817_ (.A0(\sub1.data_o[124] ),
    .A1(_2461_),
    .S(_1345_),
    .X(_2462_));
 sky130_fd_sc_hd__a32o_1 _5818_ (.A1(\mix1.data_o[124] ),
    .A2(_2325_),
    .A3(_1621_),
    .B1(_1355_),
    .B2(\sub1.data_o[124] ),
    .X(_2463_));
 sky130_fd_sc_hd__a22o_1 _5819_ (.A1(_1350_),
    .A2(_2462_),
    .B1(_2463_),
    .B2(_0678_),
    .X(_2464_));
 sky130_fd_sc_hd__mux2_1 _5820_ (.A0(\ks1.key_reg[124] ),
    .A1(net157),
    .S(_1625_),
    .X(_2465_));
 sky130_fd_sc_hd__xor2_1 _5821_ (.A(_2464_),
    .B(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__mux2_1 _5822_ (.A0(net287),
    .A1(_2466_),
    .S(_1429_),
    .X(_2467_));
 sky130_fd_sc_hd__clkbuf_1 _5823_ (.A(_2467_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _5824_ (.A0(net29),
    .A1(\mix1.data_o[125] ),
    .S(_1338_),
    .X(_2468_));
 sky130_fd_sc_hd__mux2_1 _5825_ (.A0(\sub1.data_o[125] ),
    .A1(_2468_),
    .S(_1345_),
    .X(_2469_));
 sky130_fd_sc_hd__a32o_1 _5826_ (.A1(\mix1.data_o[125] ),
    .A2(_2325_),
    .A3(_1621_),
    .B1(_1355_),
    .B2(\sub1.data_o[125] ),
    .X(_2470_));
 sky130_fd_sc_hd__a22o_1 _5827_ (.A1(_1350_),
    .A2(_2469_),
    .B1(_2470_),
    .B2(_0678_),
    .X(_2471_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(\ks1.key_reg[125] ),
    .A1(net158),
    .S(_1625_),
    .X(_2472_));
 sky130_fd_sc_hd__xor2_1 _5829_ (.A(_2471_),
    .B(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__mux2_1 _5830_ (.A0(net288),
    .A1(_2473_),
    .S(_1429_),
    .X(_2474_));
 sky130_fd_sc_hd__clkbuf_1 _5831_ (.A(_2474_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _5832_ (.A0(net30),
    .A1(\mix1.data_o[126] ),
    .S(_1338_),
    .X(_2475_));
 sky130_fd_sc_hd__mux2_1 _5833_ (.A0(\sub1.data_o[126] ),
    .A1(_2475_),
    .S(_1345_),
    .X(_2476_));
 sky130_fd_sc_hd__a32o_1 _5834_ (.A1(\mix1.data_o[126] ),
    .A2(_1306_),
    .A3(_1621_),
    .B1(_1355_),
    .B2(\sub1.data_o[126] ),
    .X(_2477_));
 sky130_fd_sc_hd__a22o_1 _5835_ (.A1(_1350_),
    .A2(_2476_),
    .B1(_2477_),
    .B2(_0678_),
    .X(_2478_));
 sky130_fd_sc_hd__mux2_1 _5836_ (.A0(\ks1.key_reg[126] ),
    .A1(net159),
    .S(_1625_),
    .X(_2479_));
 sky130_fd_sc_hd__xor2_1 _5837_ (.A(_2478_),
    .B(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__mux2_1 _5838_ (.A0(net289),
    .A1(_2480_),
    .S(_1429_),
    .X(_2481_));
 sky130_fd_sc_hd__clkbuf_1 _5839_ (.A(_2481_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _5840_ (.A0(net31),
    .A1(\mix1.data_o[127] ),
    .S(_1338_),
    .X(_2482_));
 sky130_fd_sc_hd__mux2_1 _5841_ (.A0(\sub1.data_o[127] ),
    .A1(_2482_),
    .S(_1345_),
    .X(_2483_));
 sky130_fd_sc_hd__a32o_1 _5842_ (.A1(\mix1.data_o[127] ),
    .A2(_1306_),
    .A3(_1621_),
    .B1(_1355_),
    .B2(\sub1.data_o[127] ),
    .X(_2484_));
 sky130_fd_sc_hd__a22o_1 _5843_ (.A1(_1350_),
    .A2(_2483_),
    .B1(_2484_),
    .B2(_0678_),
    .X(_2485_));
 sky130_fd_sc_hd__mux2_1 _5844_ (.A0(\ks1.key_reg[127] ),
    .A1(net160),
    .S(_1625_),
    .X(_2486_));
 sky130_fd_sc_hd__xor2_1 _5845_ (.A(_2485_),
    .B(_2486_),
    .X(_2487_));
 sky130_fd_sc_hd__mux2_1 _5846_ (.A0(net290),
    .A1(_2487_),
    .S(_1429_),
    .X(_2488_));
 sky130_fd_sc_hd__clkbuf_1 _5847_ (.A(_2488_),
    .X(_0143_));
 sky130_fd_sc_hd__clkbuf_4 _5848_ (.A(_0709_),
    .X(_2489_));
 sky130_fd_sc_hd__clkbuf_4 _5849_ (.A(_0662_),
    .X(_2490_));
 sky130_fd_sc_hd__buf_4 _5850_ (.A(_0662_),
    .X(_2491_));
 sky130_fd_sc_hd__nor2_2 _5851_ (.A(_2491_),
    .B(_2489_),
    .Y(_2492_));
 sky130_fd_sc_hd__a22o_1 _5852_ (.A1(\sub1.data_o[8] ),
    .A2(_2490_),
    .B1(_2492_),
    .B2(\sub1.data_o[72] ),
    .X(_2493_));
 sky130_fd_sc_hd__a31o_1 _5853_ (.A1(_1140_),
    .A2(_2489_),
    .A3(_1213_),
    .B1(_2493_),
    .X(_0144_));
 sky130_fd_sc_hd__a22o_1 _5854_ (.A1(\sub1.data_o[9] ),
    .A2(_2490_),
    .B1(_2492_),
    .B2(\sub1.data_o[73] ),
    .X(_2494_));
 sky130_fd_sc_hd__a31o_1 _5855_ (.A1(_1140_),
    .A2(_2489_),
    .A3(_1247_),
    .B1(_2494_),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_4 _5856_ (.A(_1139_),
    .X(_2495_));
 sky130_fd_sc_hd__a22o_1 _5857_ (.A1(\sub1.data_o[10] ),
    .A2(_2490_),
    .B1(_2492_),
    .B2(\sub1.data_o[74] ),
    .X(_2496_));
 sky130_fd_sc_hd__a31o_1 _5858_ (.A1(_2495_),
    .A2(_2489_),
    .A3(_1257_),
    .B1(_2496_),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_1 _5859_ (.A1(\sub1.data_o[11] ),
    .A2(_2490_),
    .B1(_2492_),
    .B2(\sub1.data_o[75] ),
    .X(_2497_));
 sky130_fd_sc_hd__a31o_1 _5860_ (.A1(_2495_),
    .A2(_2489_),
    .A3(_1272_),
    .B1(_2497_),
    .X(_0147_));
 sky130_fd_sc_hd__a22o_1 _5861_ (.A1(\sub1.data_o[12] ),
    .A2(_2490_),
    .B1(_2492_),
    .B2(\sub1.data_o[76] ),
    .X(_2498_));
 sky130_fd_sc_hd__a31o_1 _5862_ (.A1(_2495_),
    .A2(_2489_),
    .A3(_1278_),
    .B1(_2498_),
    .X(_0148_));
 sky130_fd_sc_hd__a22o_1 _5863_ (.A1(\sub1.data_o[13] ),
    .A2(_2490_),
    .B1(_2492_),
    .B2(\sub1.data_o[77] ),
    .X(_2499_));
 sky130_fd_sc_hd__a31o_1 _5864_ (.A1(_2495_),
    .A2(_2489_),
    .A3(_1286_),
    .B1(_2499_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_4 _5865_ (.A(_0662_),
    .X(_2500_));
 sky130_fd_sc_hd__a22o_1 _5866_ (.A1(\sub1.data_o[14] ),
    .A2(_2500_),
    .B1(_2492_),
    .B2(\sub1.data_o[78] ),
    .X(_2501_));
 sky130_fd_sc_hd__a31o_1 _5867_ (.A1(_2495_),
    .A2(_2489_),
    .A3(_1293_),
    .B1(_2501_),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_1 _5868_ (.A1(\sub1.data_o[15] ),
    .A2(_2500_),
    .B1(_2492_),
    .B2(\sub1.data_o[79] ),
    .X(_2502_));
 sky130_fd_sc_hd__a31o_1 _5869_ (.A1(_2495_),
    .A2(_2489_),
    .A3(_1300_),
    .B1(_2502_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _5870_ (.A0(\ks1.col[0] ),
    .A1(_1213_),
    .S(_0974_),
    .X(_2503_));
 sky130_fd_sc_hd__clkbuf_1 _5871_ (.A(_2503_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _5872_ (.A0(\ks1.col[1] ),
    .A1(_1247_),
    .S(_0974_),
    .X(_2504_));
 sky130_fd_sc_hd__clkbuf_1 _5873_ (.A(_2504_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _5874_ (.A0(\ks1.col[2] ),
    .A1(_1257_),
    .S(_0974_),
    .X(_2505_));
 sky130_fd_sc_hd__clkbuf_1 _5875_ (.A(_2505_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _5876_ (.A0(\ks1.col[3] ),
    .A1(_1270_),
    .S(_0974_),
    .X(_2506_));
 sky130_fd_sc_hd__clkbuf_1 _5877_ (.A(_2506_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _5878_ (.A0(\ks1.col[4] ),
    .A1(_1276_),
    .S(_0974_),
    .X(_2507_));
 sky130_fd_sc_hd__clkbuf_1 _5879_ (.A(_2507_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _5880_ (.A0(\ks1.col[5] ),
    .A1(_1282_),
    .S(_0974_),
    .X(_2508_));
 sky130_fd_sc_hd__clkbuf_1 _5881_ (.A(_2508_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(\ks1.col[6] ),
    .A1(_1293_),
    .S(_0974_),
    .X(_2509_));
 sky130_fd_sc_hd__clkbuf_1 _5883_ (.A(_2509_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _5884_ (.A0(\ks1.col[7] ),
    .A1(_1300_),
    .S(_0974_),
    .X(_2510_));
 sky130_fd_sc_hd__clkbuf_1 _5885_ (.A(_2510_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _5886_ (.A0(\ks1.col[24] ),
    .A1(_1212_),
    .S(_0850_),
    .X(_2511_));
 sky130_fd_sc_hd__clkbuf_1 _5887_ (.A(_2511_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _5888_ (.A0(net682),
    .A1(_1246_),
    .S(_0850_),
    .X(_2512_));
 sky130_fd_sc_hd__clkbuf_1 _5889_ (.A(_2512_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _5890_ (.A0(\ks1.col[26] ),
    .A1(_1256_),
    .S(_0850_),
    .X(_2513_));
 sky130_fd_sc_hd__clkbuf_1 _5891_ (.A(_2513_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _5892_ (.A0(net686),
    .A1(_1270_),
    .S(_0850_),
    .X(_2514_));
 sky130_fd_sc_hd__clkbuf_1 _5893_ (.A(_2514_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _5894_ (.A0(\ks1.col[28] ),
    .A1(_1278_),
    .S(_0850_),
    .X(_2515_));
 sky130_fd_sc_hd__clkbuf_1 _5895_ (.A(_2515_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _5896_ (.A0(\ks1.col[29] ),
    .A1(_1286_),
    .S(_0850_),
    .X(_2516_));
 sky130_fd_sc_hd__clkbuf_1 _5897_ (.A(_2516_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _5898_ (.A0(\ks1.col[30] ),
    .A1(_1292_),
    .S(_0850_),
    .X(_2517_));
 sky130_fd_sc_hd__clkbuf_1 _5899_ (.A(_2517_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _5900_ (.A0(\ks1.col[31] ),
    .A1(_1299_),
    .S(_0850_),
    .X(_2518_));
 sky130_fd_sc_hd__clkbuf_1 _5901_ (.A(_2518_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _5902_ (.A0(\ks1.col[16] ),
    .A1(_1212_),
    .S(_0649_),
    .X(_2519_));
 sky130_fd_sc_hd__clkbuf_1 _5903_ (.A(_2519_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _5904_ (.A0(net694),
    .A1(_1246_),
    .S(_0649_),
    .X(_2520_));
 sky130_fd_sc_hd__clkbuf_1 _5905_ (.A(_2520_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _5906_ (.A0(\ks1.col[18] ),
    .A1(_1256_),
    .S(_0649_),
    .X(_2521_));
 sky130_fd_sc_hd__clkbuf_1 _5907_ (.A(_2521_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _5908_ (.A0(\ks1.col[19] ),
    .A1(_1270_),
    .S(_0649_),
    .X(_2522_));
 sky130_fd_sc_hd__clkbuf_1 _5909_ (.A(_2522_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _5910_ (.A0(\ks1.col[20] ),
    .A1(_1277_),
    .S(_0649_),
    .X(_2523_));
 sky130_fd_sc_hd__clkbuf_1 _5911_ (.A(_2523_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _5912_ (.A0(\ks1.col[21] ),
    .A1(_1285_),
    .S(_0649_),
    .X(_2524_));
 sky130_fd_sc_hd__clkbuf_1 _5913_ (.A(_2524_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _5914_ (.A0(\ks1.col[22] ),
    .A1(_1292_),
    .S(_0649_),
    .X(_2525_));
 sky130_fd_sc_hd__clkbuf_1 _5915_ (.A(_2525_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _5916_ (.A0(\ks1.col[23] ),
    .A1(_1299_),
    .S(_0649_),
    .X(_2526_));
 sky130_fd_sc_hd__clkbuf_1 _5917_ (.A(_2526_),
    .X(_0175_));
 sky130_fd_sc_hd__a22oi_4 _5918_ (.A1(_0682_),
    .A2(\sub1.ready_o ),
    .B1(addroundkey_ready_o),
    .B2(_0738_),
    .Y(_2527_));
 sky130_fd_sc_hd__a2111oi_4 _5919_ (.A1(state),
    .A2(_1127_),
    .B1(_2527_),
    .C1(\mix1.state[1] ),
    .D1(\mix1.state[0] ),
    .Y(_2528_));
 sky130_fd_sc_hd__clkbuf_4 _5920_ (.A(_2528_),
    .X(_2529_));
 sky130_fd_sc_hd__clkbuf_8 _5921_ (.A(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__clkbuf_4 _5922_ (.A(_2530_),
    .X(_2531_));
 sky130_fd_sc_hd__nor2b_2 _5923_ (.A(\mix1.state[1] ),
    .B_N(\mix1.state[0] ),
    .Y(_2532_));
 sky130_fd_sc_hd__buf_4 _5924_ (.A(_2532_),
    .X(_2533_));
 sky130_fd_sc_hd__clkbuf_4 _5925_ (.A(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__clkbuf_4 _5926_ (.A(_2534_),
    .X(_2535_));
 sky130_fd_sc_hd__buf_4 _5927_ (.A(_2535_),
    .X(_2536_));
 sky130_fd_sc_hd__buf_4 _5928_ (.A(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__clkbuf_4 _5929_ (.A(_0652_),
    .X(_2538_));
 sky130_fd_sc_hd__nor2b_2 _5930_ (.A(\mix1.state[0] ),
    .B_N(\mix1.state[1] ),
    .Y(_2539_));
 sky130_fd_sc_hd__buf_4 _5931_ (.A(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__clkbuf_4 _5932_ (.A(_2540_),
    .X(_2541_));
 sky130_fd_sc_hd__clkbuf_4 _5933_ (.A(_2541_),
    .X(_2542_));
 sky130_fd_sc_hd__buf_4 _5934_ (.A(_2542_),
    .X(_2543_));
 sky130_fd_sc_hd__a22o_1 _5935_ (.A1(\sub1.data_o[16] ),
    .A2(_2538_),
    .B1(_2543_),
    .B2(\sub1.data_o[48] ),
    .X(_2544_));
 sky130_fd_sc_hd__clkbuf_4 _5936_ (.A(_0807_),
    .X(_2545_));
 sky130_fd_sc_hd__clkbuf_4 _5937_ (.A(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__buf_4 _5938_ (.A(_2546_),
    .X(_2547_));
 sky130_fd_sc_hd__a211o_1 _5939_ (.A1(\sub1.data_o[80] ),
    .A2(_2537_),
    .B1(_2544_),
    .C1(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__a21oi_1 _5940_ (.A1(\sub1.data_o[112] ),
    .A2(_2531_),
    .B1(_2548_),
    .Y(_2549_));
 sky130_fd_sc_hd__a22o_1 _5941_ (.A1(net295),
    .A2(_2538_),
    .B1(_2543_),
    .B2(net330),
    .X(_2550_));
 sky130_fd_sc_hd__a211o_1 _5942_ (.A1(net366),
    .A2(_2537_),
    .B1(_2550_),
    .C1(_1343_),
    .X(_2551_));
 sky130_fd_sc_hd__a21oi_1 _5943_ (.A1(net274),
    .A2(_2531_),
    .B1(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__nor2_4 _5944_ (.A(_2549_),
    .B(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__a22o_1 _5945_ (.A1(\sub1.data_o[88] ),
    .A2(_2536_),
    .B1(_2543_),
    .B2(\sub1.data_o[56] ),
    .X(_2554_));
 sky130_fd_sc_hd__a211o_1 _5946_ (.A1(\sub1.data_o[24] ),
    .A2(_0653_),
    .B1(_2546_),
    .C1(_2554_),
    .X(_2555_));
 sky130_fd_sc_hd__a21oi_1 _5947_ (.A1(\sub1.data_o[120] ),
    .A2(_2531_),
    .B1(_2555_),
    .Y(_2556_));
 sky130_fd_sc_hd__a22o_1 _5948_ (.A1(net374),
    .A2(_2536_),
    .B1(_2543_),
    .B2(net339),
    .X(_2557_));
 sky130_fd_sc_hd__a211o_1 _5949_ (.A1(net304),
    .A2(_0653_),
    .B1(_1342_),
    .C1(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__a21oi_1 _5950_ (.A1(net283),
    .A2(_2531_),
    .B1(_2558_),
    .Y(_2559_));
 sky130_fd_sc_hd__nor2_4 _5951_ (.A(_2556_),
    .B(_2559_),
    .Y(_2560_));
 sky130_fd_sc_hd__xor2_4 _5952_ (.A(_2553_),
    .B(_2560_),
    .X(_2561_));
 sky130_fd_sc_hd__a22o_1 _5953_ (.A1(\sub1.data_o[77] ),
    .A2(_2535_),
    .B1(_2542_),
    .B2(\sub1.data_o[45] ),
    .X(_2562_));
 sky130_fd_sc_hd__a211o_1 _5954_ (.A1(\sub1.data_o[13] ),
    .A2(_0652_),
    .B1(_2546_),
    .C1(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__a21oi_2 _5955_ (.A1(\sub1.data_o[109] ),
    .A2(_2530_),
    .B1(_2563_),
    .Y(_2564_));
 sky130_fd_sc_hd__a22o_1 _5956_ (.A1(net362),
    .A2(_2535_),
    .B1(_2542_),
    .B2(net327),
    .X(_2565_));
 sky130_fd_sc_hd__a211o_1 _5957_ (.A1(net292),
    .A2(_0652_),
    .B1(_1341_),
    .C1(_2565_),
    .X(_2566_));
 sky130_fd_sc_hd__a21oi_2 _5958_ (.A1(net270),
    .A2(_2530_),
    .B1(_2566_),
    .Y(_2567_));
 sky130_fd_sc_hd__nor2_8 _5959_ (.A(_2564_),
    .B(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__a22o_1 _5960_ (.A1(\sub1.data_o[70] ),
    .A2(_2533_),
    .B1(_2540_),
    .B2(\sub1.data_o[38] ),
    .X(_2569_));
 sky130_fd_sc_hd__a211o_1 _5961_ (.A1(\sub1.data_o[6] ),
    .A2(_0651_),
    .B1(_2545_),
    .C1(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__a21o_1 _5962_ (.A1(\sub1.data_o[102] ),
    .A2(_2529_),
    .B1(_2570_),
    .X(_2571_));
 sky130_fd_sc_hd__a22o_1 _5963_ (.A1(net355),
    .A2(_2533_),
    .B1(_2540_),
    .B2(net319),
    .X(_2572_));
 sky130_fd_sc_hd__a211o_1 _5964_ (.A1(net354),
    .A2(_0651_),
    .B1(_0798_),
    .C1(_2572_),
    .X(_2573_));
 sky130_fd_sc_hd__a21o_1 _5965_ (.A1(net263),
    .A2(_2529_),
    .B1(_2573_),
    .X(_2574_));
 sky130_fd_sc_hd__nand2_8 _5966_ (.A(_2571_),
    .B(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__buf_4 _5967_ (.A(_2529_),
    .X(_2576_));
 sky130_fd_sc_hd__clkbuf_4 _5968_ (.A(_0651_),
    .X(_2577_));
 sky130_fd_sc_hd__a22o_1 _5969_ (.A1(\sub1.data_o[85] ),
    .A2(_2534_),
    .B1(_2541_),
    .B2(\sub1.data_o[53] ),
    .X(_2578_));
 sky130_fd_sc_hd__a211o_1 _5970_ (.A1(\sub1.data_o[21] ),
    .A2(_2577_),
    .B1(_2545_),
    .C1(_2578_),
    .X(_2579_));
 sky130_fd_sc_hd__a21oi_2 _5971_ (.A1(\sub1.data_o[117] ),
    .A2(_2576_),
    .B1(_2579_),
    .Y(_2580_));
 sky130_fd_sc_hd__a22o_1 _5972_ (.A1(net371),
    .A2(_2534_),
    .B1(_2541_),
    .B2(net336),
    .X(_2581_));
 sky130_fd_sc_hd__a211o_1 _5973_ (.A1(net301),
    .A2(_2577_),
    .B1(_1341_),
    .C1(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__a21oi_2 _5974_ (.A1(net279),
    .A2(_2576_),
    .B1(_2582_),
    .Y(_2583_));
 sky130_fd_sc_hd__nor2_8 _5975_ (.A(_2580_),
    .B(_2583_),
    .Y(_2584_));
 sky130_fd_sc_hd__xnor2_2 _5976_ (.A(_2575_),
    .B(_2584_),
    .Y(_2585_));
 sky130_fd_sc_hd__xnor2_4 _5977_ (.A(_2568_),
    .B(_2585_),
    .Y(_2586_));
 sky130_fd_sc_hd__a22o_1 _5978_ (.A1(\sub1.data_o[86] ),
    .A2(_2533_),
    .B1(_2540_),
    .B2(\sub1.data_o[54] ),
    .X(_2587_));
 sky130_fd_sc_hd__a211o_1 _5979_ (.A1(\sub1.data_o[22] ),
    .A2(_2577_),
    .B1(_2545_),
    .C1(_2587_),
    .X(_2588_));
 sky130_fd_sc_hd__a21o_1 _5980_ (.A1(\sub1.data_o[118] ),
    .A2(_2529_),
    .B1(_2588_),
    .X(_2589_));
 sky130_fd_sc_hd__a22o_1 _5981_ (.A1(net372),
    .A2(_2533_),
    .B1(_2540_),
    .B2(net337),
    .X(_2590_));
 sky130_fd_sc_hd__a211o_1 _5982_ (.A1(net302),
    .A2(_0651_),
    .B1(_0798_),
    .C1(_2590_),
    .X(_2591_));
 sky130_fd_sc_hd__a21o_1 _5983_ (.A1(net280),
    .A2(_2529_),
    .B1(_2591_),
    .X(_2592_));
 sky130_fd_sc_hd__nand2_8 _5984_ (.A(_2589_),
    .B(_2592_),
    .Y(_2593_));
 sky130_fd_sc_hd__a22o_1 _5985_ (.A1(\sub1.data_o[69] ),
    .A2(_2533_),
    .B1(_2540_),
    .B2(\sub1.data_o[37] ),
    .X(_2594_));
 sky130_fd_sc_hd__a211o_1 _5986_ (.A1(\sub1.data_o[5] ),
    .A2(_2577_),
    .B1(_2545_),
    .C1(_2594_),
    .X(_2595_));
 sky130_fd_sc_hd__a21oi_1 _5987_ (.A1(\sub1.data_o[101] ),
    .A2(_2529_),
    .B1(_2595_),
    .Y(_2596_));
 sky130_fd_sc_hd__a22o_1 _5988_ (.A1(net353),
    .A2(_2533_),
    .B1(_2540_),
    .B2(net318),
    .X(_2597_));
 sky130_fd_sc_hd__a211o_1 _5989_ (.A1(net343),
    .A2(_2577_),
    .B1(_1341_),
    .C1(_2597_),
    .X(_2598_));
 sky130_fd_sc_hd__a21oi_2 _5990_ (.A1(net262),
    .A2(_2576_),
    .B1(_2598_),
    .Y(_2599_));
 sky130_fd_sc_hd__nor2_4 _5991_ (.A(_2596_),
    .B(_2599_),
    .Y(_2600_));
 sky130_fd_sc_hd__a22o_1 _5992_ (.A1(\sub1.data_o[93] ),
    .A2(_2533_),
    .B1(_2540_),
    .B2(\sub1.data_o[61] ),
    .X(_2601_));
 sky130_fd_sc_hd__a211o_1 _5993_ (.A1(\sub1.data_o[29] ),
    .A2(_2577_),
    .B1(_2545_),
    .C1(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__a21oi_2 _5994_ (.A1(\sub1.data_o[125] ),
    .A2(_2576_),
    .B1(_2602_),
    .Y(_2603_));
 sky130_fd_sc_hd__a22o_1 _5995_ (.A1(net380),
    .A2(_2534_),
    .B1(_2541_),
    .B2(net345),
    .X(_2604_));
 sky130_fd_sc_hd__a211o_1 _5996_ (.A1(net309),
    .A2(_2577_),
    .B1(_1341_),
    .C1(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__a21oi_2 _5997_ (.A1(net288),
    .A2(_2576_),
    .B1(_2605_),
    .Y(_2606_));
 sky130_fd_sc_hd__nor2_8 _5998_ (.A(_2603_),
    .B(_2606_),
    .Y(_2607_));
 sky130_fd_sc_hd__xnor2_4 _5999_ (.A(_2600_),
    .B(_2607_),
    .Y(_2608_));
 sky130_fd_sc_hd__xnor2_4 _6000_ (.A(_2593_),
    .B(_2608_),
    .Y(_2609_));
 sky130_fd_sc_hd__xnor2_2 _6001_ (.A(_2586_),
    .B(_2609_),
    .Y(_2610_));
 sky130_fd_sc_hd__or2_1 _6002_ (.A(_0682_),
    .B(_2610_),
    .X(_2611_));
 sky130_fd_sc_hd__clkbuf_4 _6003_ (.A(_2531_),
    .X(_2612_));
 sky130_fd_sc_hd__buf_4 _6004_ (.A(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__buf_4 _6005_ (.A(_2537_),
    .X(_2614_));
 sky130_fd_sc_hd__buf_4 _6006_ (.A(_2543_),
    .X(_2615_));
 sky130_fd_sc_hd__buf_4 _6007_ (.A(_2615_),
    .X(_2616_));
 sky130_fd_sc_hd__a22o_1 _6008_ (.A1(\sub1.data_o[72] ),
    .A2(_2614_),
    .B1(_2616_),
    .B2(\sub1.data_o[40] ),
    .X(_2617_));
 sky130_fd_sc_hd__a211o_1 _6009_ (.A1(\sub1.data_o[8] ),
    .A2(_0654_),
    .B1(_2547_),
    .C1(_2617_),
    .X(_2618_));
 sky130_fd_sc_hd__a21oi_1 _6010_ (.A1(\sub1.data_o[104] ),
    .A2(_2613_),
    .B1(_2618_),
    .Y(_2619_));
 sky130_fd_sc_hd__a22o_1 _6011_ (.A1(net357),
    .A2(_2614_),
    .B1(_2616_),
    .B2(net322),
    .X(_2620_));
 sky130_fd_sc_hd__a211o_1 _6012_ (.A1(net376),
    .A2(_0654_),
    .B1(_1343_),
    .C1(_2620_),
    .X(_2621_));
 sky130_fd_sc_hd__a21oi_1 _6013_ (.A1(net265),
    .A2(_2613_),
    .B1(_2621_),
    .Y(_2622_));
 sky130_fd_sc_hd__nor2_4 _6014_ (.A(_2619_),
    .B(_2622_),
    .Y(_2623_));
 sky130_fd_sc_hd__xnor2_2 _6015_ (.A(_2611_),
    .B(_2623_),
    .Y(_2624_));
 sky130_fd_sc_hd__a22o_1 _6016_ (.A1(\sub1.data_o[71] ),
    .A2(_2532_),
    .B1(_2539_),
    .B2(\sub1.data_o[39] ),
    .X(_2625_));
 sky130_fd_sc_hd__a211o_1 _6017_ (.A1(\sub1.data_o[7] ),
    .A2(_0650_),
    .B1(_0807_),
    .C1(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__a21o_1 _6018_ (.A1(\sub1.data_o[103] ),
    .A2(_2528_),
    .B1(_2626_),
    .X(_2627_));
 sky130_fd_sc_hd__a22o_1 _6019_ (.A1(net356),
    .A2(_2532_),
    .B1(_2539_),
    .B2(net320),
    .X(_2628_));
 sky130_fd_sc_hd__a211o_1 _6020_ (.A1(net365),
    .A2(_0650_),
    .B1(_0798_),
    .C1(_2628_),
    .X(_2629_));
 sky130_fd_sc_hd__a21o_1 _6021_ (.A1(net264),
    .A2(_2528_),
    .B1(_2629_),
    .X(_2630_));
 sky130_fd_sc_hd__nand2_8 _6022_ (.A(_2627_),
    .B(_2630_),
    .Y(_2631_));
 sky130_fd_sc_hd__a22o_1 _6023_ (.A1(\sub1.data_o[95] ),
    .A2(_2532_),
    .B1(_2539_),
    .B2(\sub1.data_o[63] ),
    .X(_2632_));
 sky130_fd_sc_hd__a211o_1 _6024_ (.A1(\sub1.data_o[31] ),
    .A2(_0650_),
    .B1(_0807_),
    .C1(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__a21oi_2 _6025_ (.A1(\sub1.data_o[127] ),
    .A2(_2528_),
    .B1(_2633_),
    .Y(_2634_));
 sky130_fd_sc_hd__a22o_1 _6026_ (.A1(net382),
    .A2(_2532_),
    .B1(_2539_),
    .B2(net347),
    .X(_2635_));
 sky130_fd_sc_hd__a211o_1 _6027_ (.A1(net312),
    .A2(_0651_),
    .B1(_0798_),
    .C1(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__a21oi_2 _6028_ (.A1(net290),
    .A2(_2528_),
    .B1(_2636_),
    .Y(_2637_));
 sky130_fd_sc_hd__nor2_8 _6029_ (.A(_2634_),
    .B(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__xor2_4 _6030_ (.A(_2631_),
    .B(_2638_),
    .X(_2639_));
 sky130_fd_sc_hd__xor2_2 _6031_ (.A(_2624_),
    .B(_2639_),
    .X(_2640_));
 sky130_fd_sc_hd__xnor2_4 _6032_ (.A(_2561_),
    .B(_2640_),
    .Y(_2641_));
 sky130_fd_sc_hd__clkbuf_4 _6033_ (.A(_2614_),
    .X(_2642_));
 sky130_fd_sc_hd__mux2_1 _6034_ (.A0(net568),
    .A1(_2641_),
    .S(_2642_),
    .X(_2643_));
 sky130_fd_sc_hd__clkbuf_1 _6035_ (.A(_2643_),
    .X(_0176_));
 sky130_fd_sc_hd__a22o_1 _6036_ (.A1(\sub1.data_o[94] ),
    .A2(_2535_),
    .B1(_2542_),
    .B2(\sub1.data_o[62] ),
    .X(_2644_));
 sky130_fd_sc_hd__a211o_1 _6037_ (.A1(\sub1.data_o[30] ),
    .A2(_2538_),
    .B1(_2546_),
    .C1(_2644_),
    .X(_2645_));
 sky130_fd_sc_hd__a21oi_4 _6038_ (.A1(\sub1.data_o[126] ),
    .A2(_2530_),
    .B1(_2645_),
    .Y(_2646_));
 sky130_fd_sc_hd__clkbuf_4 _6039_ (.A(_2576_),
    .X(_2647_));
 sky130_fd_sc_hd__a22o_2 _6040_ (.A1(net381),
    .A2(_2535_),
    .B1(_2542_),
    .B2(net346),
    .X(_2648_));
 sky130_fd_sc_hd__a211o_1 _6041_ (.A1(net311),
    .A2(_2538_),
    .B1(_1342_),
    .C1(_2648_),
    .X(_2649_));
 sky130_fd_sc_hd__a21oi_2 _6042_ (.A1(net289),
    .A2(_2647_),
    .B1(_2649_),
    .Y(_2650_));
 sky130_fd_sc_hd__nor2_8 _6043_ (.A(_2646_),
    .B(_2650_),
    .Y(_2651_));
 sky130_fd_sc_hd__xnor2_4 _6044_ (.A(_2575_),
    .B(_2651_),
    .Y(_2652_));
 sky130_fd_sc_hd__a22o_1 _6045_ (.A1(\sub1.data_o[87] ),
    .A2(_2534_),
    .B1(_2541_),
    .B2(\sub1.data_o[55] ),
    .X(_2653_));
 sky130_fd_sc_hd__a211o_1 _6046_ (.A1(\sub1.data_o[23] ),
    .A2(_2577_),
    .B1(_2545_),
    .C1(_2653_),
    .X(_2654_));
 sky130_fd_sc_hd__a21oi_2 _6047_ (.A1(\sub1.data_o[119] ),
    .A2(_2576_),
    .B1(_2654_),
    .Y(_2655_));
 sky130_fd_sc_hd__a22o_1 _6048_ (.A1(net373),
    .A2(_2534_),
    .B1(_2541_),
    .B2(net338),
    .X(_2656_));
 sky130_fd_sc_hd__a211o_1 _6049_ (.A1(net303),
    .A2(_2577_),
    .B1(_1341_),
    .C1(_2656_),
    .X(_2657_));
 sky130_fd_sc_hd__a21oi_2 _6050_ (.A1(net281),
    .A2(_2576_),
    .B1(_2657_),
    .Y(_2658_));
 sky130_fd_sc_hd__nor2_8 _6051_ (.A(_2655_),
    .B(_2658_),
    .Y(_2659_));
 sky130_fd_sc_hd__xor2_2 _6052_ (.A(_2631_),
    .B(_2659_),
    .X(_2660_));
 sky130_fd_sc_hd__a22o_1 _6053_ (.A1(\sub1.data_o[78] ),
    .A2(_2534_),
    .B1(_2541_),
    .B2(\sub1.data_o[46] ),
    .X(_2661_));
 sky130_fd_sc_hd__a211o_1 _6054_ (.A1(\sub1.data_o[14] ),
    .A2(_2577_),
    .B1(_2545_),
    .C1(_2661_),
    .X(_2662_));
 sky130_fd_sc_hd__a21oi_2 _6055_ (.A1(\sub1.data_o[110] ),
    .A2(_2576_),
    .B1(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__a22o_1 _6056_ (.A1(net363),
    .A2(_2534_),
    .B1(_2541_),
    .B2(net328),
    .X(_2664_));
 sky130_fd_sc_hd__a211o_1 _6057_ (.A1(net293),
    .A2(_0652_),
    .B1(_1341_),
    .C1(_2664_),
    .X(_2665_));
 sky130_fd_sc_hd__a21oi_2 _6058_ (.A1(net272),
    .A2(_2576_),
    .B1(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__nor2_8 _6059_ (.A(_2663_),
    .B(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__xnor2_2 _6060_ (.A(_2593_),
    .B(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__xnor2_2 _6061_ (.A(_2660_),
    .B(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__xor2_4 _6062_ (.A(_2652_),
    .B(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__xnor2_1 _6063_ (.A(_2610_),
    .B(_2670_),
    .Y(_2671_));
 sky130_fd_sc_hd__nand2_2 _6064_ (.A(_1218_),
    .B(_2671_),
    .Y(_2672_));
 sky130_fd_sc_hd__a22o_1 _6065_ (.A1(\sub1.data_o[89] ),
    .A2(_2535_),
    .B1(_2542_),
    .B2(\sub1.data_o[57] ),
    .X(_2673_));
 sky130_fd_sc_hd__a211o_1 _6066_ (.A1(\sub1.data_o[25] ),
    .A2(_2538_),
    .B1(_2546_),
    .C1(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__a21oi_2 _6067_ (.A1(\sub1.data_o[121] ),
    .A2(_2530_),
    .B1(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__a22o_1 _6068_ (.A1(net375),
    .A2(_2535_),
    .B1(_2542_),
    .B2(net340),
    .X(_2676_));
 sky130_fd_sc_hd__a211o_1 _6069_ (.A1(net305),
    .A2(_0652_),
    .B1(_1341_),
    .C1(_2676_),
    .X(_2677_));
 sky130_fd_sc_hd__a21oi_2 _6070_ (.A1(net284),
    .A2(_2530_),
    .B1(_2677_),
    .Y(_2678_));
 sky130_fd_sc_hd__nor2_8 _6071_ (.A(_2675_),
    .B(_2678_),
    .Y(_2679_));
 sky130_fd_sc_hd__buf_4 _6072_ (.A(_0653_),
    .X(_2680_));
 sky130_fd_sc_hd__a22o_1 _6073_ (.A1(\sub1.data_o[64] ),
    .A2(_2536_),
    .B1(_2543_),
    .B2(\sub1.data_o[32] ),
    .X(_2681_));
 sky130_fd_sc_hd__a211o_1 _6074_ (.A1(\sub1.data_o[0] ),
    .A2(_2680_),
    .B1(_2547_),
    .C1(_2681_),
    .X(_2682_));
 sky130_fd_sc_hd__a21oi_1 _6075_ (.A1(\sub1.data_o[96] ),
    .A2(_2531_),
    .B1(_2682_),
    .Y(_2683_));
 sky130_fd_sc_hd__a22o_1 _6076_ (.A1(net348),
    .A2(_2536_),
    .B1(_2543_),
    .B2(net313),
    .X(_2684_));
 sky130_fd_sc_hd__a211o_1 _6077_ (.A1(net260),
    .A2(_0653_),
    .B1(_1342_),
    .C1(_2684_),
    .X(_2685_));
 sky130_fd_sc_hd__a21oi_1 _6078_ (.A1(net383),
    .A2(_2531_),
    .B1(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__nor2_4 _6079_ (.A(_2683_),
    .B(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hd__xor2_2 _6080_ (.A(_2639_),
    .B(_2687_),
    .X(_2688_));
 sky130_fd_sc_hd__xnor2_2 _6081_ (.A(_2560_),
    .B(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__xnor2_1 _6082_ (.A(_2679_),
    .B(_2689_),
    .Y(_2690_));
 sky130_fd_sc_hd__xnor2_2 _6083_ (.A(_2672_),
    .B(_2690_),
    .Y(_2691_));
 sky130_fd_sc_hd__a22o_1 _6084_ (.A1(\sub1.data_o[73] ),
    .A2(_2535_),
    .B1(_2542_),
    .B2(\sub1.data_o[41] ),
    .X(_2692_));
 sky130_fd_sc_hd__a211o_1 _6085_ (.A1(\sub1.data_o[9] ),
    .A2(_0652_),
    .B1(_2545_),
    .C1(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__a21o_1 _6086_ (.A1(\sub1.data_o[105] ),
    .A2(_2530_),
    .B1(_2693_),
    .X(_2694_));
 sky130_fd_sc_hd__a22o_1 _6087_ (.A1(net358),
    .A2(_2535_),
    .B1(_2542_),
    .B2(net323),
    .X(_2695_));
 sky130_fd_sc_hd__a211o_1 _6088_ (.A1(net387),
    .A2(_0652_),
    .B1(_1341_),
    .C1(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__a21o_1 _6089_ (.A1(net266),
    .A2(_2530_),
    .B1(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__nand2_8 _6090_ (.A(_2694_),
    .B(_2697_),
    .Y(_2698_));
 sky130_fd_sc_hd__clkbuf_4 _6091_ (.A(_2534_),
    .X(_2699_));
 sky130_fd_sc_hd__clkbuf_4 _6092_ (.A(_2541_),
    .X(_2700_));
 sky130_fd_sc_hd__a22o_1 _6093_ (.A1(\sub1.data_o[81] ),
    .A2(_2699_),
    .B1(_2700_),
    .B2(\sub1.data_o[49] ),
    .X(_2701_));
 sky130_fd_sc_hd__a211o_1 _6094_ (.A1(\sub1.data_o[17] ),
    .A2(_2538_),
    .B1(_2546_),
    .C1(_2701_),
    .X(_2702_));
 sky130_fd_sc_hd__a21oi_1 _6095_ (.A1(\sub1.data_o[113] ),
    .A2(_2647_),
    .B1(_2702_),
    .Y(_2703_));
 sky130_fd_sc_hd__a22o_1 _6096_ (.A1(net367),
    .A2(_2699_),
    .B1(_2700_),
    .B2(net331),
    .X(_2704_));
 sky130_fd_sc_hd__a211o_1 _6097_ (.A1(net296),
    .A2(_2538_),
    .B1(_1342_),
    .C1(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__a21oi_1 _6098_ (.A1(net275),
    .A2(_2647_),
    .B1(_2705_),
    .Y(_2706_));
 sky130_fd_sc_hd__nor2_4 _6099_ (.A(_2703_),
    .B(_2706_),
    .Y(_2707_));
 sky130_fd_sc_hd__xnor2_4 _6100_ (.A(_2698_),
    .B(_2707_),
    .Y(_2708_));
 sky130_fd_sc_hd__xnor2_4 _6101_ (.A(_2691_),
    .B(_2708_),
    .Y(_2709_));
 sky130_fd_sc_hd__mux2_1 _6102_ (.A0(net584),
    .A1(_2709_),
    .S(_2642_),
    .X(_2710_));
 sky130_fd_sc_hd__clkbuf_1 _6103_ (.A(_2710_),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_1 _6104_ (.A1(\sub1.data_o[79] ),
    .A2(_2535_),
    .B1(_2542_),
    .B2(\sub1.data_o[47] ),
    .X(_2711_));
 sky130_fd_sc_hd__a211o_1 _6105_ (.A1(\sub1.data_o[15] ),
    .A2(_0652_),
    .B1(_2545_),
    .C1(_2711_),
    .X(_2712_));
 sky130_fd_sc_hd__a21oi_4 _6106_ (.A1(\sub1.data_o[111] ),
    .A2(_2530_),
    .B1(_2712_),
    .Y(_2713_));
 sky130_fd_sc_hd__a22o_1 _6107_ (.A1(net364),
    .A2(_2534_),
    .B1(_2541_),
    .B2(net329),
    .X(_2714_));
 sky130_fd_sc_hd__a211o_1 _6108_ (.A1(net294),
    .A2(_0652_),
    .B1(_1341_),
    .C1(_2714_),
    .X(_2715_));
 sky130_fd_sc_hd__a21oi_2 _6109_ (.A1(net273),
    .A2(_2530_),
    .B1(_2715_),
    .Y(_2716_));
 sky130_fd_sc_hd__nor2_8 _6110_ (.A(_2713_),
    .B(_2716_),
    .Y(_2717_));
 sky130_fd_sc_hd__xnor2_4 _6111_ (.A(_2659_),
    .B(_2717_),
    .Y(_2718_));
 sky130_fd_sc_hd__xor2_2 _6112_ (.A(_2553_),
    .B(_2718_),
    .X(_2719_));
 sky130_fd_sc_hd__xor2_1 _6113_ (.A(_2688_),
    .B(_2719_),
    .X(_2720_));
 sky130_fd_sc_hd__o21ai_1 _6114_ (.A1(_2670_),
    .A2(_2720_),
    .B1(_1217_),
    .Y(_2721_));
 sky130_fd_sc_hd__a21o_1 _6115_ (.A1(_2670_),
    .A2(_2720_),
    .B1(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__a22o_1 _6116_ (.A1(\sub1.data_o[74] ),
    .A2(_2699_),
    .B1(_2700_),
    .B2(\sub1.data_o[42] ),
    .X(_2723_));
 sky130_fd_sc_hd__a211o_1 _6117_ (.A1(\sub1.data_o[10] ),
    .A2(_2538_),
    .B1(_2546_),
    .C1(_2723_),
    .X(_2724_));
 sky130_fd_sc_hd__a21o_1 _6118_ (.A1(\sub1.data_o[106] ),
    .A2(_2647_),
    .B1(_2724_),
    .X(_2725_));
 sky130_fd_sc_hd__a22o_1 _6119_ (.A1(net359),
    .A2(_2699_),
    .B1(_2700_),
    .B2(net324),
    .X(_2726_));
 sky130_fd_sc_hd__a211o_1 _6120_ (.A1(net271),
    .A2(_2538_),
    .B1(_1342_),
    .C1(_2726_),
    .X(_2727_));
 sky130_fd_sc_hd__a21o_1 _6121_ (.A1(net267),
    .A2(_2647_),
    .B1(_2727_),
    .X(_2728_));
 sky130_fd_sc_hd__nand2_4 _6122_ (.A(_2725_),
    .B(_2728_),
    .Y(_2729_));
 sky130_fd_sc_hd__a22o_1 _6123_ (.A1(\sub1.data_o[90] ),
    .A2(_2532_),
    .B1(_2539_),
    .B2(\sub1.data_o[58] ),
    .X(_2730_));
 sky130_fd_sc_hd__a211o_1 _6124_ (.A1(\sub1.data_o[26] ),
    .A2(_0651_),
    .B1(_0807_),
    .C1(_2730_),
    .X(_2731_));
 sky130_fd_sc_hd__a21o_1 _6125_ (.A1(\sub1.data_o[122] ),
    .A2(_2529_),
    .B1(_2731_),
    .X(_2732_));
 sky130_fd_sc_hd__a22o_1 _6126_ (.A1(net377),
    .A2(_2532_),
    .B1(_2539_),
    .B2(net341),
    .X(_2733_));
 sky130_fd_sc_hd__a211o_1 _6127_ (.A1(net306),
    .A2(_0651_),
    .B1(_0798_),
    .C1(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__a21o_1 _6128_ (.A1(net285),
    .A2(_2528_),
    .B1(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__nand2_4 _6129_ (.A(_2732_),
    .B(_2735_),
    .Y(_2736_));
 sky130_fd_sc_hd__xor2_4 _6130_ (.A(_2729_),
    .B(_2736_),
    .X(_2737_));
 sky130_fd_sc_hd__xnor2_4 _6131_ (.A(_2722_),
    .B(_2737_),
    .Y(_2738_));
 sky130_fd_sc_hd__a22o_1 _6132_ (.A1(\sub1.data_o[82] ),
    .A2(_2699_),
    .B1(_2700_),
    .B2(\sub1.data_o[50] ),
    .X(_2739_));
 sky130_fd_sc_hd__a211o_1 _6133_ (.A1(\sub1.data_o[18] ),
    .A2(_0653_),
    .B1(_2546_),
    .C1(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__a21oi_1 _6134_ (.A1(\sub1.data_o[114] ),
    .A2(_2647_),
    .B1(_2740_),
    .Y(_2741_));
 sky130_fd_sc_hd__a22o_1 _6135_ (.A1(net368),
    .A2(_2699_),
    .B1(_2700_),
    .B2(net333),
    .X(_2742_));
 sky130_fd_sc_hd__a211o_1 _6136_ (.A1(net297),
    .A2(_0653_),
    .B1(_1342_),
    .C1(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__a21oi_1 _6137_ (.A1(net276),
    .A2(_2531_),
    .B1(_2743_),
    .Y(_2744_));
 sky130_fd_sc_hd__nor2_4 _6138_ (.A(_2741_),
    .B(_2744_),
    .Y(_2745_));
 sky130_fd_sc_hd__a22o_1 _6139_ (.A1(\sub1.data_o[65] ),
    .A2(_2699_),
    .B1(_2700_),
    .B2(\sub1.data_o[33] ),
    .X(_2746_));
 sky130_fd_sc_hd__a211o_1 _6140_ (.A1(\sub1.data_o[1] ),
    .A2(_2538_),
    .B1(_2546_),
    .C1(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__a21oi_1 _6141_ (.A1(\sub1.data_o[97] ),
    .A2(_2647_),
    .B1(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__a22o_1 _6142_ (.A1(net349),
    .A2(_2699_),
    .B1(_2700_),
    .B2(net314),
    .X(_2749_));
 sky130_fd_sc_hd__a211o_1 _6143_ (.A1(net299),
    .A2(_0653_),
    .B1(_1342_),
    .C1(_2749_),
    .X(_2750_));
 sky130_fd_sc_hd__a21oi_1 _6144_ (.A1(net384),
    .A2(_2647_),
    .B1(_2750_),
    .Y(_2751_));
 sky130_fd_sc_hd__nor2_4 _6145_ (.A(_2748_),
    .B(_2751_),
    .Y(_2752_));
 sky130_fd_sc_hd__xor2_4 _6146_ (.A(_2679_),
    .B(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__xnor2_4 _6147_ (.A(_2745_),
    .B(_2753_),
    .Y(_2754_));
 sky130_fd_sc_hd__xnor2_4 _6148_ (.A(_2738_),
    .B(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__mux2_1 _6149_ (.A0(net585),
    .A1(_2755_),
    .S(_2642_),
    .X(_2756_));
 sky130_fd_sc_hd__clkbuf_1 _6150_ (.A(_2756_),
    .X(_0178_));
 sky130_fd_sc_hd__xnor2_4 _6151_ (.A(_2707_),
    .B(_2752_),
    .Y(_2757_));
 sky130_fd_sc_hd__xor2_1 _6152_ (.A(_2610_),
    .B(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__xnor2_1 _6153_ (.A(_2689_),
    .B(_2758_),
    .Y(_2759_));
 sky130_fd_sc_hd__xor2_2 _6154_ (.A(_2623_),
    .B(_2719_),
    .X(_2760_));
 sky130_fd_sc_hd__o21ai_1 _6155_ (.A1(_2759_),
    .A2(_2760_),
    .B1(_1217_),
    .Y(_2761_));
 sky130_fd_sc_hd__a21o_2 _6156_ (.A1(_2759_),
    .A2(_2760_),
    .B1(_2761_),
    .X(_2762_));
 sky130_fd_sc_hd__a22o_1 _6157_ (.A1(\sub1.data_o[83] ),
    .A2(_2699_),
    .B1(_2700_),
    .B2(\sub1.data_o[51] ),
    .X(_2763_));
 sky130_fd_sc_hd__a211o_1 _6158_ (.A1(\sub1.data_o[19] ),
    .A2(_0653_),
    .B1(_2546_),
    .C1(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__a21oi_2 _6159_ (.A1(\sub1.data_o[115] ),
    .A2(_2647_),
    .B1(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__a22o_1 _6160_ (.A1(net369),
    .A2(_2699_),
    .B1(_2700_),
    .B2(net334),
    .X(_2766_));
 sky130_fd_sc_hd__a211o_1 _6161_ (.A1(net298),
    .A2(_0653_),
    .B1(_1342_),
    .C1(_2766_),
    .X(_2767_));
 sky130_fd_sc_hd__a21oi_1 _6162_ (.A1(net277),
    .A2(_2647_),
    .B1(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__nor2_4 _6163_ (.A(_2765_),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__a22o_1 _6164_ (.A1(\sub1.data_o[66] ),
    .A2(_2533_),
    .B1(_2540_),
    .B2(\sub1.data_o[34] ),
    .X(_2770_));
 sky130_fd_sc_hd__a211o_1 _6165_ (.A1(\sub1.data_o[2] ),
    .A2(_0651_),
    .B1(_0807_),
    .C1(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__a21oi_1 _6166_ (.A1(\sub1.data_o[98] ),
    .A2(_2529_),
    .B1(_2771_),
    .Y(_2772_));
 sky130_fd_sc_hd__a22o_1 _6167_ (.A1(net350),
    .A2(_2533_),
    .B1(_2540_),
    .B2(net315),
    .X(_2773_));
 sky130_fd_sc_hd__a211o_1 _6168_ (.A1(net310),
    .A2(_0651_),
    .B1(_0798_),
    .C1(_2773_),
    .X(_2774_));
 sky130_fd_sc_hd__a21oi_1 _6169_ (.A1(net385),
    .A2(_2529_),
    .B1(_2774_),
    .Y(_2775_));
 sky130_fd_sc_hd__nor2_4 _6170_ (.A(_2772_),
    .B(_2775_),
    .Y(_2776_));
 sky130_fd_sc_hd__xnor2_2 _6171_ (.A(_2736_),
    .B(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__xnor2_1 _6172_ (.A(_2639_),
    .B(_2777_),
    .Y(_2778_));
 sky130_fd_sc_hd__xnor2_2 _6173_ (.A(_2769_),
    .B(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__a22o_1 _6174_ (.A1(\sub1.data_o[91] ),
    .A2(_2536_),
    .B1(_2543_),
    .B2(\sub1.data_o[59] ),
    .X(_2780_));
 sky130_fd_sc_hd__a211o_4 _6175_ (.A1(\sub1.data_o[27] ),
    .A2(_2680_),
    .B1(_2547_),
    .C1(_2780_),
    .X(_2781_));
 sky130_fd_sc_hd__a21oi_2 _6176_ (.A1(\sub1.data_o[123] ),
    .A2(_2531_),
    .B1(_2781_),
    .Y(_2782_));
 sky130_fd_sc_hd__a22o_1 _6177_ (.A1(net378),
    .A2(_2536_),
    .B1(_2543_),
    .B2(net342),
    .X(_2783_));
 sky130_fd_sc_hd__a211o_1 _6178_ (.A1(net307),
    .A2(_2680_),
    .B1(_1342_),
    .C1(_2783_),
    .X(_2784_));
 sky130_fd_sc_hd__a21oi_2 _6179_ (.A1(net286),
    .A2(_2531_),
    .B1(_2784_),
    .Y(_2785_));
 sky130_fd_sc_hd__nor2_8 _6180_ (.A(_2782_),
    .B(_2785_),
    .Y(_2786_));
 sky130_fd_sc_hd__a22o_1 _6181_ (.A1(\sub1.data_o[75] ),
    .A2(_2536_),
    .B1(_2543_),
    .B2(\sub1.data_o[43] ),
    .X(_2787_));
 sky130_fd_sc_hd__a211o_1 _6182_ (.A1(\sub1.data_o[11] ),
    .A2(_2680_),
    .B1(_2547_),
    .C1(_2787_),
    .X(_2788_));
 sky130_fd_sc_hd__a21oi_1 _6183_ (.A1(\sub1.data_o[107] ),
    .A2(_2612_),
    .B1(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__a22o_1 _6184_ (.A1(net360),
    .A2(_2536_),
    .B1(_2615_),
    .B2(net325),
    .X(_2790_));
 sky130_fd_sc_hd__a211o_1 _6185_ (.A1(net282),
    .A2(_2680_),
    .B1(_1343_),
    .C1(_2790_),
    .X(_2791_));
 sky130_fd_sc_hd__a21oi_1 _6186_ (.A1(net268),
    .A2(_2612_),
    .B1(_2791_),
    .Y(_2792_));
 sky130_fd_sc_hd__nor2_4 _6187_ (.A(_2789_),
    .B(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__xor2_2 _6188_ (.A(_2786_),
    .B(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__xnor2_2 _6189_ (.A(_2779_),
    .B(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__xnor2_4 _6190_ (.A(_2762_),
    .B(_2795_),
    .Y(_2796_));
 sky130_fd_sc_hd__mux2_1 _6191_ (.A0(net521),
    .A1(_2796_),
    .S(_2642_),
    .X(_2797_));
 sky130_fd_sc_hd__clkbuf_1 _6192_ (.A(_2797_),
    .X(_0179_));
 sky130_fd_sc_hd__xnor2_4 _6193_ (.A(_2708_),
    .B(_2776_),
    .Y(_2798_));
 sky130_fd_sc_hd__xor2_1 _6194_ (.A(_2754_),
    .B(_2798_),
    .X(_2799_));
 sky130_fd_sc_hd__o21ai_1 _6195_ (.A1(_2671_),
    .A2(_2799_),
    .B1(_1121_),
    .Y(_2800_));
 sky130_fd_sc_hd__a21o_1 _6196_ (.A1(_2671_),
    .A2(_2799_),
    .B1(_2800_),
    .X(_2801_));
 sky130_fd_sc_hd__a22o_1 _6197_ (.A1(\sub1.data_o[92] ),
    .A2(_2537_),
    .B1(_2615_),
    .B2(\sub1.data_o[60] ),
    .X(_2802_));
 sky130_fd_sc_hd__a211o_1 _6198_ (.A1(\sub1.data_o[28] ),
    .A2(_0654_),
    .B1(_2547_),
    .C1(_2802_),
    .X(_2803_));
 sky130_fd_sc_hd__a21o_2 _6199_ (.A1(\sub1.data_o[124] ),
    .A2(_2613_),
    .B1(_2803_),
    .X(_2804_));
 sky130_fd_sc_hd__a22o_1 _6200_ (.A1(net379),
    .A2(_2537_),
    .B1(_2615_),
    .B2(net344),
    .X(_2805_));
 sky130_fd_sc_hd__a211o_1 _6201_ (.A1(net308),
    .A2(_0654_),
    .B1(_1343_),
    .C1(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__a21o_1 _6202_ (.A1(net287),
    .A2(_2612_),
    .B1(_2806_),
    .X(_2807_));
 sky130_fd_sc_hd__nand2_8 _6203_ (.A(_2804_),
    .B(_2807_),
    .Y(_2808_));
 sky130_fd_sc_hd__a22o_1 _6204_ (.A1(\sub1.data_o[84] ),
    .A2(_2537_),
    .B1(_2615_),
    .B2(\sub1.data_o[52] ),
    .X(_2809_));
 sky130_fd_sc_hd__a211o_1 _6205_ (.A1(\sub1.data_o[20] ),
    .A2(_2680_),
    .B1(_2547_),
    .C1(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__a21oi_1 _6206_ (.A1(\sub1.data_o[116] ),
    .A2(_2612_),
    .B1(_2810_),
    .Y(_2811_));
 sky130_fd_sc_hd__a22o_1 _6207_ (.A1(net370),
    .A2(_2537_),
    .B1(_2615_),
    .B2(net335),
    .X(_2812_));
 sky130_fd_sc_hd__a211o_1 _6208_ (.A1(net300),
    .A2(_0654_),
    .B1(_1343_),
    .C1(_2812_),
    .X(_2813_));
 sky130_fd_sc_hd__a21oi_1 _6209_ (.A1(net278),
    .A2(_2612_),
    .B1(_2813_),
    .Y(_2814_));
 sky130_fd_sc_hd__nor2_4 _6210_ (.A(_2811_),
    .B(_2814_),
    .Y(_2815_));
 sky130_fd_sc_hd__xnor2_4 _6211_ (.A(_2808_),
    .B(_2815_),
    .Y(_2816_));
 sky130_fd_sc_hd__xor2_2 _6212_ (.A(_2801_),
    .B(_2816_),
    .X(_2817_));
 sky130_fd_sc_hd__a22o_1 _6213_ (.A1(\sub1.data_o[67] ),
    .A2(_2536_),
    .B1(_2615_),
    .B2(\sub1.data_o[35] ),
    .X(_2818_));
 sky130_fd_sc_hd__a211o_1 _6214_ (.A1(\sub1.data_o[3] ),
    .A2(_2680_),
    .B1(_2547_),
    .C1(_2818_),
    .X(_2819_));
 sky130_fd_sc_hd__a21oi_1 _6215_ (.A1(\sub1.data_o[99] ),
    .A2(_2612_),
    .B1(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__a22o_1 _6216_ (.A1(net351),
    .A2(_2537_),
    .B1(_2615_),
    .B2(net316),
    .X(_2821_));
 sky130_fd_sc_hd__a211o_1 _6217_ (.A1(net321),
    .A2(_2680_),
    .B1(_1343_),
    .C1(_2821_),
    .X(_2822_));
 sky130_fd_sc_hd__a21oi_1 _6218_ (.A1(net386),
    .A2(_2612_),
    .B1(_2822_),
    .Y(_2823_));
 sky130_fd_sc_hd__nor2_4 _6219_ (.A(_2820_),
    .B(_2823_),
    .Y(_2824_));
 sky130_fd_sc_hd__xnor2_4 _6220_ (.A(_2786_),
    .B(_2824_),
    .Y(_2825_));
 sky130_fd_sc_hd__xor2_2 _6221_ (.A(_2639_),
    .B(_2825_),
    .X(_2826_));
 sky130_fd_sc_hd__a22o_1 _6222_ (.A1(\sub1.data_o[76] ),
    .A2(_2537_),
    .B1(_2615_),
    .B2(\sub1.data_o[44] ),
    .X(_2827_));
 sky130_fd_sc_hd__a211o_1 _6223_ (.A1(\sub1.data_o[12] ),
    .A2(_2680_),
    .B1(_2547_),
    .C1(_2827_),
    .X(_2828_));
 sky130_fd_sc_hd__a21oi_1 _6224_ (.A1(\sub1.data_o[108] ),
    .A2(_2612_),
    .B1(_2828_),
    .Y(_2829_));
 sky130_fd_sc_hd__a22o_1 _6225_ (.A1(net361),
    .A2(_2537_),
    .B1(_2615_),
    .B2(net326),
    .X(_2830_));
 sky130_fd_sc_hd__a211o_1 _6226_ (.A1(net291),
    .A2(_2680_),
    .B1(_1343_),
    .C1(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__a21oi_2 _6227_ (.A1(net269),
    .A2(_2612_),
    .B1(_2831_),
    .Y(_2832_));
 sky130_fd_sc_hd__nor2_4 _6228_ (.A(_2829_),
    .B(_2832_),
    .Y(_2833_));
 sky130_fd_sc_hd__xor2_2 _6229_ (.A(_2826_),
    .B(_2833_),
    .X(_2834_));
 sky130_fd_sc_hd__xnor2_4 _6230_ (.A(_2817_),
    .B(_2834_),
    .Y(_2835_));
 sky130_fd_sc_hd__mux2_1 _6231_ (.A0(net529),
    .A1(_2835_),
    .S(_2642_),
    .X(_2836_));
 sky130_fd_sc_hd__clkbuf_1 _6232_ (.A(_2836_),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_1 _6233_ (.A1(\sub1.data_o[68] ),
    .A2(_2614_),
    .B1(_2616_),
    .B2(\sub1.data_o[36] ),
    .X(_2837_));
 sky130_fd_sc_hd__a211o_1 _6234_ (.A1(\sub1.data_o[4] ),
    .A2(_0654_),
    .B1(_2547_),
    .C1(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__a21oi_1 _6235_ (.A1(\sub1.data_o[100] ),
    .A2(_2613_),
    .B1(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__a22o_1 _6236_ (.A1(net352),
    .A2(_2614_),
    .B1(_2616_),
    .B2(net317),
    .X(_2840_));
 sky130_fd_sc_hd__a211o_1 _6237_ (.A1(net332),
    .A2(_0654_),
    .B1(_1343_),
    .C1(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__a21oi_2 _6238_ (.A1(net261),
    .A2(_2613_),
    .B1(_2841_),
    .Y(_2842_));
 sky130_fd_sc_hd__nor2_4 _6239_ (.A(_2839_),
    .B(_2842_),
    .Y(_2843_));
 sky130_fd_sc_hd__xor2_4 _6240_ (.A(_2808_),
    .B(_2843_),
    .X(_2844_));
 sky130_fd_sc_hd__xnor2_1 _6241_ (.A(_2729_),
    .B(_2745_),
    .Y(_2845_));
 sky130_fd_sc_hd__xnor2_1 _6242_ (.A(_2718_),
    .B(_2845_),
    .Y(_2846_));
 sky130_fd_sc_hd__xor2_1 _6243_ (.A(_2779_),
    .B(_2824_),
    .X(_2847_));
 sky130_fd_sc_hd__xnor2_1 _6244_ (.A(_2846_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__o21ai_1 _6245_ (.A1(_2670_),
    .A2(_2848_),
    .B1(_1121_),
    .Y(_2849_));
 sky130_fd_sc_hd__a21o_1 _6246_ (.A1(_2670_),
    .A2(_2848_),
    .B1(_2849_),
    .X(_2850_));
 sky130_fd_sc_hd__xor2_2 _6247_ (.A(_2568_),
    .B(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__xor2_4 _6248_ (.A(_2584_),
    .B(_2607_),
    .X(_2852_));
 sky130_fd_sc_hd__xnor2_2 _6249_ (.A(_2851_),
    .B(_2852_),
    .Y(_2853_));
 sky130_fd_sc_hd__xnor2_4 _6250_ (.A(_2844_),
    .B(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__mux2_1 _6251_ (.A0(net582),
    .A1(_2854_),
    .S(_2642_),
    .X(_2855_));
 sky130_fd_sc_hd__clkbuf_1 _6252_ (.A(_2855_),
    .X(_0181_));
 sky130_fd_sc_hd__xnor2_2 _6253_ (.A(_2718_),
    .B(_2769_),
    .Y(_2856_));
 sky130_fd_sc_hd__xnor2_4 _6254_ (.A(_2793_),
    .B(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__xnor2_4 _6255_ (.A(_2815_),
    .B(_2843_),
    .Y(_2858_));
 sky130_fd_sc_hd__xor2_1 _6256_ (.A(_2826_),
    .B(_2858_),
    .X(_2859_));
 sky130_fd_sc_hd__a21oi_1 _6257_ (.A1(_2857_),
    .A2(_2859_),
    .B1(_1214_),
    .Y(_2860_));
 sky130_fd_sc_hd__o21ai_2 _6258_ (.A1(_2857_),
    .A2(_2859_),
    .B1(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__xor2_4 _6259_ (.A(_2651_),
    .B(_2667_),
    .X(_2862_));
 sky130_fd_sc_hd__xnor2_4 _6260_ (.A(_2861_),
    .B(_2862_),
    .Y(_2863_));
 sky130_fd_sc_hd__xnor2_4 _6261_ (.A(_2609_),
    .B(_2863_),
    .Y(_2864_));
 sky130_fd_sc_hd__mux2_1 _6262_ (.A0(net566),
    .A1(_2864_),
    .S(_2642_),
    .X(_2865_));
 sky130_fd_sc_hd__clkbuf_1 _6263_ (.A(_2865_),
    .X(_0182_));
 sky130_fd_sc_hd__xor2_4 _6264_ (.A(_2638_),
    .B(_2659_),
    .X(_2866_));
 sky130_fd_sc_hd__xor2_4 _6265_ (.A(_2584_),
    .B(_2600_),
    .X(_2867_));
 sky130_fd_sc_hd__xor2_2 _6266_ (.A(_2815_),
    .B(_2833_),
    .X(_2868_));
 sky130_fd_sc_hd__xnor2_1 _6267_ (.A(_2867_),
    .B(_2868_),
    .Y(_2869_));
 sky130_fd_sc_hd__a21oi_1 _6268_ (.A1(_2844_),
    .A2(_2869_),
    .B1(_1214_),
    .Y(_2870_));
 sky130_fd_sc_hd__o21ai_2 _6269_ (.A1(_2844_),
    .A2(_2869_),
    .B1(_2870_),
    .Y(_2871_));
 sky130_fd_sc_hd__xnor2_2 _6270_ (.A(_2717_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__xnor2_2 _6271_ (.A(_2652_),
    .B(_2872_),
    .Y(_2873_));
 sky130_fd_sc_hd__xnor2_4 _6272_ (.A(_2866_),
    .B(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hd__mux2_1 _6273_ (.A0(net606),
    .A1(_2874_),
    .S(_2642_),
    .X(_2875_));
 sky130_fd_sc_hd__clkbuf_1 _6274_ (.A(_2875_),
    .X(_0183_));
 sky130_fd_sc_hd__xnor2_2 _6275_ (.A(_2568_),
    .B(_2600_),
    .Y(_2876_));
 sky130_fd_sc_hd__xor2_2 _6276_ (.A(_2852_),
    .B(_2876_),
    .X(_2877_));
 sky130_fd_sc_hd__xnor2_4 _6277_ (.A(_2862_),
    .B(_2877_),
    .Y(_2878_));
 sky130_fd_sc_hd__nand2_2 _6278_ (.A(_1218_),
    .B(_2878_),
    .Y(_2879_));
 sky130_fd_sc_hd__xnor2_1 _6279_ (.A(_2561_),
    .B(_2687_),
    .Y(_2880_));
 sky130_fd_sc_hd__xnor2_2 _6280_ (.A(_2879_),
    .B(_2880_),
    .Y(_2881_));
 sky130_fd_sc_hd__xnor2_4 _6281_ (.A(_2631_),
    .B(_2717_),
    .Y(_2882_));
 sky130_fd_sc_hd__xnor2_4 _6282_ (.A(_2881_),
    .B(_2882_),
    .Y(_2883_));
 sky130_fd_sc_hd__mux2_1 _6283_ (.A0(net596),
    .A1(_2883_),
    .S(_2642_),
    .X(_2884_));
 sky130_fd_sc_hd__clkbuf_1 _6284_ (.A(_2884_),
    .X(_0184_));
 sky130_fd_sc_hd__xor2_4 _6285_ (.A(_2623_),
    .B(_2687_),
    .X(_2885_));
 sky130_fd_sc_hd__xnor2_2 _6286_ (.A(_2679_),
    .B(_2882_),
    .Y(_2886_));
 sky130_fd_sc_hd__xnor2_4 _6287_ (.A(_2885_),
    .B(_2886_),
    .Y(_2887_));
 sky130_fd_sc_hd__xnor2_4 _6288_ (.A(_2575_),
    .B(_2667_),
    .Y(_2888_));
 sky130_fd_sc_hd__xnor2_4 _6289_ (.A(_2638_),
    .B(_2888_),
    .Y(_2889_));
 sky130_fd_sc_hd__xnor2_4 _6290_ (.A(_2593_),
    .B(_2651_),
    .Y(_2890_));
 sky130_fd_sc_hd__xor2_2 _6291_ (.A(_2717_),
    .B(_2890_),
    .X(_2891_));
 sky130_fd_sc_hd__xnor2_4 _6292_ (.A(_2889_),
    .B(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__xor2_2 _6293_ (.A(_2878_),
    .B(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__nand2_2 _6294_ (.A(_1218_),
    .B(_2893_),
    .Y(_2894_));
 sky130_fd_sc_hd__xnor2_4 _6295_ (.A(_2757_),
    .B(_2894_),
    .Y(_2895_));
 sky130_fd_sc_hd__xnor2_2 _6296_ (.A(_2887_),
    .B(_2895_),
    .Y(_2896_));
 sky130_fd_sc_hd__buf_4 _6297_ (.A(_2614_),
    .X(_2897_));
 sky130_fd_sc_hd__mux2_1 _6298_ (.A0(net534),
    .A1(_2896_),
    .S(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__clkbuf_1 _6299_ (.A(_2898_),
    .X(_0185_));
 sky130_fd_sc_hd__xor2_1 _6300_ (.A(_2560_),
    .B(_2882_),
    .X(_2899_));
 sky130_fd_sc_hd__xnor2_1 _6301_ (.A(_2623_),
    .B(_2899_),
    .Y(_2900_));
 sky130_fd_sc_hd__xnor2_1 _6302_ (.A(_2866_),
    .B(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__o21ai_1 _6303_ (.A1(_2892_),
    .A2(_2901_),
    .B1(_1218_),
    .Y(_2902_));
 sky130_fd_sc_hd__a21o_2 _6304_ (.A1(_2892_),
    .A2(_2901_),
    .B1(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__xnor2_1 _6305_ (.A(_2698_),
    .B(_2752_),
    .Y(_2904_));
 sky130_fd_sc_hd__xnor2_1 _6306_ (.A(_2745_),
    .B(_2777_),
    .Y(_2905_));
 sky130_fd_sc_hd__xnor2_2 _6307_ (.A(_2904_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__xnor2_4 _6308_ (.A(_2903_),
    .B(_2906_),
    .Y(_2907_));
 sky130_fd_sc_hd__mux2_1 _6309_ (.A0(net555),
    .A1(_2907_),
    .S(_2897_),
    .X(_2908_));
 sky130_fd_sc_hd__clkbuf_1 _6310_ (.A(_2908_),
    .X(_0186_));
 sky130_fd_sc_hd__xor2_1 _6311_ (.A(_2561_),
    .B(_2698_),
    .X(_2909_));
 sky130_fd_sc_hd__xnor2_2 _6312_ (.A(_2866_),
    .B(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hd__xor2_2 _6313_ (.A(_2878_),
    .B(_2910_),
    .X(_2911_));
 sky130_fd_sc_hd__a21oi_1 _6314_ (.A1(_2887_),
    .A2(_2911_),
    .B1(_1214_),
    .Y(_2912_));
 sky130_fd_sc_hd__o21ai_4 _6315_ (.A1(_2887_),
    .A2(_2911_),
    .B1(_2912_),
    .Y(_2913_));
 sky130_fd_sc_hd__xnor2_4 _6316_ (.A(_2729_),
    .B(_2776_),
    .Y(_2914_));
 sky130_fd_sc_hd__xnor2_2 _6317_ (.A(_2882_),
    .B(_2914_),
    .Y(_2915_));
 sky130_fd_sc_hd__xnor2_1 _6318_ (.A(_2769_),
    .B(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__xnor2_2 _6319_ (.A(_2825_),
    .B(_2916_),
    .Y(_2917_));
 sky130_fd_sc_hd__xnor2_2 _6320_ (.A(_2913_),
    .B(_2917_),
    .Y(_2918_));
 sky130_fd_sc_hd__mux2_1 _6321_ (.A0(net553),
    .A1(_2918_),
    .S(_2897_),
    .X(_2919_));
 sky130_fd_sc_hd__clkbuf_1 _6322_ (.A(_2919_),
    .X(_0187_));
 sky130_fd_sc_hd__xnor2_1 _6323_ (.A(_2708_),
    .B(_2737_),
    .Y(_2920_));
 sky130_fd_sc_hd__xnor2_2 _6324_ (.A(_2753_),
    .B(_2920_),
    .Y(_2921_));
 sky130_fd_sc_hd__a21oi_1 _6325_ (.A1(_2893_),
    .A2(_2921_),
    .B1(_1214_),
    .Y(_2922_));
 sky130_fd_sc_hd__o21ai_2 _6326_ (.A1(_2893_),
    .A2(_2921_),
    .B1(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__xnor2_4 _6327_ (.A(_2858_),
    .B(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__xor2_4 _6328_ (.A(_2793_),
    .B(_2824_),
    .X(_2925_));
 sky130_fd_sc_hd__xor2_2 _6329_ (.A(_2882_),
    .B(_2925_),
    .X(_2926_));
 sky130_fd_sc_hd__xnor2_4 _6330_ (.A(_2808_),
    .B(_2926_),
    .Y(_2927_));
 sky130_fd_sc_hd__xnor2_2 _6331_ (.A(_2924_),
    .B(_2927_),
    .Y(_2928_));
 sky130_fd_sc_hd__mux2_1 _6332_ (.A0(net532),
    .A1(_2928_),
    .S(_2897_),
    .X(_2929_));
 sky130_fd_sc_hd__clkbuf_1 _6333_ (.A(_2929_),
    .X(_0188_));
 sky130_fd_sc_hd__xor2_2 _6334_ (.A(_2736_),
    .B(_2745_),
    .X(_2930_));
 sky130_fd_sc_hd__xnor2_2 _6335_ (.A(_2866_),
    .B(_2930_),
    .Y(_2931_));
 sky130_fd_sc_hd__xnor2_1 _6336_ (.A(_2794_),
    .B(_2915_),
    .Y(_2932_));
 sky130_fd_sc_hd__xor2_1 _6337_ (.A(_2931_),
    .B(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__a21oi_1 _6338_ (.A1(_2892_),
    .A2(_2933_),
    .B1(_1214_),
    .Y(_2934_));
 sky130_fd_sc_hd__o21ai_1 _6339_ (.A1(_2892_),
    .A2(_2933_),
    .B1(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__xnor2_2 _6340_ (.A(_2867_),
    .B(_2935_),
    .Y(_2936_));
 sky130_fd_sc_hd__xor2_2 _6341_ (.A(_2833_),
    .B(_2843_),
    .X(_2937_));
 sky130_fd_sc_hd__xnor2_4 _6342_ (.A(_2607_),
    .B(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__xnor2_2 _6343_ (.A(_2936_),
    .B(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__mux2_1 _6344_ (.A0(net613),
    .A1(_2939_),
    .S(_2897_),
    .X(_2940_));
 sky130_fd_sc_hd__clkbuf_1 _6345_ (.A(_2940_),
    .X(_0189_));
 sky130_fd_sc_hd__xnor2_2 _6346_ (.A(_2575_),
    .B(_2876_),
    .Y(_2941_));
 sky130_fd_sc_hd__xor2_2 _6347_ (.A(_2769_),
    .B(_2786_),
    .X(_2942_));
 sky130_fd_sc_hd__xnor2_2 _6348_ (.A(_2833_),
    .B(_2866_),
    .Y(_2943_));
 sky130_fd_sc_hd__xnor2_4 _6349_ (.A(_2942_),
    .B(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__a21oi_2 _6350_ (.A1(_2927_),
    .A2(_2944_),
    .B1(_1214_),
    .Y(_2945_));
 sky130_fd_sc_hd__o21ai_4 _6351_ (.A1(_2927_),
    .A2(_2944_),
    .B1(_2945_),
    .Y(_2946_));
 sky130_fd_sc_hd__xnor2_1 _6352_ (.A(_2890_),
    .B(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__xnor2_2 _6353_ (.A(_2941_),
    .B(_2947_),
    .Y(_2948_));
 sky130_fd_sc_hd__mux2_1 _6354_ (.A0(net602),
    .A1(_2948_),
    .S(_2897_),
    .X(_2949_));
 sky130_fd_sc_hd__clkbuf_1 _6355_ (.A(_2949_),
    .X(_0190_));
 sky130_fd_sc_hd__xnor2_4 _6356_ (.A(_2568_),
    .B(_2816_),
    .Y(_2950_));
 sky130_fd_sc_hd__a21oi_1 _6357_ (.A1(_2938_),
    .A2(_2950_),
    .B1(_1214_),
    .Y(_2951_));
 sky130_fd_sc_hd__o21ai_4 _6358_ (.A1(_2938_),
    .A2(_2950_),
    .B1(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__xnor2_1 _6359_ (.A(_2660_),
    .B(_2889_),
    .Y(_2953_));
 sky130_fd_sc_hd__xor2_2 _6360_ (.A(_2952_),
    .B(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__mux2_1 _6361_ (.A0(net597),
    .A1(_2954_),
    .S(_2897_),
    .X(_2955_));
 sky130_fd_sc_hd__clkbuf_1 _6362_ (.A(_2955_),
    .X(_0191_));
 sky130_fd_sc_hd__xnor2_1 _6363_ (.A(_2560_),
    .B(_2687_),
    .Y(_2956_));
 sky130_fd_sc_hd__xnor2_2 _6364_ (.A(_2624_),
    .B(_2956_),
    .Y(_2957_));
 sky130_fd_sc_hd__xnor2_4 _6365_ (.A(_2718_),
    .B(_2957_),
    .Y(_2958_));
 sky130_fd_sc_hd__mux2_1 _6366_ (.A0(net524),
    .A1(_2958_),
    .S(_2897_),
    .X(_2959_));
 sky130_fd_sc_hd__clkbuf_1 _6367_ (.A(_2959_),
    .X(_0192_));
 sky130_fd_sc_hd__xnor2_1 _6368_ (.A(_2753_),
    .B(_2760_),
    .Y(_2960_));
 sky130_fd_sc_hd__xnor2_1 _6369_ (.A(_2672_),
    .B(_2960_),
    .Y(_2961_));
 sky130_fd_sc_hd__xnor2_2 _6370_ (.A(_2698_),
    .B(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__mux2_1 _6371_ (.A0(net548),
    .A1(_2962_),
    .S(_2897_),
    .X(_2963_));
 sky130_fd_sc_hd__clkbuf_1 _6372_ (.A(_2963_),
    .X(_0193_));
 sky130_fd_sc_hd__xnor2_4 _6373_ (.A(_2738_),
    .B(_2798_),
    .Y(_2964_));
 sky130_fd_sc_hd__mux2_1 _6374_ (.A0(net549),
    .A1(_2964_),
    .S(_2897_),
    .X(_2965_));
 sky130_fd_sc_hd__clkbuf_1 _6375_ (.A(_2965_),
    .X(_0194_));
 sky130_fd_sc_hd__xnor2_2 _6376_ (.A(_2786_),
    .B(_2925_),
    .Y(_2966_));
 sky130_fd_sc_hd__xnor2_1 _6377_ (.A(_2762_),
    .B(_2846_),
    .Y(_2967_));
 sky130_fd_sc_hd__xnor2_2 _6378_ (.A(_2966_),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__buf_4 _6379_ (.A(_2614_),
    .X(_2969_));
 sky130_fd_sc_hd__mux2_1 _6380_ (.A0(net572),
    .A1(_2968_),
    .S(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__clkbuf_1 _6381_ (.A(_2970_),
    .X(_0195_));
 sky130_fd_sc_hd__xnor2_1 _6382_ (.A(_2801_),
    .B(_2833_),
    .Y(_2971_));
 sky130_fd_sc_hd__xnor2_1 _6383_ (.A(_2844_),
    .B(_2971_),
    .Y(_2972_));
 sky130_fd_sc_hd__xnor2_2 _6384_ (.A(_2857_),
    .B(_2972_),
    .Y(_2973_));
 sky130_fd_sc_hd__mux2_1 _6385_ (.A0(net588),
    .A1(_2973_),
    .S(_2969_),
    .X(_2974_));
 sky130_fd_sc_hd__clkbuf_1 _6386_ (.A(_2974_),
    .X(_0196_));
 sky130_fd_sc_hd__xor2_1 _6387_ (.A(_2608_),
    .B(_2851_),
    .X(_2975_));
 sky130_fd_sc_hd__xor2_2 _6388_ (.A(_2868_),
    .B(_2975_),
    .X(_2976_));
 sky130_fd_sc_hd__mux2_1 _6389_ (.A0(net525),
    .A1(_2976_),
    .S(_2969_),
    .X(_2977_));
 sky130_fd_sc_hd__clkbuf_1 _6390_ (.A(_2977_),
    .X(_0197_));
 sky130_fd_sc_hd__xnor2_2 _6391_ (.A(_2586_),
    .B(_2863_),
    .Y(_2978_));
 sky130_fd_sc_hd__mux2_1 _6392_ (.A0(net565),
    .A1(_2978_),
    .S(_2969_),
    .X(_2979_));
 sky130_fd_sc_hd__clkbuf_1 _6393_ (.A(_2979_),
    .X(_0198_));
 sky130_fd_sc_hd__xor2_1 _6394_ (.A(_2639_),
    .B(_2872_),
    .X(_2980_));
 sky130_fd_sc_hd__xnor2_2 _6395_ (.A(_2668_),
    .B(_2980_),
    .Y(_2981_));
 sky130_fd_sc_hd__mux2_1 _6396_ (.A0(net611),
    .A1(_2981_),
    .S(_2969_),
    .X(_2982_));
 sky130_fd_sc_hd__clkbuf_1 _6397_ (.A(_2982_),
    .X(_0199_));
 sky130_fd_sc_hd__xnor2_1 _6398_ (.A(_2866_),
    .B(_2885_),
    .Y(_2983_));
 sky130_fd_sc_hd__xnor2_1 _6399_ (.A(_2553_),
    .B(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__xnor2_2 _6400_ (.A(_2879_),
    .B(_2984_),
    .Y(_2985_));
 sky130_fd_sc_hd__mux2_1 _6401_ (.A0(net556),
    .A1(_2985_),
    .S(_2969_),
    .X(_2986_));
 sky130_fd_sc_hd__clkbuf_1 _6402_ (.A(_2986_),
    .X(_0200_));
 sky130_fd_sc_hd__xnor2_2 _6403_ (.A(_2895_),
    .B(_2910_),
    .Y(_2987_));
 sky130_fd_sc_hd__mux2_1 _6404_ (.A0(net633),
    .A1(_2987_),
    .S(_2969_),
    .X(_2988_));
 sky130_fd_sc_hd__clkbuf_1 _6405_ (.A(_2988_),
    .X(_0201_));
 sky130_fd_sc_hd__xnor2_1 _6406_ (.A(_2679_),
    .B(_2745_),
    .Y(_2989_));
 sky130_fd_sc_hd__xnor2_1 _6407_ (.A(_2707_),
    .B(_2989_),
    .Y(_2990_));
 sky130_fd_sc_hd__xnor2_2 _6408_ (.A(_2914_),
    .B(_2990_),
    .Y(_2991_));
 sky130_fd_sc_hd__xor2_4 _6409_ (.A(_2903_),
    .B(_2991_),
    .X(_2992_));
 sky130_fd_sc_hd__mux2_1 _6410_ (.A0(net576),
    .A1(_2992_),
    .S(_2969_),
    .X(_2993_));
 sky130_fd_sc_hd__clkbuf_1 _6411_ (.A(_2993_),
    .X(_0202_));
 sky130_fd_sc_hd__xnor2_1 _6412_ (.A(_2769_),
    .B(_2925_),
    .Y(_2994_));
 sky130_fd_sc_hd__xnor2_2 _6413_ (.A(_2931_),
    .B(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__xnor2_2 _6414_ (.A(_2913_),
    .B(_2995_),
    .Y(_2996_));
 sky130_fd_sc_hd__mux2_1 _6415_ (.A0(net601),
    .A1(_2996_),
    .S(_2969_),
    .X(_2997_));
 sky130_fd_sc_hd__clkbuf_1 _6416_ (.A(_2997_),
    .X(_0203_));
 sky130_fd_sc_hd__xnor2_2 _6417_ (.A(_2924_),
    .B(_2944_),
    .Y(_2998_));
 sky130_fd_sc_hd__mux2_1 _6418_ (.A0(net591),
    .A1(_2998_),
    .S(_2969_),
    .X(_2999_));
 sky130_fd_sc_hd__clkbuf_1 _6419_ (.A(_2999_),
    .X(_0204_));
 sky130_fd_sc_hd__xnor2_2 _6420_ (.A(_2936_),
    .B(_2950_),
    .Y(_3000_));
 sky130_fd_sc_hd__mux2_1 _6421_ (.A0(net527),
    .A1(_3000_),
    .S(_2614_),
    .X(_3001_));
 sky130_fd_sc_hd__clkbuf_1 _6422_ (.A(_3001_),
    .X(_0205_));
 sky130_fd_sc_hd__xor2_2 _6423_ (.A(_2593_),
    .B(_2888_),
    .X(_3002_));
 sky130_fd_sc_hd__xnor2_4 _6424_ (.A(_2852_),
    .B(_3002_),
    .Y(_3003_));
 sky130_fd_sc_hd__xnor2_4 _6425_ (.A(_2946_),
    .B(_3003_),
    .Y(_3004_));
 sky130_fd_sc_hd__mux2_1 _6426_ (.A0(net547),
    .A1(_3004_),
    .S(_2614_),
    .X(_3005_));
 sky130_fd_sc_hd__clkbuf_1 _6427_ (.A(_3005_),
    .X(_0206_));
 sky130_fd_sc_hd__xnor2_1 _6428_ (.A(_2659_),
    .B(_2890_),
    .Y(_3006_));
 sky130_fd_sc_hd__xnor2_1 _6429_ (.A(_2882_),
    .B(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__xnor2_2 _6430_ (.A(_2952_),
    .B(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__mux2_1 _6431_ (.A0(net554),
    .A1(_3008_),
    .S(_2614_),
    .X(_3009_));
 sky130_fd_sc_hd__clkbuf_1 _6432_ (.A(_3009_),
    .X(_0207_));
 sky130_fd_sc_hd__buf_4 _6433_ (.A(_2616_),
    .X(_3010_));
 sky130_fd_sc_hd__mux2_1 _6434_ (.A0(net608),
    .A1(_2641_),
    .S(_3010_),
    .X(_3011_));
 sky130_fd_sc_hd__clkbuf_1 _6435_ (.A(_3011_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _6436_ (.A0(net605),
    .A1(_2709_),
    .S(_3010_),
    .X(_3012_));
 sky130_fd_sc_hd__clkbuf_1 _6437_ (.A(_3012_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _6438_ (.A0(net559),
    .A1(_2755_),
    .S(_3010_),
    .X(_3013_));
 sky130_fd_sc_hd__clkbuf_1 _6439_ (.A(_3013_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _6440_ (.A0(net550),
    .A1(_2796_),
    .S(_3010_),
    .X(_3014_));
 sky130_fd_sc_hd__clkbuf_1 _6441_ (.A(_3014_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _6442_ (.A0(net587),
    .A1(_2835_),
    .S(_3010_),
    .X(_3015_));
 sky130_fd_sc_hd__clkbuf_1 _6443_ (.A(_3015_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _6444_ (.A0(net583),
    .A1(_2854_),
    .S(_3010_),
    .X(_3016_));
 sky130_fd_sc_hd__clkbuf_1 _6445_ (.A(_3016_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _6446_ (.A0(net544),
    .A1(_2864_),
    .S(_3010_),
    .X(_3017_));
 sky130_fd_sc_hd__clkbuf_1 _6447_ (.A(_3017_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _6448_ (.A0(net577),
    .A1(_2874_),
    .S(_3010_),
    .X(_3018_));
 sky130_fd_sc_hd__clkbuf_1 _6449_ (.A(_3018_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _6450_ (.A0(net546),
    .A1(_2883_),
    .S(_3010_),
    .X(_3019_));
 sky130_fd_sc_hd__clkbuf_1 _6451_ (.A(_3019_),
    .X(_0216_));
 sky130_fd_sc_hd__buf_4 _6452_ (.A(_2616_),
    .X(_3020_));
 sky130_fd_sc_hd__mux2_1 _6453_ (.A0(net531),
    .A1(_2896_),
    .S(_3020_),
    .X(_3021_));
 sky130_fd_sc_hd__clkbuf_1 _6454_ (.A(_3021_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _6455_ (.A0(net557),
    .A1(_2907_),
    .S(_3020_),
    .X(_3022_));
 sky130_fd_sc_hd__clkbuf_1 _6456_ (.A(_3022_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _6457_ (.A0(net578),
    .A1(_2918_),
    .S(_3020_),
    .X(_3023_));
 sky130_fd_sc_hd__clkbuf_1 _6458_ (.A(_3023_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _6459_ (.A0(net609),
    .A1(_2928_),
    .S(_3020_),
    .X(_3024_));
 sky130_fd_sc_hd__clkbuf_1 _6460_ (.A(_3024_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _6461_ (.A0(net533),
    .A1(_2939_),
    .S(_3020_),
    .X(_3025_));
 sky130_fd_sc_hd__clkbuf_1 _6462_ (.A(_3025_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _6463_ (.A0(net619),
    .A1(_2948_),
    .S(_3020_),
    .X(_3026_));
 sky130_fd_sc_hd__clkbuf_1 _6464_ (.A(_3026_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _6465_ (.A0(net618),
    .A1(_2954_),
    .S(_3020_),
    .X(_3027_));
 sky130_fd_sc_hd__clkbuf_1 _6466_ (.A(_3027_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _6467_ (.A0(net600),
    .A1(_2958_),
    .S(_3020_),
    .X(_3028_));
 sky130_fd_sc_hd__clkbuf_1 _6468_ (.A(_3028_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _6469_ (.A0(net579),
    .A1(_2962_),
    .S(_3020_),
    .X(_3029_));
 sky130_fd_sc_hd__clkbuf_1 _6470_ (.A(_3029_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _6471_ (.A0(net594),
    .A1(_2964_),
    .S(_3020_),
    .X(_3030_));
 sky130_fd_sc_hd__clkbuf_1 _6472_ (.A(_3030_),
    .X(_0226_));
 sky130_fd_sc_hd__buf_4 _6473_ (.A(_2616_),
    .X(_3031_));
 sky130_fd_sc_hd__mux2_1 _6474_ (.A0(net536),
    .A1(_2968_),
    .S(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__clkbuf_1 _6475_ (.A(_3032_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _6476_ (.A0(net573),
    .A1(_2973_),
    .S(_3031_),
    .X(_3033_));
 sky130_fd_sc_hd__clkbuf_1 _6477_ (.A(_3033_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _6478_ (.A0(net545),
    .A1(_2976_),
    .S(_3031_),
    .X(_3034_));
 sky130_fd_sc_hd__clkbuf_1 _6479_ (.A(_3034_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _6480_ (.A0(net589),
    .A1(_2978_),
    .S(_3031_),
    .X(_3035_));
 sky130_fd_sc_hd__clkbuf_1 _6481_ (.A(_3035_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _6482_ (.A0(net623),
    .A1(_2981_),
    .S(_3031_),
    .X(_3036_));
 sky130_fd_sc_hd__clkbuf_1 _6483_ (.A(_3036_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _6484_ (.A0(net552),
    .A1(_2985_),
    .S(_3031_),
    .X(_3037_));
 sky130_fd_sc_hd__clkbuf_1 _6485_ (.A(_3037_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _6486_ (.A0(net560),
    .A1(_2987_),
    .S(_3031_),
    .X(_3038_));
 sky130_fd_sc_hd__clkbuf_1 _6487_ (.A(_3038_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _6488_ (.A0(net558),
    .A1(_2992_),
    .S(_3031_),
    .X(_3039_));
 sky130_fd_sc_hd__clkbuf_1 _6489_ (.A(_3039_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _6490_ (.A0(net530),
    .A1(_2996_),
    .S(_3031_),
    .X(_3040_));
 sky130_fd_sc_hd__clkbuf_1 _6491_ (.A(_3040_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _6492_ (.A0(net604),
    .A1(_2998_),
    .S(_3031_),
    .X(_3041_));
 sky130_fd_sc_hd__clkbuf_1 _6493_ (.A(_3041_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _6494_ (.A0(net603),
    .A1(_3000_),
    .S(_2616_),
    .X(_3042_));
 sky130_fd_sc_hd__clkbuf_1 _6495_ (.A(_3042_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _6496_ (.A0(net535),
    .A1(_3004_),
    .S(_2616_),
    .X(_3043_));
 sky130_fd_sc_hd__clkbuf_1 _6497_ (.A(_3043_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _6498_ (.A0(net599),
    .A1(_3008_),
    .S(_2616_),
    .X(_3044_));
 sky130_fd_sc_hd__clkbuf_1 _6499_ (.A(_3044_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _6500_ (.A0(\sub1.data_o[120] ),
    .A1(_1212_),
    .S(_0911_),
    .X(_3045_));
 sky130_fd_sc_hd__clkbuf_1 _6501_ (.A(_3045_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _6502_ (.A0(\sub1.data_o[121] ),
    .A1(_1246_),
    .S(_0911_),
    .X(_3046_));
 sky130_fd_sc_hd__clkbuf_1 _6503_ (.A(_3046_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _6504_ (.A0(\sub1.data_o[122] ),
    .A1(_1256_),
    .S(_0911_),
    .X(_3047_));
 sky130_fd_sc_hd__clkbuf_1 _6505_ (.A(_3047_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _6506_ (.A0(\sub1.data_o[123] ),
    .A1(_1272_),
    .S(_0911_),
    .X(_3048_));
 sky130_fd_sc_hd__clkbuf_1 _6507_ (.A(_3048_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _6508_ (.A0(\sub1.data_o[124] ),
    .A1(_1277_),
    .S(_0911_),
    .X(_3049_));
 sky130_fd_sc_hd__clkbuf_1 _6509_ (.A(_3049_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _6510_ (.A0(\sub1.data_o[125] ),
    .A1(_1285_),
    .S(_0911_),
    .X(_3050_));
 sky130_fd_sc_hd__clkbuf_1 _6511_ (.A(_3050_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _6512_ (.A0(\sub1.data_o[126] ),
    .A1(_1292_),
    .S(_0911_),
    .X(_3051_));
 sky130_fd_sc_hd__clkbuf_1 _6513_ (.A(_3051_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _6514_ (.A0(\sub1.data_o[127] ),
    .A1(_1299_),
    .S(_0911_),
    .X(_3052_));
 sky130_fd_sc_hd__clkbuf_1 _6515_ (.A(_3052_),
    .X(_0247_));
 sky130_fd_sc_hd__buf_4 _6516_ (.A(_1218_),
    .X(_3053_));
 sky130_fd_sc_hd__mux2_1 _6517_ (.A0(\sub1.data_o[32] ),
    .A1(\sub1.data_o[96] ),
    .S(_3053_),
    .X(_3054_));
 sky130_fd_sc_hd__buf_4 _6518_ (.A(_0662_),
    .X(_3055_));
 sky130_fd_sc_hd__mux2_1 _6519_ (.A0(\sub1.data_o[0] ),
    .A1(_3054_),
    .S(_3055_),
    .X(_3056_));
 sky130_fd_sc_hd__clkbuf_1 _6520_ (.A(_3056_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _6521_ (.A0(\sub1.data_o[33] ),
    .A1(\sub1.data_o[97] ),
    .S(_3053_),
    .X(_3057_));
 sky130_fd_sc_hd__mux2_1 _6522_ (.A0(\sub1.data_o[1] ),
    .A1(_3057_),
    .S(_3055_),
    .X(_3058_));
 sky130_fd_sc_hd__clkbuf_1 _6523_ (.A(_3058_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _6524_ (.A0(\sub1.data_o[34] ),
    .A1(\sub1.data_o[98] ),
    .S(_3053_),
    .X(_3059_));
 sky130_fd_sc_hd__mux2_1 _6525_ (.A0(\sub1.data_o[2] ),
    .A1(_3059_),
    .S(_3055_),
    .X(_3060_));
 sky130_fd_sc_hd__clkbuf_1 _6526_ (.A(_3060_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _6527_ (.A0(\sub1.data_o[35] ),
    .A1(\sub1.data_o[99] ),
    .S(_3053_),
    .X(_3061_));
 sky130_fd_sc_hd__mux2_1 _6528_ (.A0(\sub1.data_o[3] ),
    .A1(_3061_),
    .S(_3055_),
    .X(_3062_));
 sky130_fd_sc_hd__clkbuf_1 _6529_ (.A(_3062_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _6530_ (.A0(\sub1.data_o[36] ),
    .A1(\sub1.data_o[100] ),
    .S(_3053_),
    .X(_3063_));
 sky130_fd_sc_hd__mux2_1 _6531_ (.A0(\sub1.data_o[4] ),
    .A1(_3063_),
    .S(_2491_),
    .X(_3064_));
 sky130_fd_sc_hd__clkbuf_1 _6532_ (.A(_3064_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _6533_ (.A0(\sub1.data_o[37] ),
    .A1(\sub1.data_o[101] ),
    .S(_3053_),
    .X(_3065_));
 sky130_fd_sc_hd__mux2_1 _6534_ (.A0(\sub1.data_o[5] ),
    .A1(_3065_),
    .S(_2491_),
    .X(_3066_));
 sky130_fd_sc_hd__clkbuf_1 _6535_ (.A(_3066_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _6536_ (.A0(\sub1.data_o[38] ),
    .A1(\sub1.data_o[102] ),
    .S(_1218_),
    .X(_3067_));
 sky130_fd_sc_hd__mux2_1 _6537_ (.A0(\sub1.data_o[6] ),
    .A1(_3067_),
    .S(_2491_),
    .X(_3068_));
 sky130_fd_sc_hd__clkbuf_1 _6538_ (.A(_3068_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _6539_ (.A0(\sub1.data_o[39] ),
    .A1(\sub1.data_o[103] ),
    .S(_1218_),
    .X(_3069_));
 sky130_fd_sc_hd__mux2_1 _6540_ (.A0(\sub1.data_o[7] ),
    .A1(_3069_),
    .S(_2491_),
    .X(_3070_));
 sky130_fd_sc_hd__clkbuf_1 _6541_ (.A(_3070_),
    .X(_0255_));
 sky130_fd_sc_hd__clkbuf_4 _6542_ (.A(_0712_),
    .X(_3071_));
 sky130_fd_sc_hd__nor2_2 _6543_ (.A(_2491_),
    .B(_0712_),
    .Y(_3072_));
 sky130_fd_sc_hd__a22o_1 _6544_ (.A1(\sub1.data_o[72] ),
    .A2(_2500_),
    .B1(_3072_),
    .B2(\sub1.data_o[8] ),
    .X(_3073_));
 sky130_fd_sc_hd__a31o_1 _6545_ (.A1(_2495_),
    .A2(_3071_),
    .A3(_1213_),
    .B1(_3073_),
    .X(_0256_));
 sky130_fd_sc_hd__a22o_1 _6546_ (.A1(\sub1.data_o[73] ),
    .A2(_2500_),
    .B1(_3072_),
    .B2(\sub1.data_o[9] ),
    .X(_3074_));
 sky130_fd_sc_hd__a31o_1 _6547_ (.A1(_2495_),
    .A2(_3071_),
    .A3(_1247_),
    .B1(_3074_),
    .X(_0257_));
 sky130_fd_sc_hd__a22o_1 _6548_ (.A1(\sub1.data_o[74] ),
    .A2(_2500_),
    .B1(_3072_),
    .B2(\sub1.data_o[10] ),
    .X(_3075_));
 sky130_fd_sc_hd__a31o_1 _6549_ (.A1(_2495_),
    .A2(_3071_),
    .A3(_1257_),
    .B1(_3075_),
    .X(_0258_));
 sky130_fd_sc_hd__a22o_1 _6550_ (.A1(\sub1.data_o[75] ),
    .A2(_2500_),
    .B1(_3072_),
    .B2(\sub1.data_o[11] ),
    .X(_3076_));
 sky130_fd_sc_hd__a31o_1 _6551_ (.A1(_2495_),
    .A2(_3071_),
    .A3(_1272_),
    .B1(_3076_),
    .X(_0259_));
 sky130_fd_sc_hd__clkbuf_4 _6552_ (.A(_1139_),
    .X(_3077_));
 sky130_fd_sc_hd__a22o_1 _6553_ (.A1(\sub1.data_o[76] ),
    .A2(_2500_),
    .B1(_3072_),
    .B2(\sub1.data_o[12] ),
    .X(_3078_));
 sky130_fd_sc_hd__a31o_1 _6554_ (.A1(_3077_),
    .A2(_3071_),
    .A3(_1278_),
    .B1(_3078_),
    .X(_0260_));
 sky130_fd_sc_hd__a22o_1 _6555_ (.A1(\sub1.data_o[77] ),
    .A2(_2500_),
    .B1(_3072_),
    .B2(\sub1.data_o[13] ),
    .X(_3079_));
 sky130_fd_sc_hd__a31o_1 _6556_ (.A1(_3077_),
    .A2(_3071_),
    .A3(_1286_),
    .B1(_3079_),
    .X(_0261_));
 sky130_fd_sc_hd__a22o_1 _6557_ (.A1(\sub1.data_o[78] ),
    .A2(_2500_),
    .B1(_3072_),
    .B2(\sub1.data_o[14] ),
    .X(_3080_));
 sky130_fd_sc_hd__a31o_1 _6558_ (.A1(_3077_),
    .A2(_3071_),
    .A3(_1293_),
    .B1(_3080_),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _6559_ (.A1(\sub1.data_o[79] ),
    .A2(_2500_),
    .B1(_3072_),
    .B2(\sub1.data_o[15] ),
    .X(_3081_));
 sky130_fd_sc_hd__a31o_1 _6560_ (.A1(_3077_),
    .A2(_3071_),
    .A3(_1300_),
    .B1(_3081_),
    .X(_0263_));
 sky130_fd_sc_hd__nor2_2 _6561_ (.A(_0662_),
    .B(_0953_),
    .Y(_3082_));
 sky130_fd_sc_hd__mux2_1 _6562_ (.A0(\sub1.data_o[112] ),
    .A1(\sub1.data_o[48] ),
    .S(_1219_),
    .X(_3083_));
 sky130_fd_sc_hd__a22o_1 _6563_ (.A1(\sub1.data_o[16] ),
    .A2(_3082_),
    .B1(_3083_),
    .B2(\sub1.next_ready_o ),
    .X(_3084_));
 sky130_fd_sc_hd__a31o_1 _6564_ (.A1(_3077_),
    .A2(_0953_),
    .A3(_1213_),
    .B1(_3084_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _6565_ (.A0(\sub1.data_o[113] ),
    .A1(\sub1.data_o[49] ),
    .S(_1219_),
    .X(_3085_));
 sky130_fd_sc_hd__a22o_1 _6566_ (.A1(\sub1.data_o[17] ),
    .A2(_3082_),
    .B1(_3085_),
    .B2(\sub1.next_ready_o ),
    .X(_3086_));
 sky130_fd_sc_hd__a31o_1 _6567_ (.A1(_3077_),
    .A2(_0953_),
    .A3(_1247_),
    .B1(_3086_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _6568_ (.A0(\sub1.data_o[114] ),
    .A1(\sub1.data_o[50] ),
    .S(_1219_),
    .X(_3087_));
 sky130_fd_sc_hd__a22o_1 _6569_ (.A1(\sub1.data_o[18] ),
    .A2(_3082_),
    .B1(_3087_),
    .B2(\sub1.next_ready_o ),
    .X(_3088_));
 sky130_fd_sc_hd__a31o_1 _6570_ (.A1(_3077_),
    .A2(_0953_),
    .A3(_1257_),
    .B1(_3088_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _6571_ (.A0(\sub1.data_o[115] ),
    .A1(\sub1.data_o[51] ),
    .S(_1219_),
    .X(_3089_));
 sky130_fd_sc_hd__a22o_1 _6572_ (.A1(\sub1.data_o[19] ),
    .A2(_3082_),
    .B1(_3089_),
    .B2(\sub1.next_ready_o ),
    .X(_3090_));
 sky130_fd_sc_hd__a31o_1 _6573_ (.A1(_3077_),
    .A2(_0953_),
    .A3(_1272_),
    .B1(_3090_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _6574_ (.A0(\sub1.data_o[116] ),
    .A1(\sub1.data_o[52] ),
    .S(_1219_),
    .X(_3091_));
 sky130_fd_sc_hd__a22o_1 _6575_ (.A1(\sub1.data_o[20] ),
    .A2(_3082_),
    .B1(_3091_),
    .B2(\sub1.next_ready_o ),
    .X(_3092_));
 sky130_fd_sc_hd__a31o_1 _6576_ (.A1(_3077_),
    .A2(_0953_),
    .A3(_1278_),
    .B1(_3092_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _6577_ (.A0(\sub1.data_o[117] ),
    .A1(\sub1.data_o[53] ),
    .S(_1219_),
    .X(_3093_));
 sky130_fd_sc_hd__a22o_1 _6578_ (.A1(\sub1.data_o[21] ),
    .A2(_3082_),
    .B1(_3093_),
    .B2(\sub1.next_ready_o ),
    .X(_3094_));
 sky130_fd_sc_hd__a31o_1 _6579_ (.A1(_3077_),
    .A2(_0953_),
    .A3(_1286_),
    .B1(_3094_),
    .X(_0269_));
 sky130_fd_sc_hd__clkbuf_4 _6580_ (.A(_1139_),
    .X(_3095_));
 sky130_fd_sc_hd__mux2_1 _6581_ (.A0(\sub1.data_o[118] ),
    .A1(\sub1.data_o[54] ),
    .S(_1219_),
    .X(_3096_));
 sky130_fd_sc_hd__a22o_1 _6582_ (.A1(\sub1.data_o[22] ),
    .A2(_3082_),
    .B1(_3096_),
    .B2(\sub1.next_ready_o ),
    .X(_3097_));
 sky130_fd_sc_hd__a31o_1 _6583_ (.A1(_3095_),
    .A2(_0953_),
    .A3(_1293_),
    .B1(_3097_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _6584_ (.A0(\sub1.data_o[119] ),
    .A1(\sub1.data_o[55] ),
    .S(_1219_),
    .X(_3098_));
 sky130_fd_sc_hd__a22o_1 _6585_ (.A1(\sub1.data_o[23] ),
    .A2(_3082_),
    .B1(_3098_),
    .B2(\sub1.next_ready_o ),
    .X(_3099_));
 sky130_fd_sc_hd__a31o_1 _6586_ (.A1(_3095_),
    .A2(_0953_),
    .A3(_1300_),
    .B1(_3099_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _6587_ (.A0(\sub1.data_o[24] ),
    .A1(_1212_),
    .S(_0927_),
    .X(_3100_));
 sky130_fd_sc_hd__clkbuf_1 _6588_ (.A(_3100_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _6589_ (.A0(\sub1.data_o[25] ),
    .A1(_1246_),
    .S(_0927_),
    .X(_3101_));
 sky130_fd_sc_hd__clkbuf_1 _6590_ (.A(_3101_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _6591_ (.A0(\sub1.data_o[26] ),
    .A1(_1256_),
    .S(_0927_),
    .X(_3102_));
 sky130_fd_sc_hd__clkbuf_1 _6592_ (.A(_3102_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _6593_ (.A0(\sub1.data_o[27] ),
    .A1(_1271_),
    .S(_0927_),
    .X(_3103_));
 sky130_fd_sc_hd__clkbuf_1 _6594_ (.A(_3103_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _6595_ (.A0(\sub1.data_o[28] ),
    .A1(_1277_),
    .S(_0927_),
    .X(_3104_));
 sky130_fd_sc_hd__clkbuf_1 _6596_ (.A(_3104_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _6597_ (.A0(\sub1.data_o[29] ),
    .A1(_1285_),
    .S(_0927_),
    .X(_3105_));
 sky130_fd_sc_hd__clkbuf_1 _6598_ (.A(_3105_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _6599_ (.A0(\sub1.data_o[30] ),
    .A1(_1292_),
    .S(_0927_),
    .X(_3106_));
 sky130_fd_sc_hd__clkbuf_1 _6600_ (.A(_3106_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _6601_ (.A0(\sub1.data_o[31] ),
    .A1(_1299_),
    .S(_0927_),
    .X(_3107_));
 sky130_fd_sc_hd__clkbuf_1 _6602_ (.A(_3107_),
    .X(_0279_));
 sky130_fd_sc_hd__nand2_4 _6603_ (.A(_1214_),
    .B(_0661_),
    .Y(_3108_));
 sky130_fd_sc_hd__mux2_1 _6604_ (.A0(\sub1.data_o[64] ),
    .A1(_1212_),
    .S(_3108_),
    .X(_3109_));
 sky130_fd_sc_hd__or2_1 _6605_ (.A(_0661_),
    .B(_0713_),
    .X(_3110_));
 sky130_fd_sc_hd__clkbuf_4 _6606_ (.A(_3110_),
    .X(_3111_));
 sky130_fd_sc_hd__mux2_1 _6607_ (.A0(\sub1.data_o[32] ),
    .A1(_3109_),
    .S(_3111_),
    .X(_3112_));
 sky130_fd_sc_hd__clkbuf_1 _6608_ (.A(_3112_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _6609_ (.A0(\sub1.data_o[65] ),
    .A1(_1246_),
    .S(_3108_),
    .X(_3113_));
 sky130_fd_sc_hd__mux2_1 _6610_ (.A0(\sub1.data_o[33] ),
    .A1(_3113_),
    .S(_3111_),
    .X(_3114_));
 sky130_fd_sc_hd__clkbuf_1 _6611_ (.A(_3114_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _6612_ (.A0(\sub1.data_o[66] ),
    .A1(_1256_),
    .S(_3108_),
    .X(_3115_));
 sky130_fd_sc_hd__mux2_1 _6613_ (.A0(\sub1.data_o[34] ),
    .A1(_3115_),
    .S(_3111_),
    .X(_3116_));
 sky130_fd_sc_hd__clkbuf_1 _6614_ (.A(_3116_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _6615_ (.A0(\sub1.data_o[67] ),
    .A1(_1271_),
    .S(_3108_),
    .X(_3117_));
 sky130_fd_sc_hd__mux2_1 _6616_ (.A0(\sub1.data_o[35] ),
    .A1(_3117_),
    .S(_3111_),
    .X(_3118_));
 sky130_fd_sc_hd__clkbuf_1 _6617_ (.A(_3118_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _6618_ (.A0(\sub1.data_o[68] ),
    .A1(_1277_),
    .S(_3108_),
    .X(_3119_));
 sky130_fd_sc_hd__mux2_1 _6619_ (.A0(\sub1.data_o[36] ),
    .A1(_3119_),
    .S(_3111_),
    .X(_3120_));
 sky130_fd_sc_hd__clkbuf_1 _6620_ (.A(_3120_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _6621_ (.A0(\sub1.data_o[69] ),
    .A1(_1285_),
    .S(_3108_),
    .X(_3121_));
 sky130_fd_sc_hd__mux2_1 _6622_ (.A0(\sub1.data_o[37] ),
    .A1(_3121_),
    .S(_3111_),
    .X(_3122_));
 sky130_fd_sc_hd__clkbuf_1 _6623_ (.A(_3122_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _6624_ (.A0(\sub1.data_o[70] ),
    .A1(_1292_),
    .S(_3108_),
    .X(_3123_));
 sky130_fd_sc_hd__mux2_1 _6625_ (.A0(\sub1.data_o[38] ),
    .A1(_3123_),
    .S(_3111_),
    .X(_3124_));
 sky130_fd_sc_hd__clkbuf_1 _6626_ (.A(_3124_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _6627_ (.A0(\sub1.data_o[71] ),
    .A1(_1299_),
    .S(_3108_),
    .X(_3125_));
 sky130_fd_sc_hd__mux2_1 _6628_ (.A0(\sub1.data_o[39] ),
    .A1(_3125_),
    .S(_3111_),
    .X(_3126_));
 sky130_fd_sc_hd__clkbuf_1 _6629_ (.A(_3126_),
    .X(_0287_));
 sky130_fd_sc_hd__buf_2 _6630_ (.A(_0662_),
    .X(_3127_));
 sky130_fd_sc_hd__nor2_2 _6631_ (.A(_2491_),
    .B(_0967_),
    .Y(_3128_));
 sky130_fd_sc_hd__a22o_1 _6632_ (.A1(\sub1.data_o[104] ),
    .A2(_3127_),
    .B1(_3128_),
    .B2(\sub1.data_o[40] ),
    .X(_3129_));
 sky130_fd_sc_hd__a31o_1 _6633_ (.A1(_3095_),
    .A2(_0967_),
    .A3(_1213_),
    .B1(_3129_),
    .X(_0288_));
 sky130_fd_sc_hd__a22o_1 _6634_ (.A1(\sub1.data_o[105] ),
    .A2(_3127_),
    .B1(_3128_),
    .B2(\sub1.data_o[41] ),
    .X(_3130_));
 sky130_fd_sc_hd__a31o_1 _6635_ (.A1(_3095_),
    .A2(_0967_),
    .A3(_1247_),
    .B1(_3130_),
    .X(_0289_));
 sky130_fd_sc_hd__a22o_1 _6636_ (.A1(\sub1.data_o[106] ),
    .A2(_3127_),
    .B1(_3128_),
    .B2(\sub1.data_o[42] ),
    .X(_3131_));
 sky130_fd_sc_hd__a31o_1 _6637_ (.A1(_3095_),
    .A2(_0967_),
    .A3(_1257_),
    .B1(_3131_),
    .X(_0290_));
 sky130_fd_sc_hd__a22o_1 _6638_ (.A1(\sub1.data_o[107] ),
    .A2(_3127_),
    .B1(_3128_),
    .B2(\sub1.data_o[43] ),
    .X(_3132_));
 sky130_fd_sc_hd__a31o_1 _6639_ (.A1(_3095_),
    .A2(_0967_),
    .A3(_1272_),
    .B1(_3132_),
    .X(_0291_));
 sky130_fd_sc_hd__a22o_1 _6640_ (.A1(\sub1.data_o[108] ),
    .A2(_3127_),
    .B1(_3128_),
    .B2(\sub1.data_o[44] ),
    .X(_3133_));
 sky130_fd_sc_hd__a31o_1 _6641_ (.A1(_3095_),
    .A2(_0967_),
    .A3(_1278_),
    .B1(_3133_),
    .X(_0292_));
 sky130_fd_sc_hd__a22o_1 _6642_ (.A1(\sub1.data_o[109] ),
    .A2(_3127_),
    .B1(_3128_),
    .B2(\sub1.data_o[45] ),
    .X(_3134_));
 sky130_fd_sc_hd__a31o_1 _6643_ (.A1(_3095_),
    .A2(_0967_),
    .A3(_1286_),
    .B1(_3134_),
    .X(_0293_));
 sky130_fd_sc_hd__a22o_1 _6644_ (.A1(\sub1.data_o[110] ),
    .A2(_3127_),
    .B1(_3128_),
    .B2(\sub1.data_o[46] ),
    .X(_3135_));
 sky130_fd_sc_hd__a31o_1 _6645_ (.A1(_3095_),
    .A2(_0967_),
    .A3(_1293_),
    .B1(_3135_),
    .X(_0294_));
 sky130_fd_sc_hd__a22o_1 _6646_ (.A1(\sub1.data_o[111] ),
    .A2(_3127_),
    .B1(_3128_),
    .B2(\sub1.data_o[47] ),
    .X(_3136_));
 sky130_fd_sc_hd__a31o_1 _6647_ (.A1(_3095_),
    .A2(_0967_),
    .A3(_1300_),
    .B1(_3136_),
    .X(_0295_));
 sky130_fd_sc_hd__clkbuf_4 _6648_ (.A(_1139_),
    .X(_3137_));
 sky130_fd_sc_hd__nor2_2 _6649_ (.A(_0662_),
    .B(_0970_),
    .Y(_3138_));
 sky130_fd_sc_hd__buf_4 _6650_ (.A(_1218_),
    .X(_3139_));
 sky130_fd_sc_hd__mux2_1 _6651_ (.A0(\sub1.data_o[16] ),
    .A1(\sub1.data_o[80] ),
    .S(_3139_),
    .X(_3140_));
 sky130_fd_sc_hd__clkbuf_4 _6652_ (.A(_2491_),
    .X(_3141_));
 sky130_fd_sc_hd__a22o_1 _6653_ (.A1(\sub1.data_o[48] ),
    .A2(_3138_),
    .B1(_3140_),
    .B2(_3141_),
    .X(_3142_));
 sky130_fd_sc_hd__a31o_1 _6654_ (.A1(_3137_),
    .A2(_0970_),
    .A3(_1213_),
    .B1(_3142_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _6655_ (.A0(\sub1.data_o[17] ),
    .A1(\sub1.data_o[81] ),
    .S(_3139_),
    .X(_3143_));
 sky130_fd_sc_hd__a22o_1 _6656_ (.A1(\sub1.data_o[49] ),
    .A2(_3138_),
    .B1(_3143_),
    .B2(_3141_),
    .X(_3144_));
 sky130_fd_sc_hd__a31o_1 _6657_ (.A1(_3137_),
    .A2(_0970_),
    .A3(_1247_),
    .B1(_3144_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _6658_ (.A0(\sub1.data_o[18] ),
    .A1(\sub1.data_o[82] ),
    .S(_3139_),
    .X(_3145_));
 sky130_fd_sc_hd__a22o_1 _6659_ (.A1(\sub1.data_o[50] ),
    .A2(_3138_),
    .B1(_3145_),
    .B2(_3141_),
    .X(_3146_));
 sky130_fd_sc_hd__a31o_1 _6660_ (.A1(_3137_),
    .A2(_0970_),
    .A3(_1257_),
    .B1(_3146_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _6661_ (.A0(\sub1.data_o[19] ),
    .A1(\sub1.data_o[83] ),
    .S(_3139_),
    .X(_3147_));
 sky130_fd_sc_hd__a22o_1 _6662_ (.A1(\sub1.data_o[51] ),
    .A2(_3138_),
    .B1(_3147_),
    .B2(_3141_),
    .X(_3148_));
 sky130_fd_sc_hd__a31o_1 _6663_ (.A1(_3137_),
    .A2(_0970_),
    .A3(_1272_),
    .B1(_3148_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _6664_ (.A0(\sub1.data_o[20] ),
    .A1(\sub1.data_o[84] ),
    .S(_3139_),
    .X(_3149_));
 sky130_fd_sc_hd__a22o_1 _6665_ (.A1(\sub1.data_o[52] ),
    .A2(_3138_),
    .B1(_3149_),
    .B2(_3141_),
    .X(_3150_));
 sky130_fd_sc_hd__a31o_1 _6666_ (.A1(_3137_),
    .A2(_0970_),
    .A3(_1278_),
    .B1(_3150_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _6667_ (.A0(\sub1.data_o[21] ),
    .A1(\sub1.data_o[85] ),
    .S(_3139_),
    .X(_3151_));
 sky130_fd_sc_hd__a22o_1 _6668_ (.A1(\sub1.data_o[53] ),
    .A2(_3138_),
    .B1(_3151_),
    .B2(_3141_),
    .X(_3152_));
 sky130_fd_sc_hd__a31o_1 _6669_ (.A1(_3137_),
    .A2(_0970_),
    .A3(_1286_),
    .B1(_3152_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _6670_ (.A0(\sub1.data_o[22] ),
    .A1(\sub1.data_o[86] ),
    .S(_3139_),
    .X(_3153_));
 sky130_fd_sc_hd__a22o_1 _6671_ (.A1(\sub1.data_o[54] ),
    .A2(_3138_),
    .B1(_3153_),
    .B2(_3141_),
    .X(_3154_));
 sky130_fd_sc_hd__a31o_1 _6672_ (.A1(_3137_),
    .A2(_0970_),
    .A3(_1293_),
    .B1(_3154_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _6673_ (.A0(\sub1.data_o[23] ),
    .A1(\sub1.data_o[87] ),
    .S(_3139_),
    .X(_3155_));
 sky130_fd_sc_hd__a22o_1 _6674_ (.A1(\sub1.data_o[55] ),
    .A2(_3138_),
    .B1(_3155_),
    .B2(_3141_),
    .X(_3156_));
 sky130_fd_sc_hd__a31o_1 _6675_ (.A1(_3137_),
    .A2(_0970_),
    .A3(_1300_),
    .B1(_3156_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _6676_ (.A0(\sub1.data_o[56] ),
    .A1(_1212_),
    .S(_0929_),
    .X(_3157_));
 sky130_fd_sc_hd__clkbuf_1 _6677_ (.A(_3157_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _6678_ (.A0(\sub1.data_o[57] ),
    .A1(_1246_),
    .S(_0929_),
    .X(_3158_));
 sky130_fd_sc_hd__clkbuf_1 _6679_ (.A(_3158_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _6680_ (.A0(\sub1.data_o[58] ),
    .A1(_1256_),
    .S(_0929_),
    .X(_3159_));
 sky130_fd_sc_hd__clkbuf_1 _6681_ (.A(_3159_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _6682_ (.A0(\sub1.data_o[59] ),
    .A1(_1271_),
    .S(_0929_),
    .X(_3160_));
 sky130_fd_sc_hd__clkbuf_1 _6683_ (.A(_3160_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _6684_ (.A0(\sub1.data_o[60] ),
    .A1(_1277_),
    .S(_0929_),
    .X(_3161_));
 sky130_fd_sc_hd__clkbuf_1 _6685_ (.A(_3161_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _6686_ (.A0(\sub1.data_o[61] ),
    .A1(_1285_),
    .S(_0929_),
    .X(_3162_));
 sky130_fd_sc_hd__clkbuf_1 _6687_ (.A(_3162_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _6688_ (.A0(\sub1.data_o[62] ),
    .A1(_1292_),
    .S(_0929_),
    .X(_3163_));
 sky130_fd_sc_hd__clkbuf_1 _6689_ (.A(_3163_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _6690_ (.A0(\sub1.data_o[63] ),
    .A1(_1299_),
    .S(_0929_),
    .X(_3164_));
 sky130_fd_sc_hd__clkbuf_1 _6691_ (.A(_3164_),
    .X(_0311_));
 sky130_fd_sc_hd__nor2_2 _6692_ (.A(_0662_),
    .B(_0961_),
    .Y(_3165_));
 sky130_fd_sc_hd__mux2_1 _6693_ (.A0(\sub1.data_o[96] ),
    .A1(\sub1.data_o[32] ),
    .S(_3139_),
    .X(_3166_));
 sky130_fd_sc_hd__a22o_1 _6694_ (.A1(\sub1.data_o[64] ),
    .A2(_3165_),
    .B1(_3166_),
    .B2(_3141_),
    .X(_3167_));
 sky130_fd_sc_hd__a31o_1 _6695_ (.A1(_3137_),
    .A2(_0961_),
    .A3(_1213_),
    .B1(_3167_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _6696_ (.A0(\sub1.data_o[97] ),
    .A1(\sub1.data_o[33] ),
    .S(_3139_),
    .X(_3168_));
 sky130_fd_sc_hd__a22o_1 _6697_ (.A1(\sub1.data_o[65] ),
    .A2(_3165_),
    .B1(_3168_),
    .B2(_3141_),
    .X(_3169_));
 sky130_fd_sc_hd__a31o_1 _6698_ (.A1(_3137_),
    .A2(_0961_),
    .A3(_1247_),
    .B1(_3169_),
    .X(_0313_));
 sky130_fd_sc_hd__clkbuf_4 _6699_ (.A(_1139_),
    .X(_3170_));
 sky130_fd_sc_hd__buf_4 _6700_ (.A(_1218_),
    .X(_3171_));
 sky130_fd_sc_hd__mux2_1 _6701_ (.A0(\sub1.data_o[98] ),
    .A1(\sub1.data_o[34] ),
    .S(_3171_),
    .X(_3172_));
 sky130_fd_sc_hd__buf_2 _6702_ (.A(_2491_),
    .X(_3173_));
 sky130_fd_sc_hd__a22o_1 _6703_ (.A1(\sub1.data_o[66] ),
    .A2(_3165_),
    .B1(_3172_),
    .B2(_3173_),
    .X(_3174_));
 sky130_fd_sc_hd__a31o_1 _6704_ (.A1(_3170_),
    .A2(_0961_),
    .A3(_1257_),
    .B1(_3174_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _6705_ (.A0(\sub1.data_o[99] ),
    .A1(\sub1.data_o[35] ),
    .S(_3171_),
    .X(_3175_));
 sky130_fd_sc_hd__a22o_1 _6706_ (.A1(\sub1.data_o[67] ),
    .A2(_3165_),
    .B1(_3175_),
    .B2(_3173_),
    .X(_3176_));
 sky130_fd_sc_hd__a31o_1 _6707_ (.A1(_3170_),
    .A2(_0961_),
    .A3(_1272_),
    .B1(_3176_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _6708_ (.A0(\sub1.data_o[100] ),
    .A1(\sub1.data_o[36] ),
    .S(_3171_),
    .X(_3177_));
 sky130_fd_sc_hd__a22o_1 _6709_ (.A1(\sub1.data_o[68] ),
    .A2(_3165_),
    .B1(_3177_),
    .B2(_3173_),
    .X(_3178_));
 sky130_fd_sc_hd__a31o_1 _6710_ (.A1(_3170_),
    .A2(_0961_),
    .A3(_1278_),
    .B1(_3178_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _6711_ (.A0(\sub1.data_o[101] ),
    .A1(\sub1.data_o[37] ),
    .S(_3171_),
    .X(_3179_));
 sky130_fd_sc_hd__a22o_1 _6712_ (.A1(\sub1.data_o[69] ),
    .A2(_3165_),
    .B1(_3179_),
    .B2(_3173_),
    .X(_3180_));
 sky130_fd_sc_hd__a31o_1 _6713_ (.A1(_3170_),
    .A2(_0961_),
    .A3(_1286_),
    .B1(_3180_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _6714_ (.A0(\sub1.data_o[102] ),
    .A1(\sub1.data_o[38] ),
    .S(_3171_),
    .X(_3181_));
 sky130_fd_sc_hd__a22o_1 _6715_ (.A1(\sub1.data_o[70] ),
    .A2(_3165_),
    .B1(_3181_),
    .B2(_3173_),
    .X(_3182_));
 sky130_fd_sc_hd__a31o_1 _6716_ (.A1(_3170_),
    .A2(_0961_),
    .A3(_1293_),
    .B1(_3182_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _6717_ (.A0(\sub1.data_o[103] ),
    .A1(\sub1.data_o[39] ),
    .S(_3171_),
    .X(_3183_));
 sky130_fd_sc_hd__a22o_1 _6718_ (.A1(\sub1.data_o[71] ),
    .A2(_3165_),
    .B1(_3183_),
    .B2(_3173_),
    .X(_3184_));
 sky130_fd_sc_hd__a31o_1 _6719_ (.A1(_3170_),
    .A2(_0961_),
    .A3(_1300_),
    .B1(_3184_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _6720_ (.A0(\mix1.data_o[0] ),
    .A1(_2641_),
    .S(\mix1.next_ready_o ),
    .X(_3185_));
 sky130_fd_sc_hd__clkbuf_1 _6721_ (.A(_3185_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _6722_ (.A0(\mix1.data_o[1] ),
    .A1(_2709_),
    .S(\mix1.next_ready_o ),
    .X(_3186_));
 sky130_fd_sc_hd__clkbuf_1 _6723_ (.A(_3186_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _6724_ (.A0(\mix1.data_o[2] ),
    .A1(_2755_),
    .S(\mix1.next_ready_o ),
    .X(_3187_));
 sky130_fd_sc_hd__clkbuf_1 _6725_ (.A(_3187_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _6726_ (.A0(\mix1.data_o[3] ),
    .A1(_2796_),
    .S(\mix1.next_ready_o ),
    .X(_3188_));
 sky130_fd_sc_hd__clkbuf_1 _6727_ (.A(_3188_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _6728_ (.A0(\mix1.data_o[4] ),
    .A1(_2835_),
    .S(\mix1.next_ready_o ),
    .X(_3189_));
 sky130_fd_sc_hd__clkbuf_1 _6729_ (.A(_3189_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _6730_ (.A0(\mix1.data_o[5] ),
    .A1(_2854_),
    .S(\mix1.next_ready_o ),
    .X(_3190_));
 sky130_fd_sc_hd__clkbuf_1 _6731_ (.A(_3190_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _6732_ (.A0(\mix1.data_o[6] ),
    .A1(_2864_),
    .S(\mix1.next_ready_o ),
    .X(_3191_));
 sky130_fd_sc_hd__clkbuf_1 _6733_ (.A(_3191_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _6734_ (.A0(\mix1.data_o[7] ),
    .A1(_2874_),
    .S(\mix1.next_ready_o ),
    .X(_3192_));
 sky130_fd_sc_hd__clkbuf_1 _6735_ (.A(_3192_),
    .X(_0327_));
 sky130_fd_sc_hd__mux2_1 _6736_ (.A0(\mix1.data_o[8] ),
    .A1(_2883_),
    .S(\mix1.next_ready_o ),
    .X(_3193_));
 sky130_fd_sc_hd__clkbuf_1 _6737_ (.A(_3193_),
    .X(_0328_));
 sky130_fd_sc_hd__buf_4 _6738_ (.A(_0654_),
    .X(_3194_));
 sky130_fd_sc_hd__buf_4 _6739_ (.A(_3194_),
    .X(_3195_));
 sky130_fd_sc_hd__mux2_1 _6740_ (.A0(\mix1.data_o[9] ),
    .A1(_2896_),
    .S(_3195_),
    .X(_3196_));
 sky130_fd_sc_hd__clkbuf_1 _6741_ (.A(_3196_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _6742_ (.A0(\mix1.data_o[10] ),
    .A1(_2907_),
    .S(_3195_),
    .X(_3197_));
 sky130_fd_sc_hd__clkbuf_1 _6743_ (.A(_3197_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _6744_ (.A0(\mix1.data_o[11] ),
    .A1(_2918_),
    .S(_3195_),
    .X(_3198_));
 sky130_fd_sc_hd__clkbuf_1 _6745_ (.A(_3198_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _6746_ (.A0(\mix1.data_o[12] ),
    .A1(_2928_),
    .S(_3195_),
    .X(_3199_));
 sky130_fd_sc_hd__clkbuf_1 _6747_ (.A(_3199_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _6748_ (.A0(\mix1.data_o[13] ),
    .A1(_2939_),
    .S(_3195_),
    .X(_3200_));
 sky130_fd_sc_hd__clkbuf_1 _6749_ (.A(_3200_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _6750_ (.A0(\mix1.data_o[14] ),
    .A1(_2948_),
    .S(_3195_),
    .X(_3201_));
 sky130_fd_sc_hd__clkbuf_1 _6751_ (.A(_3201_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _6752_ (.A0(\mix1.data_o[15] ),
    .A1(_2954_),
    .S(_3195_),
    .X(_3202_));
 sky130_fd_sc_hd__clkbuf_1 _6753_ (.A(_3202_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _6754_ (.A0(\mix1.data_o[16] ),
    .A1(_2958_),
    .S(_3195_),
    .X(_3203_));
 sky130_fd_sc_hd__clkbuf_1 _6755_ (.A(_3203_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _6756_ (.A0(\mix1.data_o[17] ),
    .A1(_2962_),
    .S(_3195_),
    .X(_3204_));
 sky130_fd_sc_hd__clkbuf_1 _6757_ (.A(_3204_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _6758_ (.A0(\mix1.data_o[18] ),
    .A1(_2964_),
    .S(_3195_),
    .X(_3205_));
 sky130_fd_sc_hd__clkbuf_1 _6759_ (.A(_3205_),
    .X(_0338_));
 sky130_fd_sc_hd__buf_2 _6760_ (.A(_0654_),
    .X(_3206_));
 sky130_fd_sc_hd__buf_4 _6761_ (.A(_3206_),
    .X(_3207_));
 sky130_fd_sc_hd__mux2_1 _6762_ (.A0(\mix1.data_o[19] ),
    .A1(_2968_),
    .S(_3207_),
    .X(_3208_));
 sky130_fd_sc_hd__clkbuf_1 _6763_ (.A(_3208_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _6764_ (.A0(\mix1.data_o[20] ),
    .A1(_2973_),
    .S(_3207_),
    .X(_3209_));
 sky130_fd_sc_hd__clkbuf_1 _6765_ (.A(_3209_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _6766_ (.A0(\mix1.data_o[21] ),
    .A1(_2976_),
    .S(_3207_),
    .X(_3210_));
 sky130_fd_sc_hd__clkbuf_1 _6767_ (.A(_3210_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _6768_ (.A0(\mix1.data_o[22] ),
    .A1(_2978_),
    .S(_3207_),
    .X(_3211_));
 sky130_fd_sc_hd__clkbuf_1 _6769_ (.A(_3211_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _6770_ (.A0(\mix1.data_o[23] ),
    .A1(_2981_),
    .S(_3207_),
    .X(_3212_));
 sky130_fd_sc_hd__clkbuf_1 _6771_ (.A(_3212_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _6772_ (.A0(\mix1.data_o[24] ),
    .A1(_2985_),
    .S(_3207_),
    .X(_3213_));
 sky130_fd_sc_hd__clkbuf_1 _6773_ (.A(_3213_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _6774_ (.A0(\mix1.data_o[25] ),
    .A1(_2987_),
    .S(_3207_),
    .X(_3214_));
 sky130_fd_sc_hd__clkbuf_1 _6775_ (.A(_3214_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _6776_ (.A0(\mix1.data_o[26] ),
    .A1(_2992_),
    .S(_3207_),
    .X(_3215_));
 sky130_fd_sc_hd__clkbuf_1 _6777_ (.A(_3215_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _6778_ (.A0(\mix1.data_o[27] ),
    .A1(_2996_),
    .S(_3207_),
    .X(_3216_));
 sky130_fd_sc_hd__clkbuf_1 _6779_ (.A(_3216_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _6780_ (.A0(\mix1.data_o[28] ),
    .A1(_2998_),
    .S(_3207_),
    .X(_3217_));
 sky130_fd_sc_hd__clkbuf_1 _6781_ (.A(_3217_),
    .X(_0348_));
 sky130_fd_sc_hd__buf_4 _6782_ (.A(_3206_),
    .X(_3218_));
 sky130_fd_sc_hd__mux2_1 _6783_ (.A0(\mix1.data_o[29] ),
    .A1(_3000_),
    .S(_3218_),
    .X(_3219_));
 sky130_fd_sc_hd__clkbuf_1 _6784_ (.A(_3219_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _6785_ (.A0(\mix1.data_o[30] ),
    .A1(_3004_),
    .S(_3218_),
    .X(_3220_));
 sky130_fd_sc_hd__clkbuf_1 _6786_ (.A(_3220_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _6787_ (.A0(\mix1.data_o[31] ),
    .A1(_3008_),
    .S(_3218_),
    .X(_3221_));
 sky130_fd_sc_hd__clkbuf_1 _6788_ (.A(_3221_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _6789_ (.A0(\mix1.data_o[32] ),
    .A1(net608),
    .S(_3218_),
    .X(_3222_));
 sky130_fd_sc_hd__clkbuf_1 _6790_ (.A(_3222_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _6791_ (.A0(\mix1.data_o[33] ),
    .A1(net605),
    .S(_3218_),
    .X(_3223_));
 sky130_fd_sc_hd__clkbuf_1 _6792_ (.A(_3223_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _6793_ (.A0(\mix1.data_o[34] ),
    .A1(net559),
    .S(_3218_),
    .X(_3224_));
 sky130_fd_sc_hd__clkbuf_1 _6794_ (.A(_3224_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _6795_ (.A0(\mix1.data_o[35] ),
    .A1(net550),
    .S(_3218_),
    .X(_3225_));
 sky130_fd_sc_hd__clkbuf_1 _6796_ (.A(_3225_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _6797_ (.A0(\mix1.data_o[36] ),
    .A1(net587),
    .S(_3218_),
    .X(_3226_));
 sky130_fd_sc_hd__clkbuf_1 _6798_ (.A(_3226_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _6799_ (.A0(\mix1.data_o[37] ),
    .A1(net583),
    .S(_3218_),
    .X(_3227_));
 sky130_fd_sc_hd__clkbuf_1 _6800_ (.A(_3227_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _6801_ (.A0(\mix1.data_o[38] ),
    .A1(net544),
    .S(_3218_),
    .X(_3228_));
 sky130_fd_sc_hd__clkbuf_1 _6802_ (.A(_3228_),
    .X(_0358_));
 sky130_fd_sc_hd__buf_4 _6803_ (.A(_3206_),
    .X(_3229_));
 sky130_fd_sc_hd__mux2_1 _6804_ (.A0(\mix1.data_o[39] ),
    .A1(net577),
    .S(_3229_),
    .X(_3230_));
 sky130_fd_sc_hd__clkbuf_1 _6805_ (.A(_3230_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _6806_ (.A0(\mix1.data_o[40] ),
    .A1(net546),
    .S(_3229_),
    .X(_3231_));
 sky130_fd_sc_hd__clkbuf_1 _6807_ (.A(_3231_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _6808_ (.A0(\mix1.data_o[41] ),
    .A1(net531),
    .S(_3229_),
    .X(_3232_));
 sky130_fd_sc_hd__clkbuf_1 _6809_ (.A(_3232_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _6810_ (.A0(\mix1.data_o[42] ),
    .A1(net557),
    .S(_3229_),
    .X(_3233_));
 sky130_fd_sc_hd__clkbuf_1 _6811_ (.A(_3233_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _6812_ (.A0(\mix1.data_o[43] ),
    .A1(\mix1.data_reg[43] ),
    .S(_3229_),
    .X(_3234_));
 sky130_fd_sc_hd__clkbuf_1 _6813_ (.A(_3234_),
    .X(_0363_));
 sky130_fd_sc_hd__mux2_1 _6814_ (.A0(\mix1.data_o[44] ),
    .A1(net609),
    .S(_3229_),
    .X(_3235_));
 sky130_fd_sc_hd__clkbuf_1 _6815_ (.A(_3235_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _6816_ (.A0(\mix1.data_o[45] ),
    .A1(net533),
    .S(_3229_),
    .X(_3236_));
 sky130_fd_sc_hd__clkbuf_1 _6817_ (.A(_3236_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _6818_ (.A0(\mix1.data_o[46] ),
    .A1(net619),
    .S(_3229_),
    .X(_3237_));
 sky130_fd_sc_hd__clkbuf_1 _6819_ (.A(_3237_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _6820_ (.A0(\mix1.data_o[47] ),
    .A1(net618),
    .S(_3229_),
    .X(_3238_));
 sky130_fd_sc_hd__clkbuf_1 _6821_ (.A(_3238_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _6822_ (.A0(\mix1.data_o[48] ),
    .A1(net600),
    .S(_3229_),
    .X(_3239_));
 sky130_fd_sc_hd__clkbuf_1 _6823_ (.A(_3239_),
    .X(_0368_));
 sky130_fd_sc_hd__buf_4 _6824_ (.A(_3206_),
    .X(_3240_));
 sky130_fd_sc_hd__mux2_1 _6825_ (.A0(\mix1.data_o[49] ),
    .A1(net579),
    .S(_3240_),
    .X(_3241_));
 sky130_fd_sc_hd__clkbuf_1 _6826_ (.A(_3241_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _6827_ (.A0(\mix1.data_o[50] ),
    .A1(net594),
    .S(_3240_),
    .X(_3242_));
 sky130_fd_sc_hd__clkbuf_1 _6828_ (.A(_3242_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _6829_ (.A0(\mix1.data_o[51] ),
    .A1(net536),
    .S(_3240_),
    .X(_3243_));
 sky130_fd_sc_hd__clkbuf_1 _6830_ (.A(_3243_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _6831_ (.A0(\mix1.data_o[52] ),
    .A1(net573),
    .S(_3240_),
    .X(_3244_));
 sky130_fd_sc_hd__clkbuf_1 _6832_ (.A(_3244_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _6833_ (.A0(\mix1.data_o[53] ),
    .A1(net545),
    .S(_3240_),
    .X(_3245_));
 sky130_fd_sc_hd__clkbuf_1 _6834_ (.A(_3245_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _6835_ (.A0(\mix1.data_o[54] ),
    .A1(net589),
    .S(_3240_),
    .X(_3246_));
 sky130_fd_sc_hd__clkbuf_1 _6836_ (.A(_3246_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _6837_ (.A0(\mix1.data_o[55] ),
    .A1(net623),
    .S(_3240_),
    .X(_3247_));
 sky130_fd_sc_hd__clkbuf_1 _6838_ (.A(_3247_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _6839_ (.A0(\mix1.data_o[56] ),
    .A1(net552),
    .S(_3240_),
    .X(_3248_));
 sky130_fd_sc_hd__clkbuf_1 _6840_ (.A(_3248_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _6841_ (.A0(\mix1.data_o[57] ),
    .A1(net560),
    .S(_3240_),
    .X(_3249_));
 sky130_fd_sc_hd__clkbuf_1 _6842_ (.A(_3249_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _6843_ (.A0(\mix1.data_o[58] ),
    .A1(net558),
    .S(_3240_),
    .X(_3250_));
 sky130_fd_sc_hd__clkbuf_1 _6844_ (.A(_3250_),
    .X(_0378_));
 sky130_fd_sc_hd__buf_4 _6845_ (.A(_3206_),
    .X(_3251_));
 sky130_fd_sc_hd__mux2_1 _6846_ (.A0(\mix1.data_o[59] ),
    .A1(net530),
    .S(_3251_),
    .X(_3252_));
 sky130_fd_sc_hd__clkbuf_1 _6847_ (.A(_3252_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _6848_ (.A0(\mix1.data_o[60] ),
    .A1(net604),
    .S(_3251_),
    .X(_3253_));
 sky130_fd_sc_hd__clkbuf_1 _6849_ (.A(_3253_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _6850_ (.A0(\mix1.data_o[61] ),
    .A1(net603),
    .S(_3251_),
    .X(_3254_));
 sky130_fd_sc_hd__clkbuf_1 _6851_ (.A(_3254_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _6852_ (.A0(\mix1.data_o[62] ),
    .A1(net535),
    .S(_3251_),
    .X(_3255_));
 sky130_fd_sc_hd__clkbuf_1 _6853_ (.A(_3255_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _6854_ (.A0(\mix1.data_o[63] ),
    .A1(net599),
    .S(_3251_),
    .X(_3256_));
 sky130_fd_sc_hd__clkbuf_1 _6855_ (.A(_3256_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _6856_ (.A0(\mix1.data_o[64] ),
    .A1(net568),
    .S(_3251_),
    .X(_3257_));
 sky130_fd_sc_hd__clkbuf_1 _6857_ (.A(_3257_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _6858_ (.A0(\mix1.data_o[65] ),
    .A1(net584),
    .S(_3251_),
    .X(_3258_));
 sky130_fd_sc_hd__clkbuf_1 _6859_ (.A(_3258_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _6860_ (.A0(\mix1.data_o[66] ),
    .A1(net585),
    .S(_3251_),
    .X(_3259_));
 sky130_fd_sc_hd__clkbuf_1 _6861_ (.A(_3259_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _6862_ (.A0(\mix1.data_o[67] ),
    .A1(net521),
    .S(_3251_),
    .X(_3260_));
 sky130_fd_sc_hd__clkbuf_1 _6863_ (.A(_3260_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _6864_ (.A0(\mix1.data_o[68] ),
    .A1(net529),
    .S(_3251_),
    .X(_3261_));
 sky130_fd_sc_hd__clkbuf_1 _6865_ (.A(_3261_),
    .X(_0388_));
 sky130_fd_sc_hd__buf_4 _6866_ (.A(_3206_),
    .X(_3262_));
 sky130_fd_sc_hd__mux2_1 _6867_ (.A0(\mix1.data_o[69] ),
    .A1(net582),
    .S(_3262_),
    .X(_3263_));
 sky130_fd_sc_hd__clkbuf_1 _6868_ (.A(_3263_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _6869_ (.A0(\mix1.data_o[70] ),
    .A1(net566),
    .S(_3262_),
    .X(_3264_));
 sky130_fd_sc_hd__clkbuf_1 _6870_ (.A(_3264_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _6871_ (.A0(\mix1.data_o[71] ),
    .A1(net606),
    .S(_3262_),
    .X(_3265_));
 sky130_fd_sc_hd__clkbuf_1 _6872_ (.A(_3265_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _6873_ (.A0(\mix1.data_o[72] ),
    .A1(net596),
    .S(_3262_),
    .X(_3266_));
 sky130_fd_sc_hd__clkbuf_1 _6874_ (.A(_3266_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _6875_ (.A0(\mix1.data_o[73] ),
    .A1(net534),
    .S(_3262_),
    .X(_3267_));
 sky130_fd_sc_hd__clkbuf_1 _6876_ (.A(_3267_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _6877_ (.A0(\mix1.data_o[74] ),
    .A1(net555),
    .S(_3262_),
    .X(_3268_));
 sky130_fd_sc_hd__clkbuf_1 _6878_ (.A(_3268_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _6879_ (.A0(\mix1.data_o[75] ),
    .A1(net553),
    .S(_3262_),
    .X(_3269_));
 sky130_fd_sc_hd__clkbuf_1 _6880_ (.A(_3269_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _6881_ (.A0(\mix1.data_o[76] ),
    .A1(net532),
    .S(_3262_),
    .X(_3270_));
 sky130_fd_sc_hd__clkbuf_1 _6882_ (.A(_3270_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _6883_ (.A0(\mix1.data_o[77] ),
    .A1(net613),
    .S(_3262_),
    .X(_3271_));
 sky130_fd_sc_hd__clkbuf_1 _6884_ (.A(_3271_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _6885_ (.A0(\mix1.data_o[78] ),
    .A1(net602),
    .S(_3262_),
    .X(_3272_));
 sky130_fd_sc_hd__clkbuf_1 _6886_ (.A(_3272_),
    .X(_0398_));
 sky130_fd_sc_hd__buf_4 _6887_ (.A(_3206_),
    .X(_3273_));
 sky130_fd_sc_hd__mux2_1 _6888_ (.A0(\mix1.data_o[79] ),
    .A1(net597),
    .S(_3273_),
    .X(_3274_));
 sky130_fd_sc_hd__clkbuf_1 _6889_ (.A(_3274_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _6890_ (.A0(\mix1.data_o[80] ),
    .A1(net524),
    .S(_3273_),
    .X(_3275_));
 sky130_fd_sc_hd__clkbuf_1 _6891_ (.A(_3275_),
    .X(_0400_));
 sky130_fd_sc_hd__mux2_1 _6892_ (.A0(\mix1.data_o[81] ),
    .A1(net548),
    .S(_3273_),
    .X(_3276_));
 sky130_fd_sc_hd__clkbuf_1 _6893_ (.A(_3276_),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _6894_ (.A0(\mix1.data_o[82] ),
    .A1(net549),
    .S(_3273_),
    .X(_3277_));
 sky130_fd_sc_hd__clkbuf_1 _6895_ (.A(_3277_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _6896_ (.A0(\mix1.data_o[83] ),
    .A1(net572),
    .S(_3273_),
    .X(_3278_));
 sky130_fd_sc_hd__clkbuf_1 _6897_ (.A(_3278_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _6898_ (.A0(\mix1.data_o[84] ),
    .A1(net588),
    .S(_3273_),
    .X(_3279_));
 sky130_fd_sc_hd__clkbuf_1 _6899_ (.A(_3279_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2_1 _6900_ (.A0(\mix1.data_o[85] ),
    .A1(net525),
    .S(_3273_),
    .X(_3280_));
 sky130_fd_sc_hd__clkbuf_1 _6901_ (.A(_3280_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _6902_ (.A0(\mix1.data_o[86] ),
    .A1(net565),
    .S(_3273_),
    .X(_3281_));
 sky130_fd_sc_hd__clkbuf_1 _6903_ (.A(_3281_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _6904_ (.A0(\mix1.data_o[87] ),
    .A1(net611),
    .S(_3273_),
    .X(_3282_));
 sky130_fd_sc_hd__clkbuf_1 _6905_ (.A(_3282_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _6906_ (.A0(\mix1.data_o[88] ),
    .A1(net556),
    .S(_3273_),
    .X(_3283_));
 sky130_fd_sc_hd__clkbuf_1 _6907_ (.A(_3283_),
    .X(_0408_));
 sky130_fd_sc_hd__buf_4 _6908_ (.A(_3206_),
    .X(_3284_));
 sky130_fd_sc_hd__mux2_1 _6909_ (.A0(\mix1.data_o[89] ),
    .A1(\mix1.data_reg[89] ),
    .S(_3284_),
    .X(_3285_));
 sky130_fd_sc_hd__clkbuf_1 _6910_ (.A(_3285_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _6911_ (.A0(\mix1.data_o[90] ),
    .A1(net576),
    .S(_3284_),
    .X(_3286_));
 sky130_fd_sc_hd__clkbuf_1 _6912_ (.A(_3286_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _6913_ (.A0(\mix1.data_o[91] ),
    .A1(net601),
    .S(_3284_),
    .X(_3287_));
 sky130_fd_sc_hd__clkbuf_1 _6914_ (.A(_3287_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _6915_ (.A0(\mix1.data_o[92] ),
    .A1(net591),
    .S(_3284_),
    .X(_3288_));
 sky130_fd_sc_hd__clkbuf_1 _6916_ (.A(_3288_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _6917_ (.A0(\mix1.data_o[93] ),
    .A1(net527),
    .S(_3284_),
    .X(_3289_));
 sky130_fd_sc_hd__clkbuf_1 _6918_ (.A(_3289_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _6919_ (.A0(\mix1.data_o[94] ),
    .A1(net547),
    .S(_3284_),
    .X(_3290_));
 sky130_fd_sc_hd__clkbuf_1 _6920_ (.A(_3290_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _6921_ (.A0(\mix1.data_o[95] ),
    .A1(net554),
    .S(_3284_),
    .X(_3291_));
 sky130_fd_sc_hd__clkbuf_1 _6922_ (.A(_3291_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _6923_ (.A0(\mix1.data_o[96] ),
    .A1(net538),
    .S(_3284_),
    .X(_3292_));
 sky130_fd_sc_hd__clkbuf_1 _6924_ (.A(_3292_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _6925_ (.A0(\mix1.data_o[97] ),
    .A1(net542),
    .S(_3284_),
    .X(_3293_));
 sky130_fd_sc_hd__clkbuf_1 _6926_ (.A(_3293_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _6927_ (.A0(\mix1.data_o[98] ),
    .A1(net543),
    .S(_3284_),
    .X(_3294_));
 sky130_fd_sc_hd__clkbuf_1 _6928_ (.A(_3294_),
    .X(_0418_));
 sky130_fd_sc_hd__buf_4 _6929_ (.A(_3206_),
    .X(_3295_));
 sky130_fd_sc_hd__mux2_1 _6930_ (.A0(\mix1.data_o[99] ),
    .A1(net541),
    .S(_3295_),
    .X(_3296_));
 sky130_fd_sc_hd__clkbuf_1 _6931_ (.A(_3296_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _6932_ (.A0(\mix1.data_o[100] ),
    .A1(net562),
    .S(_3295_),
    .X(_3297_));
 sky130_fd_sc_hd__clkbuf_1 _6933_ (.A(_3297_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _6934_ (.A0(\mix1.data_o[101] ),
    .A1(net561),
    .S(_3295_),
    .X(_3298_));
 sky130_fd_sc_hd__clkbuf_1 _6935_ (.A(_3298_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_1 _6936_ (.A0(\mix1.data_o[102] ),
    .A1(net551),
    .S(_3295_),
    .X(_3299_));
 sky130_fd_sc_hd__clkbuf_1 _6937_ (.A(_3299_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _6938_ (.A0(\mix1.data_o[103] ),
    .A1(net563),
    .S(_3295_),
    .X(_3300_));
 sky130_fd_sc_hd__clkbuf_1 _6939_ (.A(_3300_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _6940_ (.A0(\mix1.data_o[104] ),
    .A1(net539),
    .S(_3295_),
    .X(_3301_));
 sky130_fd_sc_hd__clkbuf_1 _6941_ (.A(_3301_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _6942_ (.A0(\mix1.data_o[105] ),
    .A1(net537),
    .S(_3295_),
    .X(_3302_));
 sky130_fd_sc_hd__clkbuf_1 _6943_ (.A(_3302_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _6944_ (.A0(\mix1.data_o[106] ),
    .A1(net564),
    .S(_3295_),
    .X(_3303_));
 sky130_fd_sc_hd__clkbuf_1 _6945_ (.A(_3303_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _6946_ (.A0(\mix1.data_o[107] ),
    .A1(net574),
    .S(_3295_),
    .X(_3304_));
 sky130_fd_sc_hd__clkbuf_1 _6947_ (.A(_3304_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _6948_ (.A0(\mix1.data_o[108] ),
    .A1(net598),
    .S(_3295_),
    .X(_3305_));
 sky130_fd_sc_hd__clkbuf_1 _6949_ (.A(_3305_),
    .X(_0428_));
 sky130_fd_sc_hd__buf_4 _6950_ (.A(_3206_),
    .X(_3306_));
 sky130_fd_sc_hd__mux2_1 _6951_ (.A0(\mix1.data_o[109] ),
    .A1(net590),
    .S(_3306_),
    .X(_3307_));
 sky130_fd_sc_hd__clkbuf_1 _6952_ (.A(_3307_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _6953_ (.A0(\mix1.data_o[110] ),
    .A1(net701),
    .S(_3306_),
    .X(_3308_));
 sky130_fd_sc_hd__clkbuf_1 _6954_ (.A(_3308_),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_1 _6955_ (.A0(\mix1.data_o[111] ),
    .A1(net627),
    .S(_3306_),
    .X(_3309_));
 sky130_fd_sc_hd__clkbuf_1 _6956_ (.A(_3309_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _6957_ (.A0(\mix1.data_o[112] ),
    .A1(net569),
    .S(_3306_),
    .X(_3310_));
 sky130_fd_sc_hd__clkbuf_1 _6958_ (.A(_3310_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _6959_ (.A0(\mix1.data_o[113] ),
    .A1(net571),
    .S(_3306_),
    .X(_3311_));
 sky130_fd_sc_hd__clkbuf_1 _6960_ (.A(_3311_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _6961_ (.A0(\mix1.data_o[114] ),
    .A1(\mix1.data_reg[114] ),
    .S(_3306_),
    .X(_3312_));
 sky130_fd_sc_hd__clkbuf_1 _6962_ (.A(_3312_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _6963_ (.A0(\mix1.data_o[115] ),
    .A1(net622),
    .S(_3306_),
    .X(_3313_));
 sky130_fd_sc_hd__clkbuf_1 _6964_ (.A(_3313_),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _6965_ (.A0(\mix1.data_o[116] ),
    .A1(net570),
    .S(_3306_),
    .X(_3314_));
 sky130_fd_sc_hd__clkbuf_1 _6966_ (.A(_3314_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _6967_ (.A0(\mix1.data_o[117] ),
    .A1(net526),
    .S(_3306_),
    .X(_3315_));
 sky130_fd_sc_hd__clkbuf_1 _6968_ (.A(_3315_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _6969_ (.A0(\mix1.data_o[118] ),
    .A1(net610),
    .S(_3306_),
    .X(_3316_));
 sky130_fd_sc_hd__clkbuf_1 _6970_ (.A(_3316_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _6971_ (.A0(\mix1.data_o[119] ),
    .A1(net616),
    .S(_3194_),
    .X(_3317_));
 sky130_fd_sc_hd__clkbuf_1 _6972_ (.A(_3317_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _6973_ (.A0(\mix1.data_o[120] ),
    .A1(net575),
    .S(_3194_),
    .X(_3318_));
 sky130_fd_sc_hd__clkbuf_1 _6974_ (.A(_3318_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _6975_ (.A0(\mix1.data_o[121] ),
    .A1(net595),
    .S(_3194_),
    .X(_3319_));
 sky130_fd_sc_hd__clkbuf_1 _6976_ (.A(_3319_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _6977_ (.A0(\mix1.data_o[122] ),
    .A1(net580),
    .S(_3194_),
    .X(_3320_));
 sky130_fd_sc_hd__clkbuf_1 _6978_ (.A(_3320_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _6979_ (.A0(\mix1.data_o[123] ),
    .A1(net567),
    .S(_3194_),
    .X(_3321_));
 sky130_fd_sc_hd__clkbuf_1 _6980_ (.A(_3321_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _6981_ (.A0(\mix1.data_o[124] ),
    .A1(net593),
    .S(_3194_),
    .X(_3322_));
 sky130_fd_sc_hd__clkbuf_1 _6982_ (.A(_3322_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _6983_ (.A0(\mix1.data_o[125] ),
    .A1(net586),
    .S(_3194_),
    .X(_3323_));
 sky130_fd_sc_hd__clkbuf_1 _6984_ (.A(_3323_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _6985_ (.A0(\mix1.data_o[126] ),
    .A1(net540),
    .S(_3194_),
    .X(_3324_));
 sky130_fd_sc_hd__clkbuf_1 _6986_ (.A(_3324_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _6987_ (.A0(\mix1.data_o[127] ),
    .A1(net581),
    .S(_3194_),
    .X(_3325_));
 sky130_fd_sc_hd__clkbuf_1 _6988_ (.A(_3325_),
    .X(_0447_));
 sky130_fd_sc_hd__inv_2 _6989_ (.A(_0719_),
    .Y(_3326_));
 sky130_fd_sc_hd__a211oi_1 _6990_ (.A1(_3326_),
    .A2(_0720_),
    .B1(_0655_),
    .C1(\sub1.next_ready_o ),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_1 _6991_ (.A(_0691_),
    .B(_0705_),
    .Y(_0449_));
 sky130_fd_sc_hd__xnor2_1 _6992_ (.A(\sub1.state[2] ),
    .B(_0686_),
    .Y(_0450_));
 sky130_fd_sc_hd__o21a_1 _6993_ (.A1(_0699_),
    .A2(_0686_),
    .B1(_0657_),
    .X(_3327_));
 sky130_fd_sc_hd__or2_1 _6994_ (.A(_2489_),
    .B(_3327_),
    .X(_3328_));
 sky130_fd_sc_hd__clkbuf_1 _6995_ (.A(_3328_),
    .X(_0451_));
 sky130_fd_sc_hd__o21ai_1 _6996_ (.A1(net497),
    .A2(_3071_),
    .B1(_0658_),
    .Y(_3329_));
 sky130_fd_sc_hd__a21oi_1 _6997_ (.A1(net497),
    .A2(_3071_),
    .B1(_3329_),
    .Y(_0452_));
 sky130_fd_sc_hd__nor2_2 _6998_ (.A(_0662_),
    .B(_0947_),
    .Y(_3330_));
 sky130_fd_sc_hd__mux2_1 _6999_ (.A0(\sub1.data_o[48] ),
    .A1(\sub1.data_o[112] ),
    .S(_3171_),
    .X(_3331_));
 sky130_fd_sc_hd__a22o_1 _7000_ (.A1(\sub1.data_o[80] ),
    .A2(_3330_),
    .B1(_3331_),
    .B2(_3173_),
    .X(_3332_));
 sky130_fd_sc_hd__a31o_1 _7001_ (.A1(_3170_),
    .A2(_0947_),
    .A3(_1213_),
    .B1(_3332_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _7002_ (.A0(\sub1.data_o[49] ),
    .A1(\sub1.data_o[113] ),
    .S(_3171_),
    .X(_3333_));
 sky130_fd_sc_hd__a22o_1 _7003_ (.A1(\sub1.data_o[81] ),
    .A2(_3330_),
    .B1(_3333_),
    .B2(_3173_),
    .X(_3334_));
 sky130_fd_sc_hd__a31o_1 _7004_ (.A1(_3170_),
    .A2(_0947_),
    .A3(_1247_),
    .B1(_3334_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _7005_ (.A0(\sub1.data_o[50] ),
    .A1(\sub1.data_o[114] ),
    .S(_3171_),
    .X(_3335_));
 sky130_fd_sc_hd__a22o_1 _7006_ (.A1(\sub1.data_o[82] ),
    .A2(_3330_),
    .B1(_3335_),
    .B2(_3173_),
    .X(_3336_));
 sky130_fd_sc_hd__a31o_1 _7007_ (.A1(_3170_),
    .A2(_0947_),
    .A3(_1257_),
    .B1(_3336_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _7008_ (.A0(\sub1.data_o[51] ),
    .A1(\sub1.data_o[115] ),
    .S(_3171_),
    .X(_3337_));
 sky130_fd_sc_hd__a22o_1 _7009_ (.A1(\sub1.data_o[83] ),
    .A2(_3330_),
    .B1(_3337_),
    .B2(_3173_),
    .X(_3338_));
 sky130_fd_sc_hd__a31o_1 _7010_ (.A1(_3170_),
    .A2(_0947_),
    .A3(_1272_),
    .B1(_3338_),
    .X(_0456_));
 sky130_fd_sc_hd__clkbuf_4 _7011_ (.A(_1139_),
    .X(_3339_));
 sky130_fd_sc_hd__mux2_1 _7012_ (.A0(\sub1.data_o[52] ),
    .A1(\sub1.data_o[116] ),
    .S(_3053_),
    .X(_3340_));
 sky130_fd_sc_hd__a22o_1 _7013_ (.A1(\sub1.data_o[84] ),
    .A2(_3330_),
    .B1(_3340_),
    .B2(_2490_),
    .X(_3341_));
 sky130_fd_sc_hd__a31o_1 _7014_ (.A1(_3339_),
    .A2(_0947_),
    .A3(_1278_),
    .B1(_3341_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _7015_ (.A0(\sub1.data_o[53] ),
    .A1(\sub1.data_o[117] ),
    .S(_3053_),
    .X(_3342_));
 sky130_fd_sc_hd__a22o_1 _7016_ (.A1(\sub1.data_o[85] ),
    .A2(_3330_),
    .B1(_3342_),
    .B2(_2490_),
    .X(_3343_));
 sky130_fd_sc_hd__a31o_1 _7017_ (.A1(_3339_),
    .A2(_0947_),
    .A3(_1286_),
    .B1(_3343_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _7018_ (.A0(\sub1.data_o[54] ),
    .A1(\sub1.data_o[118] ),
    .S(_3053_),
    .X(_3344_));
 sky130_fd_sc_hd__a22o_1 _7019_ (.A1(\sub1.data_o[86] ),
    .A2(_3330_),
    .B1(_3344_),
    .B2(_2490_),
    .X(_3345_));
 sky130_fd_sc_hd__a31o_1 _7020_ (.A1(_3339_),
    .A2(_0947_),
    .A3(_1293_),
    .B1(_3345_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _7021_ (.A0(\sub1.data_o[55] ),
    .A1(\sub1.data_o[119] ),
    .S(_3053_),
    .X(_3346_));
 sky130_fd_sc_hd__a22o_1 _7022_ (.A1(\sub1.data_o[87] ),
    .A2(_3330_),
    .B1(_3346_),
    .B2(_2490_),
    .X(_3347_));
 sky130_fd_sc_hd__a31o_1 _7023_ (.A1(_3339_),
    .A2(_0947_),
    .A3(_1300_),
    .B1(_3347_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _7024_ (.A0(\sub1.data_o[88] ),
    .A1(_1212_),
    .S(_0903_),
    .X(_3348_));
 sky130_fd_sc_hd__clkbuf_1 _7025_ (.A(_3348_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _7026_ (.A0(\sub1.data_o[89] ),
    .A1(_1246_),
    .S(_0903_),
    .X(_3349_));
 sky130_fd_sc_hd__clkbuf_1 _7027_ (.A(_3349_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _7028_ (.A0(\sub1.data_o[90] ),
    .A1(_1256_),
    .S(_0903_),
    .X(_3350_));
 sky130_fd_sc_hd__clkbuf_1 _7029_ (.A(_3350_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _7030_ (.A0(\sub1.data_o[91] ),
    .A1(_1271_),
    .S(_0903_),
    .X(_3351_));
 sky130_fd_sc_hd__clkbuf_1 _7031_ (.A(_3351_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _7032_ (.A0(\sub1.data_o[92] ),
    .A1(_1277_),
    .S(_0903_),
    .X(_3352_));
 sky130_fd_sc_hd__clkbuf_1 _7033_ (.A(_3352_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _7034_ (.A0(\sub1.data_o[93] ),
    .A1(_1285_),
    .S(_0903_),
    .X(_3353_));
 sky130_fd_sc_hd__clkbuf_1 _7035_ (.A(_3353_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _7036_ (.A0(\sub1.data_o[94] ),
    .A1(_1292_),
    .S(_0903_),
    .X(_3354_));
 sky130_fd_sc_hd__clkbuf_1 _7037_ (.A(_3354_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _7038_ (.A0(\sub1.data_o[95] ),
    .A1(_1299_),
    .S(_0903_),
    .X(_3355_));
 sky130_fd_sc_hd__clkbuf_1 _7039_ (.A(_3355_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _7040_ (.A0(_1212_),
    .A1(\sub1.data_o[64] ),
    .S(_1216_),
    .X(_3356_));
 sky130_fd_sc_hd__or2_1 _7041_ (.A(_0661_),
    .B(_0727_),
    .X(_3357_));
 sky130_fd_sc_hd__clkbuf_4 _7042_ (.A(_3357_),
    .X(_3358_));
 sky130_fd_sc_hd__mux2_1 _7043_ (.A0(\sub1.data_o[96] ),
    .A1(_3356_),
    .S(_3358_),
    .X(_3359_));
 sky130_fd_sc_hd__clkbuf_1 _7044_ (.A(_3359_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _7045_ (.A0(_1246_),
    .A1(\sub1.data_o[65] ),
    .S(_1216_),
    .X(_3360_));
 sky130_fd_sc_hd__mux2_1 _7046_ (.A0(\sub1.data_o[97] ),
    .A1(_3360_),
    .S(_3358_),
    .X(_3361_));
 sky130_fd_sc_hd__clkbuf_1 _7047_ (.A(_3361_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _7048_ (.A0(_1256_),
    .A1(\sub1.data_o[66] ),
    .S(_1215_),
    .X(_3362_));
 sky130_fd_sc_hd__mux2_1 _7049_ (.A0(\sub1.data_o[98] ),
    .A1(_3362_),
    .S(_3358_),
    .X(_3363_));
 sky130_fd_sc_hd__clkbuf_1 _7050_ (.A(_3363_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _7051_ (.A0(_1271_),
    .A1(\sub1.data_o[67] ),
    .S(_1215_),
    .X(_3364_));
 sky130_fd_sc_hd__mux2_1 _7052_ (.A0(\sub1.data_o[99] ),
    .A1(_3364_),
    .S(_3358_),
    .X(_3365_));
 sky130_fd_sc_hd__clkbuf_1 _7053_ (.A(_3365_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _7054_ (.A0(_1277_),
    .A1(\sub1.data_o[68] ),
    .S(_1215_),
    .X(_3366_));
 sky130_fd_sc_hd__mux2_1 _7055_ (.A0(\sub1.data_o[100] ),
    .A1(_3366_),
    .S(_3358_),
    .X(_3367_));
 sky130_fd_sc_hd__clkbuf_1 _7056_ (.A(_3367_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _7057_ (.A0(_1285_),
    .A1(\sub1.data_o[69] ),
    .S(_1215_),
    .X(_3368_));
 sky130_fd_sc_hd__mux2_1 _7058_ (.A0(\sub1.data_o[101] ),
    .A1(_3368_),
    .S(_3358_),
    .X(_3369_));
 sky130_fd_sc_hd__clkbuf_1 _7059_ (.A(_3369_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _7060_ (.A0(_1292_),
    .A1(\sub1.data_o[70] ),
    .S(_1215_),
    .X(_3370_));
 sky130_fd_sc_hd__mux2_1 _7061_ (.A0(\sub1.data_o[102] ),
    .A1(_3370_),
    .S(_3358_),
    .X(_3371_));
 sky130_fd_sc_hd__clkbuf_1 _7062_ (.A(_3371_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _7063_ (.A0(_1299_),
    .A1(\sub1.data_o[71] ),
    .S(_1215_),
    .X(_3372_));
 sky130_fd_sc_hd__mux2_1 _7064_ (.A0(\sub1.data_o[103] ),
    .A1(_3372_),
    .S(_3358_),
    .X(_3373_));
 sky130_fd_sc_hd__clkbuf_1 _7065_ (.A(_3373_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_4 _7066_ (.A(_0754_),
    .X(_3374_));
 sky130_fd_sc_hd__clkbuf_4 _7067_ (.A(_3374_),
    .X(_3375_));
 sky130_fd_sc_hd__buf_4 _7068_ (.A(_0810_),
    .X(_3376_));
 sky130_fd_sc_hd__clkbuf_8 _7069_ (.A(_3376_),
    .X(_3377_));
 sky130_fd_sc_hd__mux2_2 _7070_ (.A0(\ks1.key_reg[96] ),
    .A1(net253),
    .S(_3377_),
    .X(_3378_));
 sky130_fd_sc_hd__xor2_4 _7071_ (.A(\ks1.col[0] ),
    .B(_3378_),
    .X(_3379_));
 sky130_fd_sc_hd__buf_6 _7072_ (.A(_0810_),
    .X(_3380_));
 sky130_fd_sc_hd__clkbuf_8 _7073_ (.A(_3380_),
    .X(_3381_));
 sky130_fd_sc_hd__clkbuf_8 _7074_ (.A(_3381_),
    .X(_3382_));
 sky130_fd_sc_hd__mux2_1 _7075_ (.A0(\ks1.key_reg[64] ),
    .A1(net218),
    .S(_3382_),
    .X(_3383_));
 sky130_fd_sc_hd__xor2_2 _7076_ (.A(_3379_),
    .B(_3383_),
    .X(_3384_));
 sky130_fd_sc_hd__buf_4 _7077_ (.A(_3381_),
    .X(_3385_));
 sky130_fd_sc_hd__buf_4 _7078_ (.A(_3385_),
    .X(_3386_));
 sky130_fd_sc_hd__mux2_1 _7079_ (.A0(\ks1.key_reg[32] ),
    .A1(net183),
    .S(_3386_),
    .X(_3387_));
 sky130_fd_sc_hd__xor2_2 _7080_ (.A(_3384_),
    .B(_3387_),
    .X(_3388_));
 sky130_fd_sc_hd__or2_1 _7081_ (.A(_0934_),
    .B(_3388_),
    .X(_3389_));
 sky130_fd_sc_hd__clkbuf_4 _7082_ (.A(_0754_),
    .X(_3390_));
 sky130_fd_sc_hd__a21oi_1 _7083_ (.A1(_0934_),
    .A2(_3388_),
    .B1(_3390_),
    .Y(_3391_));
 sky130_fd_sc_hd__a22o_1 _7084_ (.A1(net512),
    .A2(_3375_),
    .B1(_3389_),
    .B2(_3391_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_2 _7085_ (.A0(\ks1.key_reg[97] ),
    .A1(net254),
    .S(_3377_),
    .X(_3392_));
 sky130_fd_sc_hd__xor2_4 _7086_ (.A(\ks1.col[1] ),
    .B(_3392_),
    .X(_3393_));
 sky130_fd_sc_hd__mux2_1 _7087_ (.A0(\ks1.key_reg[65] ),
    .A1(net219),
    .S(_3382_),
    .X(_3394_));
 sky130_fd_sc_hd__xor2_2 _7088_ (.A(_3393_),
    .B(_3394_),
    .X(_3395_));
 sky130_fd_sc_hd__mux2_1 _7089_ (.A0(\ks1.key_reg[33] ),
    .A1(net184),
    .S(_3386_),
    .X(_3396_));
 sky130_fd_sc_hd__xor2_2 _7090_ (.A(_3395_),
    .B(_3396_),
    .X(_3397_));
 sky130_fd_sc_hd__or2_1 _7091_ (.A(_0768_),
    .B(_3397_),
    .X(_3398_));
 sky130_fd_sc_hd__clkbuf_4 _7092_ (.A(_0754_),
    .X(_3399_));
 sky130_fd_sc_hd__a21oi_1 _7093_ (.A1(_0768_),
    .A2(_3397_),
    .B1(_3399_),
    .Y(_3400_));
 sky130_fd_sc_hd__a22o_1 _7094_ (.A1(net518),
    .A2(_3375_),
    .B1(_3398_),
    .B2(_3400_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_2 _7095_ (.A0(\ks1.key_reg[98] ),
    .A1(net255),
    .S(_3377_),
    .X(_3401_));
 sky130_fd_sc_hd__xor2_4 _7096_ (.A(\ks1.col[2] ),
    .B(_3401_),
    .X(_3402_));
 sky130_fd_sc_hd__mux2_1 _7097_ (.A0(\ks1.key_reg[66] ),
    .A1(net220),
    .S(_3382_),
    .X(_3403_));
 sky130_fd_sc_hd__xor2_2 _7098_ (.A(_3402_),
    .B(_3403_),
    .X(_3404_));
 sky130_fd_sc_hd__mux2_1 _7099_ (.A0(\ks1.key_reg[34] ),
    .A1(net185),
    .S(_3386_),
    .X(_3405_));
 sky130_fd_sc_hd__xor2_1 _7100_ (.A(_3404_),
    .B(_3405_),
    .X(_3406_));
 sky130_fd_sc_hd__or2_1 _7101_ (.A(_1057_),
    .B(_3406_),
    .X(_3407_));
 sky130_fd_sc_hd__a21oi_1 _7102_ (.A1(_1057_),
    .A2(_3406_),
    .B1(_3399_),
    .Y(_3408_));
 sky130_fd_sc_hd__a22o_1 _7103_ (.A1(net522),
    .A2(_3375_),
    .B1(_3407_),
    .B2(_3408_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _7104_ (.A0(\ks1.key_reg[99] ),
    .A1(net256),
    .S(_3377_),
    .X(_3409_));
 sky130_fd_sc_hd__xor2_2 _7105_ (.A(\ks1.col[3] ),
    .B(_3409_),
    .X(_3410_));
 sky130_fd_sc_hd__mux2_1 _7106_ (.A0(\ks1.key_reg[67] ),
    .A1(net221),
    .S(_3382_),
    .X(_3411_));
 sky130_fd_sc_hd__xor2_1 _7107_ (.A(_3410_),
    .B(_3411_),
    .X(_3412_));
 sky130_fd_sc_hd__mux2_1 _7108_ (.A0(\ks1.key_reg[35] ),
    .A1(net186),
    .S(_3386_),
    .X(_3413_));
 sky130_fd_sc_hd__xor2_1 _7109_ (.A(_3412_),
    .B(_3413_),
    .X(_3414_));
 sky130_fd_sc_hd__or2_1 _7110_ (.A(_0853_),
    .B(_3414_),
    .X(_3415_));
 sky130_fd_sc_hd__a21oi_1 _7111_ (.A1(_0853_),
    .A2(_3414_),
    .B1(_3399_),
    .Y(_3416_));
 sky130_fd_sc_hd__a22o_1 _7112_ (.A1(net502),
    .A2(_3375_),
    .B1(_3415_),
    .B2(_3416_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _7113_ (.A0(\ks1.key_reg[100] ),
    .A1(net131),
    .S(_3377_),
    .X(_3417_));
 sky130_fd_sc_hd__xor2_2 _7114_ (.A(\ks1.col[4] ),
    .B(_3417_),
    .X(_3418_));
 sky130_fd_sc_hd__clkbuf_8 _7115_ (.A(_3381_),
    .X(_3419_));
 sky130_fd_sc_hd__mux2_1 _7116_ (.A0(\ks1.key_reg[68] ),
    .A1(net222),
    .S(_3419_),
    .X(_3420_));
 sky130_fd_sc_hd__xor2_2 _7117_ (.A(_3418_),
    .B(_3420_),
    .X(_3421_));
 sky130_fd_sc_hd__mux2_1 _7118_ (.A0(\ks1.key_reg[36] ),
    .A1(net187),
    .S(_3386_),
    .X(_3422_));
 sky130_fd_sc_hd__xor2_2 _7119_ (.A(_3421_),
    .B(_3422_),
    .X(_3423_));
 sky130_fd_sc_hd__or2_1 _7120_ (.A(_0890_),
    .B(_3423_),
    .X(_3424_));
 sky130_fd_sc_hd__a21oi_1 _7121_ (.A1(_0890_),
    .A2(_3423_),
    .B1(_3399_),
    .Y(_3425_));
 sky130_fd_sc_hd__a22o_1 _7122_ (.A1(net516),
    .A2(_3375_),
    .B1(_3424_),
    .B2(_3425_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _7123_ (.A0(\ks1.key_reg[101] ),
    .A1(net132),
    .S(_3377_),
    .X(_3426_));
 sky130_fd_sc_hd__xor2_2 _7124_ (.A(\ks1.col[5] ),
    .B(_3426_),
    .X(_3427_));
 sky130_fd_sc_hd__mux2_1 _7125_ (.A0(\ks1.key_reg[69] ),
    .A1(net223),
    .S(_3419_),
    .X(_3428_));
 sky130_fd_sc_hd__xor2_2 _7126_ (.A(_3427_),
    .B(_3428_),
    .X(_3429_));
 sky130_fd_sc_hd__mux2_1 _7127_ (.A0(\ks1.key_reg[37] ),
    .A1(net188),
    .S(_3386_),
    .X(_3430_));
 sky130_fd_sc_hd__xor2_2 _7128_ (.A(_3429_),
    .B(_3430_),
    .X(_3431_));
 sky130_fd_sc_hd__or2_1 _7129_ (.A(_0977_),
    .B(_3431_),
    .X(_3432_));
 sky130_fd_sc_hd__a21oi_1 _7130_ (.A1(_0977_),
    .A2(_3431_),
    .B1(_3399_),
    .Y(_3433_));
 sky130_fd_sc_hd__a22o_1 _7131_ (.A1(net511),
    .A2(_3375_),
    .B1(_3432_),
    .B2(_3433_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_2 _7132_ (.A0(\ks1.key_reg[102] ),
    .A1(net133),
    .S(_3377_),
    .X(_3434_));
 sky130_fd_sc_hd__xor2_4 _7133_ (.A(\ks1.col[6] ),
    .B(_3434_),
    .X(_3435_));
 sky130_fd_sc_hd__mux2_1 _7134_ (.A0(\ks1.key_reg[70] ),
    .A1(net225),
    .S(_3419_),
    .X(_3436_));
 sky130_fd_sc_hd__xor2_2 _7135_ (.A(_3435_),
    .B(_3436_),
    .X(_3437_));
 sky130_fd_sc_hd__mux2_1 _7136_ (.A0(\ks1.key_reg[38] ),
    .A1(net189),
    .S(_3386_),
    .X(_3438_));
 sky130_fd_sc_hd__xor2_1 _7137_ (.A(_3437_),
    .B(_3438_),
    .X(_3439_));
 sky130_fd_sc_hd__or2_1 _7138_ (.A(_0812_),
    .B(_3439_),
    .X(_3440_));
 sky130_fd_sc_hd__a21oi_1 _7139_ (.A1(_0812_),
    .A2(_3439_),
    .B1(_3399_),
    .Y(_3441_));
 sky130_fd_sc_hd__a22o_1 _7140_ (.A1(net513),
    .A2(_3375_),
    .B1(_3440_),
    .B2(_3441_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _7141_ (.A0(\ks1.key_reg[103] ),
    .A1(net134),
    .S(_3377_),
    .X(_3442_));
 sky130_fd_sc_hd__xor2_2 _7142_ (.A(\ks1.col[7] ),
    .B(_3442_),
    .X(_3443_));
 sky130_fd_sc_hd__mux2_1 _7143_ (.A0(\ks1.key_reg[71] ),
    .A1(net226),
    .S(_3419_),
    .X(_3444_));
 sky130_fd_sc_hd__xor2_2 _7144_ (.A(_3443_),
    .B(_3444_),
    .X(_3445_));
 sky130_fd_sc_hd__mux2_1 _7145_ (.A0(\ks1.key_reg[39] ),
    .A1(net190),
    .S(_3386_),
    .X(_3446_));
 sky130_fd_sc_hd__xor2_2 _7146_ (.A(_3445_),
    .B(_3446_),
    .X(_3447_));
 sky130_fd_sc_hd__or2_1 _7147_ (.A(_1017_),
    .B(_3447_),
    .X(_3448_));
 sky130_fd_sc_hd__a21oi_1 _7148_ (.A1(_1017_),
    .A2(_3447_),
    .B1(_3399_),
    .Y(_3449_));
 sky130_fd_sc_hd__a22o_1 _7149_ (.A1(net509),
    .A2(_3375_),
    .B1(_3448_),
    .B2(_3449_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _7150_ (.A0(\ks1.key_reg[104] ),
    .A1(net135),
    .S(_0810_),
    .X(_3450_));
 sky130_fd_sc_hd__xnor2_2 _7151_ (.A(_1212_),
    .B(_3450_),
    .Y(_3451_));
 sky130_fd_sc_hd__buf_4 _7152_ (.A(_3376_),
    .X(_3452_));
 sky130_fd_sc_hd__mux2_1 _7153_ (.A0(\ks1.key_reg[72] ),
    .A1(net227),
    .S(_3452_),
    .X(_3453_));
 sky130_fd_sc_hd__xnor2_1 _7154_ (.A(_3451_),
    .B(_3453_),
    .Y(_3454_));
 sky130_fd_sc_hd__buf_4 _7155_ (.A(_3381_),
    .X(_3455_));
 sky130_fd_sc_hd__mux2_1 _7156_ (.A0(\ks1.key_reg[40] ),
    .A1(net192),
    .S(_3455_),
    .X(_3456_));
 sky130_fd_sc_hd__xnor2_1 _7157_ (.A(_3454_),
    .B(_3456_),
    .Y(_3457_));
 sky130_fd_sc_hd__xnor2_1 _7158_ (.A(_0935_),
    .B(_3457_),
    .Y(_3458_));
 sky130_fd_sc_hd__buf_4 _7159_ (.A(_1112_),
    .X(_3459_));
 sky130_fd_sc_hd__mux2_1 _7160_ (.A0(net650),
    .A1(_3458_),
    .S(_3459_),
    .X(_3460_));
 sky130_fd_sc_hd__clkbuf_1 _7161_ (.A(_3460_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _7162_ (.A0(\ks1.key_reg[105] ),
    .A1(net136),
    .S(_3376_),
    .X(_3461_));
 sky130_fd_sc_hd__xor2_2 _7163_ (.A(_1246_),
    .B(_3461_),
    .X(_3462_));
 sky130_fd_sc_hd__mux2_1 _7164_ (.A0(\ks1.key_reg[73] ),
    .A1(net228),
    .S(_3381_),
    .X(_3463_));
 sky130_fd_sc_hd__xor2_2 _7165_ (.A(_3462_),
    .B(_3463_),
    .X(_3464_));
 sky130_fd_sc_hd__mux2_1 _7166_ (.A0(\ks1.key_reg[41] ),
    .A1(net193),
    .S(_3382_),
    .X(_3465_));
 sky130_fd_sc_hd__xnor2_2 _7167_ (.A(_3464_),
    .B(_3465_),
    .Y(_3466_));
 sky130_fd_sc_hd__xnor2_1 _7168_ (.A(_0762_),
    .B(_3466_),
    .Y(_3467_));
 sky130_fd_sc_hd__mux2_1 _7169_ (.A0(net674),
    .A1(_3467_),
    .S(_3459_),
    .X(_3468_));
 sky130_fd_sc_hd__clkbuf_1 _7170_ (.A(_3468_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _7171_ (.A0(\ks1.key_reg[42] ),
    .A1(net194),
    .S(_3385_),
    .X(_3469_));
 sky130_fd_sc_hd__mux2_1 _7172_ (.A0(\ks1.key_reg[74] ),
    .A1(net229),
    .S(_3382_),
    .X(_3470_));
 sky130_fd_sc_hd__mux2_1 _7173_ (.A0(\ks1.key_reg[106] ),
    .A1(net137),
    .S(_3452_),
    .X(_3471_));
 sky130_fd_sc_hd__xor2_2 _7174_ (.A(_1256_),
    .B(_3471_),
    .X(_3472_));
 sky130_fd_sc_hd__xor2_1 _7175_ (.A(_3470_),
    .B(_3472_),
    .X(_3473_));
 sky130_fd_sc_hd__xor2_1 _7176_ (.A(_3469_),
    .B(_3473_),
    .X(_3474_));
 sky130_fd_sc_hd__or2_1 _7177_ (.A(_1058_),
    .B(_3474_),
    .X(_3475_));
 sky130_fd_sc_hd__a21oi_1 _7178_ (.A1(_1058_),
    .A2(_3474_),
    .B1(_3399_),
    .Y(_3476_));
 sky130_fd_sc_hd__a22o_1 _7179_ (.A1(net495),
    .A2(_3375_),
    .B1(_3475_),
    .B2(_3476_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _7180_ (.A0(\ks1.key_reg[43] ),
    .A1(net195),
    .S(_3385_),
    .X(_3477_));
 sky130_fd_sc_hd__mux2_1 _7181_ (.A0(\ks1.key_reg[75] ),
    .A1(net230),
    .S(_3382_),
    .X(_3478_));
 sky130_fd_sc_hd__mux2_1 _7182_ (.A0(\ks1.key_reg[107] ),
    .A1(net138),
    .S(_3377_),
    .X(_3479_));
 sky130_fd_sc_hd__xnor2_2 _7183_ (.A(_1271_),
    .B(_3479_),
    .Y(_3480_));
 sky130_fd_sc_hd__xnor2_2 _7184_ (.A(_3478_),
    .B(_3480_),
    .Y(_3481_));
 sky130_fd_sc_hd__xor2_2 _7185_ (.A(_3477_),
    .B(_3481_),
    .X(_3482_));
 sky130_fd_sc_hd__or2_1 _7186_ (.A(_0851_),
    .B(_3482_),
    .X(_3483_));
 sky130_fd_sc_hd__a21oi_1 _7187_ (.A1(_0851_),
    .A2(_3482_),
    .B1(_3399_),
    .Y(_3484_));
 sky130_fd_sc_hd__a22o_1 _7188_ (.A1(net506),
    .A2(_3375_),
    .B1(_3483_),
    .B2(_3484_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _7189_ (.A0(\ks1.key_reg[108] ),
    .A1(net139),
    .S(_0810_),
    .X(_3485_));
 sky130_fd_sc_hd__xnor2_1 _7190_ (.A(_1277_),
    .B(_3485_),
    .Y(_3486_));
 sky130_fd_sc_hd__mux2_1 _7191_ (.A0(\ks1.key_reg[76] ),
    .A1(net231),
    .S(_3452_),
    .X(_3487_));
 sky130_fd_sc_hd__xnor2_1 _7192_ (.A(_3486_),
    .B(_3487_),
    .Y(_3488_));
 sky130_fd_sc_hd__mux2_1 _7193_ (.A0(\ks1.key_reg[44] ),
    .A1(net196),
    .S(_3382_),
    .X(_3489_));
 sky130_fd_sc_hd__xnor2_1 _7194_ (.A(_3488_),
    .B(_3489_),
    .Y(_3490_));
 sky130_fd_sc_hd__xnor2_1 _7195_ (.A(_0892_),
    .B(_3490_),
    .Y(_3491_));
 sky130_fd_sc_hd__mux2_1 _7196_ (.A0(net625),
    .A1(_3491_),
    .S(_3459_),
    .X(_3492_));
 sky130_fd_sc_hd__clkbuf_1 _7197_ (.A(_3492_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _7198_ (.A0(\ks1.key_reg[45] ),
    .A1(net197),
    .S(_3455_),
    .X(_3493_));
 sky130_fd_sc_hd__mux2_2 _7199_ (.A0(\ks1.key_reg[77] ),
    .A1(net232),
    .S(_3381_),
    .X(_3494_));
 sky130_fd_sc_hd__mux2_2 _7200_ (.A0(\ks1.key_reg[109] ),
    .A1(net140),
    .S(_3380_),
    .X(_3495_));
 sky130_fd_sc_hd__xor2_4 _7201_ (.A(_1285_),
    .B(_3495_),
    .X(_3496_));
 sky130_fd_sc_hd__xnor2_4 _7202_ (.A(_3494_),
    .B(_3496_),
    .Y(_3497_));
 sky130_fd_sc_hd__xor2_2 _7203_ (.A(_3493_),
    .B(_3497_),
    .X(_3498_));
 sky130_fd_sc_hd__nor2_1 _7204_ (.A(_0976_),
    .B(_3498_),
    .Y(_3499_));
 sky130_fd_sc_hd__a21o_1 _7205_ (.A1(_0976_),
    .A2(_3498_),
    .B1(_3374_),
    .X(_3500_));
 sky130_fd_sc_hd__o22a_1 _7206_ (.A1(net500),
    .A2(\ks1.next_ready_o ),
    .B1(_3499_),
    .B2(_3500_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_2 _7207_ (.A0(\ks1.key_reg[110] ),
    .A1(net142),
    .S(_0810_),
    .X(_3501_));
 sky130_fd_sc_hd__xnor2_4 _7208_ (.A(_1292_),
    .B(_3501_),
    .Y(_3502_));
 sky130_fd_sc_hd__mux2_2 _7209_ (.A0(\ks1.key_reg[78] ),
    .A1(net233),
    .S(_3452_),
    .X(_3503_));
 sky130_fd_sc_hd__xor2_4 _7210_ (.A(_3502_),
    .B(_3503_),
    .X(_3504_));
 sky130_fd_sc_hd__mux2_2 _7211_ (.A0(\ks1.key_reg[46] ),
    .A1(net198),
    .S(_3455_),
    .X(_3505_));
 sky130_fd_sc_hd__xor2_4 _7212_ (.A(_3504_),
    .B(_3505_),
    .X(_3506_));
 sky130_fd_sc_hd__xnor2_1 _7213_ (.A(_0813_),
    .B(_3506_),
    .Y(_3507_));
 sky130_fd_sc_hd__mux2_1 _7214_ (.A0(net649),
    .A1(_3507_),
    .S(_3459_),
    .X(_3508_));
 sky130_fd_sc_hd__clkbuf_1 _7215_ (.A(_3508_),
    .X(_0491_));
 sky130_fd_sc_hd__clkbuf_4 _7216_ (.A(_3374_),
    .X(_3509_));
 sky130_fd_sc_hd__mux2_1 _7217_ (.A0(\ks1.key_reg[47] ),
    .A1(net199),
    .S(_3386_),
    .X(_3510_));
 sky130_fd_sc_hd__mux2_1 _7218_ (.A0(\ks1.key_reg[111] ),
    .A1(net143),
    .S(_3377_),
    .X(_3511_));
 sky130_fd_sc_hd__xor2_2 _7219_ (.A(_1299_),
    .B(_3511_),
    .X(_3512_));
 sky130_fd_sc_hd__mux2_1 _7220_ (.A0(\ks1.key_reg[79] ),
    .A1(net234),
    .S(_3382_),
    .X(_3513_));
 sky130_fd_sc_hd__xnor2_2 _7221_ (.A(_3512_),
    .B(_3513_),
    .Y(_3514_));
 sky130_fd_sc_hd__xnor2_1 _7222_ (.A(_3510_),
    .B(_3514_),
    .Y(_3515_));
 sky130_fd_sc_hd__nand2_1 _7223_ (.A(_1019_),
    .B(_3515_),
    .Y(_3516_));
 sky130_fd_sc_hd__o21a_1 _7224_ (.A1(_1019_),
    .A2(_3515_),
    .B1(_1113_),
    .X(_3517_));
 sky130_fd_sc_hd__a22o_1 _7225_ (.A1(net510),
    .A2(_3509_),
    .B1(_3516_),
    .B2(_3517_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_2 _7226_ (.A0(\ks1.key_reg[112] ),
    .A1(net144),
    .S(_3380_),
    .X(_3518_));
 sky130_fd_sc_hd__xor2_4 _7227_ (.A(\ks1.col[16] ),
    .B(_3518_),
    .X(_3519_));
 sky130_fd_sc_hd__mux2_1 _7228_ (.A0(\ks1.key_reg[80] ),
    .A1(net236),
    .S(_3419_),
    .X(_3520_));
 sky130_fd_sc_hd__xor2_1 _7229_ (.A(_3519_),
    .B(_3520_),
    .X(_3521_));
 sky130_fd_sc_hd__mux2_1 _7230_ (.A0(\ks1.key_reg[48] ),
    .A1(net200),
    .S(_3386_),
    .X(_3522_));
 sky130_fd_sc_hd__xor2_1 _7231_ (.A(_3521_),
    .B(_3522_),
    .X(_3523_));
 sky130_fd_sc_hd__or2_1 _7232_ (.A(_0933_),
    .B(_3523_),
    .X(_3524_));
 sky130_fd_sc_hd__a21oi_1 _7233_ (.A1(_0933_),
    .A2(_3523_),
    .B1(_3399_),
    .Y(_3525_));
 sky130_fd_sc_hd__a22o_1 _7234_ (.A1(net515),
    .A2(_3509_),
    .B1(_3524_),
    .B2(_3525_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _7235_ (.A0(\ks1.key_reg[113] ),
    .A1(net145),
    .S(_3380_),
    .X(_3526_));
 sky130_fd_sc_hd__xor2_2 _7236_ (.A(\ks1.col[17] ),
    .B(_3526_),
    .X(_3527_));
 sky130_fd_sc_hd__mux2_1 _7237_ (.A0(\ks1.key_reg[81] ),
    .A1(net237),
    .S(_3419_),
    .X(_3528_));
 sky130_fd_sc_hd__xor2_2 _7238_ (.A(_3527_),
    .B(_3528_),
    .X(_3529_));
 sky130_fd_sc_hd__mux2_1 _7239_ (.A0(\ks1.key_reg[49] ),
    .A1(net201),
    .S(_3385_),
    .X(_3530_));
 sky130_fd_sc_hd__xor2_2 _7240_ (.A(_3529_),
    .B(_3530_),
    .X(_3531_));
 sky130_fd_sc_hd__or2_1 _7241_ (.A(_0764_),
    .B(_3531_),
    .X(_3532_));
 sky130_fd_sc_hd__a21oi_1 _7242_ (.A1(_0764_),
    .A2(_3531_),
    .B1(_3374_),
    .Y(_3533_));
 sky130_fd_sc_hd__a22o_1 _7243_ (.A1(net517),
    .A2(_3509_),
    .B1(_3532_),
    .B2(_3533_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _7244_ (.A0(\ks1.key_reg[114] ),
    .A1(net146),
    .S(_3380_),
    .X(_3534_));
 sky130_fd_sc_hd__xor2_2 _7245_ (.A(\ks1.col[18] ),
    .B(_3534_),
    .X(_3535_));
 sky130_fd_sc_hd__mux2_1 _7246_ (.A0(\ks1.key_reg[82] ),
    .A1(net238),
    .S(_3419_),
    .X(_3536_));
 sky130_fd_sc_hd__xor2_2 _7247_ (.A(_3535_),
    .B(_3536_),
    .X(_3537_));
 sky130_fd_sc_hd__mux2_1 _7248_ (.A0(\ks1.key_reg[50] ),
    .A1(net203),
    .S(_3385_),
    .X(_3538_));
 sky130_fd_sc_hd__xor2_1 _7249_ (.A(_3537_),
    .B(_3538_),
    .X(_3539_));
 sky130_fd_sc_hd__or2_1 _7250_ (.A(_1059_),
    .B(_3539_),
    .X(_3540_));
 sky130_fd_sc_hd__a21oi_1 _7251_ (.A1(_1059_),
    .A2(_3539_),
    .B1(_3374_),
    .Y(_3541_));
 sky130_fd_sc_hd__a22o_1 _7252_ (.A1(net523),
    .A2(_3509_),
    .B1(_3540_),
    .B2(_3541_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _7253_ (.A0(\ks1.key_reg[115] ),
    .A1(net147),
    .S(_3380_),
    .X(_3542_));
 sky130_fd_sc_hd__xor2_1 _7254_ (.A(\ks1.col[19] ),
    .B(_3542_),
    .X(_3543_));
 sky130_fd_sc_hd__mux2_1 _7255_ (.A0(\ks1.key_reg[83] ),
    .A1(net239),
    .S(_3419_),
    .X(_3544_));
 sky130_fd_sc_hd__xor2_1 _7256_ (.A(_3543_),
    .B(_3544_),
    .X(_3545_));
 sky130_fd_sc_hd__mux2_1 _7257_ (.A0(\ks1.key_reg[51] ),
    .A1(net204),
    .S(_3385_),
    .X(_3546_));
 sky130_fd_sc_hd__xor2_1 _7258_ (.A(_3545_),
    .B(_3546_),
    .X(_3547_));
 sky130_fd_sc_hd__or2_1 _7259_ (.A(_0852_),
    .B(_3547_),
    .X(_3548_));
 sky130_fd_sc_hd__a21oi_1 _7260_ (.A1(_0852_),
    .A2(_3547_),
    .B1(_3374_),
    .Y(_3549_));
 sky130_fd_sc_hd__a22o_1 _7261_ (.A1(net499),
    .A2(_3509_),
    .B1(_3548_),
    .B2(_3549_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_2 _7262_ (.A0(\ks1.key_reg[116] ),
    .A1(net148),
    .S(_3380_),
    .X(_3550_));
 sky130_fd_sc_hd__xor2_4 _7263_ (.A(\ks1.col[20] ),
    .B(_3550_),
    .X(_3551_));
 sky130_fd_sc_hd__mux2_2 _7264_ (.A0(\ks1.key_reg[84] ),
    .A1(net240),
    .S(_3419_),
    .X(_3552_));
 sky130_fd_sc_hd__xor2_4 _7265_ (.A(_3551_),
    .B(_3552_),
    .X(_3553_));
 sky130_fd_sc_hd__mux2_1 _7266_ (.A0(\ks1.key_reg[52] ),
    .A1(net205),
    .S(_3385_),
    .X(_3554_));
 sky130_fd_sc_hd__xor2_1 _7267_ (.A(_3553_),
    .B(_3554_),
    .X(_3555_));
 sky130_fd_sc_hd__or2_1 _7268_ (.A(_0891_),
    .B(_3555_),
    .X(_3556_));
 sky130_fd_sc_hd__a21oi_1 _7269_ (.A1(_0891_),
    .A2(_3555_),
    .B1(_3374_),
    .Y(_3557_));
 sky130_fd_sc_hd__a22o_1 _7270_ (.A1(net496),
    .A2(_3509_),
    .B1(_3556_),
    .B2(_3557_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _7271_ (.A0(\ks1.key_reg[117] ),
    .A1(net149),
    .S(_3380_),
    .X(_3558_));
 sky130_fd_sc_hd__xor2_1 _7272_ (.A(\ks1.col[21] ),
    .B(_3558_),
    .X(_3559_));
 sky130_fd_sc_hd__mux2_1 _7273_ (.A0(\ks1.key_reg[85] ),
    .A1(net241),
    .S(_3419_),
    .X(_3560_));
 sky130_fd_sc_hd__xor2_1 _7274_ (.A(_3559_),
    .B(_3560_),
    .X(_3561_));
 sky130_fd_sc_hd__mux2_1 _7275_ (.A0(\ks1.key_reg[53] ),
    .A1(net206),
    .S(_3385_),
    .X(_3562_));
 sky130_fd_sc_hd__xor2_1 _7276_ (.A(_3561_),
    .B(_3562_),
    .X(_3563_));
 sky130_fd_sc_hd__or2_1 _7277_ (.A(_0975_),
    .B(_3563_),
    .X(_3564_));
 sky130_fd_sc_hd__a21oi_1 _7278_ (.A1(_0975_),
    .A2(_3563_),
    .B1(_3374_),
    .Y(_3565_));
 sky130_fd_sc_hd__a22o_1 _7279_ (.A1(net498),
    .A2(_3509_),
    .B1(_3564_),
    .B2(_3565_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _7280_ (.A0(\ks1.key_reg[118] ),
    .A1(net150),
    .S(_3380_),
    .X(_3566_));
 sky130_fd_sc_hd__xor2_2 _7281_ (.A(\ks1.col[22] ),
    .B(_3566_),
    .X(_3567_));
 sky130_fd_sc_hd__mux2_1 _7282_ (.A0(\ks1.key_reg[86] ),
    .A1(net242),
    .S(_3381_),
    .X(_3568_));
 sky130_fd_sc_hd__xor2_2 _7283_ (.A(_3567_),
    .B(_3568_),
    .X(_3569_));
 sky130_fd_sc_hd__mux2_1 _7284_ (.A0(\ks1.key_reg[54] ),
    .A1(net207),
    .S(_3385_),
    .X(_3570_));
 sky130_fd_sc_hd__xor2_2 _7285_ (.A(_3569_),
    .B(_3570_),
    .X(_3571_));
 sky130_fd_sc_hd__or2_1 _7286_ (.A(_0811_),
    .B(_3571_),
    .X(_3572_));
 sky130_fd_sc_hd__a21oi_1 _7287_ (.A1(_0811_),
    .A2(_3571_),
    .B1(_3374_),
    .Y(_3573_));
 sky130_fd_sc_hd__a22o_1 _7288_ (.A1(net504),
    .A2(_3509_),
    .B1(_3572_),
    .B2(_3573_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _7289_ (.A0(\ks1.key_reg[119] ),
    .A1(net151),
    .S(_3380_),
    .X(_3574_));
 sky130_fd_sc_hd__xor2_2 _7290_ (.A(\ks1.col[23] ),
    .B(_3574_),
    .X(_3575_));
 sky130_fd_sc_hd__mux2_1 _7291_ (.A0(\ks1.key_reg[87] ),
    .A1(net243),
    .S(_3381_),
    .X(_3576_));
 sky130_fd_sc_hd__xor2_2 _7292_ (.A(_3575_),
    .B(_3576_),
    .X(_3577_));
 sky130_fd_sc_hd__mux2_1 _7293_ (.A0(\ks1.key_reg[55] ),
    .A1(net208),
    .S(_3385_),
    .X(_3578_));
 sky130_fd_sc_hd__xor2_2 _7294_ (.A(_3577_),
    .B(_3578_),
    .X(_3579_));
 sky130_fd_sc_hd__or2_1 _7295_ (.A(_1018_),
    .B(_3579_),
    .X(_3580_));
 sky130_fd_sc_hd__a21oi_1 _7296_ (.A1(_1018_),
    .A2(_3579_),
    .B1(_3374_),
    .Y(_3581_));
 sky130_fd_sc_hd__a22o_1 _7297_ (.A1(net503),
    .A2(_3509_),
    .B1(_3580_),
    .B2(_3581_),
    .X(_0500_));
 sky130_fd_sc_hd__nand2_1 _7298_ (.A(\ks1.ready_o ),
    .B(_0669_),
    .Y(_3582_));
 sky130_fd_sc_hd__nor2_1 _7299_ (.A(_0674_),
    .B(_3582_),
    .Y(_3583_));
 sky130_fd_sc_hd__o221ai_4 _7300_ (.A1(\addroundkey_round[1] ),
    .A2(_3583_),
    .B1(_1132_),
    .B2(_0750_),
    .C1(_0748_),
    .Y(_3584_));
 sky130_fd_sc_hd__a31oi_4 _7301_ (.A1(\addroundkey_round[2] ),
    .A2(_0748_),
    .A3(_0750_),
    .B1(_1135_),
    .Y(_3585_));
 sky130_fd_sc_hd__o21a_1 _7302_ (.A1(_0674_),
    .A2(_3582_),
    .B1(\addroundkey_round[0] ),
    .X(_3586_));
 sky130_fd_sc_hd__or3_2 _7303_ (.A(_0759_),
    .B(_1130_),
    .C(_3586_),
    .X(_3587_));
 sky130_fd_sc_hd__and3_1 _7304_ (.A(_3584_),
    .B(_3585_),
    .C(_3587_),
    .X(_3588_));
 sky130_fd_sc_hd__xnor2_2 _7305_ (.A(\ks1.col[24] ),
    .B(_3588_),
    .Y(_3589_));
 sky130_fd_sc_hd__mux2_1 _7306_ (.A0(\ks1.key_reg[120] ),
    .A1(net153),
    .S(_3376_),
    .X(_3590_));
 sky130_fd_sc_hd__xor2_2 _7307_ (.A(_3589_),
    .B(_3590_),
    .X(_3591_));
 sky130_fd_sc_hd__mux2_1 _7308_ (.A0(\ks1.key_reg[88] ),
    .A1(net244),
    .S(_3452_),
    .X(_3592_));
 sky130_fd_sc_hd__xnor2_2 _7309_ (.A(_3591_),
    .B(_3592_),
    .Y(_3593_));
 sky130_fd_sc_hd__mux2_1 _7310_ (.A0(\ks1.key_reg[56] ),
    .A1(net209),
    .S(_3455_),
    .X(_3594_));
 sky130_fd_sc_hd__xnor2_1 _7311_ (.A(_3593_),
    .B(_3594_),
    .Y(_3595_));
 sky130_fd_sc_hd__xnor2_1 _7312_ (.A(_0937_),
    .B(_3595_),
    .Y(_3596_));
 sky130_fd_sc_hd__mux2_1 _7313_ (.A0(\ks1.key_reg[24] ),
    .A1(_3596_),
    .S(_3459_),
    .X(_3597_));
 sky130_fd_sc_hd__clkbuf_1 _7314_ (.A(_3597_),
    .X(_0501_));
 sky130_fd_sc_hd__xnor2_1 _7315_ (.A(_3584_),
    .B(_3587_),
    .Y(_3598_));
 sky130_fd_sc_hd__a31oi_2 _7316_ (.A1(\addroundkey_round[3] ),
    .A2(_0748_),
    .A3(_0750_),
    .B1(_1137_),
    .Y(_3599_));
 sky130_fd_sc_hd__nand2_1 _7317_ (.A(_3587_),
    .B(_3599_),
    .Y(_3600_));
 sky130_fd_sc_hd__and3_1 _7318_ (.A(_3585_),
    .B(_3598_),
    .C(_3600_),
    .X(_3601_));
 sky130_fd_sc_hd__xor2_2 _7319_ (.A(\ks1.col[25] ),
    .B(_3601_),
    .X(_3602_));
 sky130_fd_sc_hd__mux2_1 _7320_ (.A0(\ks1.key_reg[121] ),
    .A1(net154),
    .S(_3376_),
    .X(_3603_));
 sky130_fd_sc_hd__xnor2_2 _7321_ (.A(_3602_),
    .B(_3603_),
    .Y(_3604_));
 sky130_fd_sc_hd__mux2_1 _7322_ (.A0(\ks1.key_reg[89] ),
    .A1(net245),
    .S(_3381_),
    .X(_3605_));
 sky130_fd_sc_hd__xor2_2 _7323_ (.A(_3604_),
    .B(_3605_),
    .X(_3606_));
 sky130_fd_sc_hd__mux2_1 _7324_ (.A0(\ks1.key_reg[57] ),
    .A1(net210),
    .S(_3455_),
    .X(_3607_));
 sky130_fd_sc_hd__xor2_1 _7325_ (.A(_3606_),
    .B(_3607_),
    .X(_3608_));
 sky130_fd_sc_hd__xnor2_1 _7326_ (.A(_0770_),
    .B(_3608_),
    .Y(_3609_));
 sky130_fd_sc_hd__mux2_1 _7327_ (.A0(net612),
    .A1(_3609_),
    .S(_3459_),
    .X(_3610_));
 sky130_fd_sc_hd__clkbuf_1 _7328_ (.A(_3610_),
    .X(_0502_));
 sky130_fd_sc_hd__inv_2 _7329_ (.A(_3585_),
    .Y(_3611_));
 sky130_fd_sc_hd__or2_1 _7330_ (.A(_3587_),
    .B(_3599_),
    .X(_3612_));
 sky130_fd_sc_hd__and2_1 _7331_ (.A(_3600_),
    .B(_3612_),
    .X(_3613_));
 sky130_fd_sc_hd__or3_2 _7332_ (.A(_3584_),
    .B(_3611_),
    .C(_3613_),
    .X(_3614_));
 sky130_fd_sc_hd__xnor2_2 _7333_ (.A(\ks1.col[26] ),
    .B(_3614_),
    .Y(_3615_));
 sky130_fd_sc_hd__mux2_1 _7334_ (.A0(\ks1.key_reg[122] ),
    .A1(net155),
    .S(_3376_),
    .X(_3616_));
 sky130_fd_sc_hd__xnor2_2 _7335_ (.A(_3615_),
    .B(_3616_),
    .Y(_3617_));
 sky130_fd_sc_hd__mux2_1 _7336_ (.A0(\ks1.key_reg[90] ),
    .A1(net247),
    .S(_3381_),
    .X(_3618_));
 sky130_fd_sc_hd__xor2_2 _7337_ (.A(_3617_),
    .B(_3618_),
    .X(_3619_));
 sky130_fd_sc_hd__mux2_1 _7338_ (.A0(\ks1.key_reg[58] ),
    .A1(net211),
    .S(_3455_),
    .X(_3620_));
 sky130_fd_sc_hd__xor2_2 _7339_ (.A(_3619_),
    .B(_3620_),
    .X(_3621_));
 sky130_fd_sc_hd__xnor2_1 _7340_ (.A(_1061_),
    .B(_3621_),
    .Y(_3622_));
 sky130_fd_sc_hd__mux2_1 _7341_ (.A0(net661),
    .A1(_3622_),
    .S(_3459_),
    .X(_3623_));
 sky130_fd_sc_hd__clkbuf_1 _7342_ (.A(_3623_),
    .X(_0503_));
 sky130_fd_sc_hd__xor2_1 _7343_ (.A(_3585_),
    .B(_3599_),
    .X(_3624_));
 sky130_fd_sc_hd__and3_2 _7344_ (.A(_3584_),
    .B(_3613_),
    .C(_3624_),
    .X(_3625_));
 sky130_fd_sc_hd__xnor2_4 _7345_ (.A(\ks1.col[27] ),
    .B(_3625_),
    .Y(_3626_));
 sky130_fd_sc_hd__mux2_2 _7346_ (.A0(\ks1.key_reg[123] ),
    .A1(net156),
    .S(_0810_),
    .X(_3627_));
 sky130_fd_sc_hd__xor2_4 _7347_ (.A(_3626_),
    .B(_3627_),
    .X(_3628_));
 sky130_fd_sc_hd__mux2_2 _7348_ (.A0(\ks1.key_reg[91] ),
    .A1(net248),
    .S(_3452_),
    .X(_3629_));
 sky130_fd_sc_hd__xnor2_4 _7349_ (.A(_3628_),
    .B(_3629_),
    .Y(_3630_));
 sky130_fd_sc_hd__mux2_1 _7350_ (.A0(\ks1.key_reg[59] ),
    .A1(net212),
    .S(_3382_),
    .X(_3631_));
 sky130_fd_sc_hd__xnor2_2 _7351_ (.A(_3630_),
    .B(_3631_),
    .Y(_3632_));
 sky130_fd_sc_hd__xnor2_1 _7352_ (.A(_0854_),
    .B(_3632_),
    .Y(_3633_));
 sky130_fd_sc_hd__mux2_1 _7353_ (.A0(net624),
    .A1(_3633_),
    .S(_3459_),
    .X(_3634_));
 sky130_fd_sc_hd__clkbuf_1 _7354_ (.A(_3634_),
    .X(_0504_));
 sky130_fd_sc_hd__o211a_1 _7355_ (.A1(_3585_),
    .A2(_3587_),
    .B1(_3598_),
    .C1(_3624_),
    .X(_3635_));
 sky130_fd_sc_hd__xor2_4 _7356_ (.A(\ks1.col[28] ),
    .B(_3635_),
    .X(_3636_));
 sky130_fd_sc_hd__mux2_2 _7357_ (.A0(\ks1.key_reg[124] ),
    .A1(net157),
    .S(_3376_),
    .X(_3637_));
 sky130_fd_sc_hd__xnor2_4 _7358_ (.A(_3636_),
    .B(_3637_),
    .Y(_3638_));
 sky130_fd_sc_hd__mux2_2 _7359_ (.A0(\ks1.key_reg[92] ),
    .A1(net249),
    .S(_3452_),
    .X(_3639_));
 sky130_fd_sc_hd__xor2_4 _7360_ (.A(_3638_),
    .B(_3639_),
    .X(_3640_));
 sky130_fd_sc_hd__mux2_1 _7361_ (.A0(\ks1.key_reg[60] ),
    .A1(net214),
    .S(_3455_),
    .X(_3641_));
 sky130_fd_sc_hd__xor2_2 _7362_ (.A(_3640_),
    .B(_3641_),
    .X(_3642_));
 sky130_fd_sc_hd__xnor2_1 _7363_ (.A(_0894_),
    .B(_3642_),
    .Y(_3643_));
 sky130_fd_sc_hd__mux2_1 _7364_ (.A0(net699),
    .A1(_3643_),
    .S(_3459_),
    .X(_3644_));
 sky130_fd_sc_hd__clkbuf_1 _7365_ (.A(_3644_),
    .X(_0505_));
 sky130_fd_sc_hd__or3b_1 _7366_ (.A(_3584_),
    .B(_3587_),
    .C_N(_3624_),
    .X(_3645_));
 sky130_fd_sc_hd__xnor2_2 _7367_ (.A(\ks1.col[29] ),
    .B(_3645_),
    .Y(_3646_));
 sky130_fd_sc_hd__mux2_2 _7368_ (.A0(\ks1.key_reg[125] ),
    .A1(net158),
    .S(_3376_),
    .X(_3647_));
 sky130_fd_sc_hd__xnor2_4 _7369_ (.A(_3646_),
    .B(_3647_),
    .Y(_3648_));
 sky130_fd_sc_hd__mux2_2 _7370_ (.A0(\ks1.key_reg[93] ),
    .A1(net250),
    .S(_3452_),
    .X(_3649_));
 sky130_fd_sc_hd__xor2_4 _7371_ (.A(_3648_),
    .B(_3649_),
    .X(_3650_));
 sky130_fd_sc_hd__mux2_1 _7372_ (.A0(\ks1.key_reg[61] ),
    .A1(net215),
    .S(_3455_),
    .X(_3651_));
 sky130_fd_sc_hd__xor2_2 _7373_ (.A(_3650_),
    .B(_3651_),
    .X(_3652_));
 sky130_fd_sc_hd__xnor2_1 _7374_ (.A(_0979_),
    .B(_3652_),
    .Y(_3653_));
 sky130_fd_sc_hd__mux2_1 _7375_ (.A0(net675),
    .A1(_3653_),
    .S(_3459_),
    .X(_3654_));
 sky130_fd_sc_hd__clkbuf_1 _7376_ (.A(_3654_),
    .X(_0506_));
 sky130_fd_sc_hd__or3_1 _7377_ (.A(_3584_),
    .B(_3585_),
    .C(_3600_),
    .X(_3655_));
 sky130_fd_sc_hd__xnor2_2 _7378_ (.A(\ks1.col[30] ),
    .B(_3655_),
    .Y(_3656_));
 sky130_fd_sc_hd__mux2_1 _7379_ (.A0(\ks1.key_reg[126] ),
    .A1(net159),
    .S(_3376_),
    .X(_3657_));
 sky130_fd_sc_hd__xnor2_2 _7380_ (.A(_3656_),
    .B(_3657_),
    .Y(_3658_));
 sky130_fd_sc_hd__mux2_1 _7381_ (.A0(\ks1.key_reg[94] ),
    .A1(net251),
    .S(_3452_),
    .X(_3659_));
 sky130_fd_sc_hd__xor2_2 _7382_ (.A(_3658_),
    .B(_3659_),
    .X(_3660_));
 sky130_fd_sc_hd__mux2_1 _7383_ (.A0(\ks1.key_reg[62] ),
    .A1(net216),
    .S(_3455_),
    .X(_3661_));
 sky130_fd_sc_hd__xor2_2 _7384_ (.A(_3660_),
    .B(_3661_),
    .X(_3662_));
 sky130_fd_sc_hd__xnor2_1 _7385_ (.A(_0816_),
    .B(_3662_),
    .Y(_3663_));
 sky130_fd_sc_hd__buf_4 _7386_ (.A(_1112_),
    .X(_3664_));
 sky130_fd_sc_hd__mux2_1 _7387_ (.A0(net643),
    .A1(_3663_),
    .S(_3664_),
    .X(_3665_));
 sky130_fd_sc_hd__clkbuf_1 _7388_ (.A(_3665_),
    .X(_0507_));
 sky130_fd_sc_hd__or4b_2 _7389_ (.A(_3611_),
    .B(_3587_),
    .C(_3599_),
    .D_N(_3584_),
    .X(_3666_));
 sky130_fd_sc_hd__xnor2_4 _7390_ (.A(\ks1.col[31] ),
    .B(_3666_),
    .Y(_3667_));
 sky130_fd_sc_hd__mux2_2 _7391_ (.A0(\ks1.key_reg[127] ),
    .A1(net160),
    .S(_3376_),
    .X(_3668_));
 sky130_fd_sc_hd__xnor2_4 _7392_ (.A(_3667_),
    .B(_3668_),
    .Y(_3669_));
 sky130_fd_sc_hd__mux2_2 _7393_ (.A0(\ks1.key_reg[95] ),
    .A1(net252),
    .S(_3452_),
    .X(_3670_));
 sky130_fd_sc_hd__xor2_4 _7394_ (.A(_3669_),
    .B(_3670_),
    .X(_3671_));
 sky130_fd_sc_hd__mux2_1 _7395_ (.A0(\ks1.key_reg[63] ),
    .A1(net217),
    .S(_3455_),
    .X(_3672_));
 sky130_fd_sc_hd__xor2_2 _7396_ (.A(_3671_),
    .B(_3672_),
    .X(_3673_));
 sky130_fd_sc_hd__xnor2_1 _7397_ (.A(_1021_),
    .B(_3673_),
    .Y(_3674_));
 sky130_fd_sc_hd__mux2_1 _7398_ (.A0(net693),
    .A1(_3674_),
    .S(_3664_),
    .X(_3675_));
 sky130_fd_sc_hd__clkbuf_1 _7399_ (.A(_3675_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _7400_ (.A0(net654),
    .A1(_3388_),
    .S(_3664_),
    .X(_3676_));
 sky130_fd_sc_hd__clkbuf_1 _7401_ (.A(_3676_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _7402_ (.A0(net657),
    .A1(_3397_),
    .S(_3664_),
    .X(_3677_));
 sky130_fd_sc_hd__clkbuf_1 _7403_ (.A(_3677_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _7404_ (.A0(net663),
    .A1(_3406_),
    .S(_3664_),
    .X(_3678_));
 sky130_fd_sc_hd__clkbuf_1 _7405_ (.A(_3678_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _7406_ (.A0(net702),
    .A1(_3414_),
    .S(_3664_),
    .X(_3679_));
 sky130_fd_sc_hd__clkbuf_1 _7407_ (.A(_3679_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _7408_ (.A0(net677),
    .A1(_3423_),
    .S(_3664_),
    .X(_3680_));
 sky130_fd_sc_hd__clkbuf_1 _7409_ (.A(_3680_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _7410_ (.A0(net698),
    .A1(_3431_),
    .S(_3664_),
    .X(_3681_));
 sky130_fd_sc_hd__clkbuf_1 _7411_ (.A(_3681_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _7412_ (.A0(net639),
    .A1(_3439_),
    .S(_3664_),
    .X(_3682_));
 sky130_fd_sc_hd__clkbuf_1 _7413_ (.A(_3682_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _7414_ (.A0(net648),
    .A1(_3447_),
    .S(_3664_),
    .X(_3683_));
 sky130_fd_sc_hd__clkbuf_1 _7415_ (.A(_3683_),
    .X(_0516_));
 sky130_fd_sc_hd__buf_4 _7416_ (.A(_0754_),
    .X(_3684_));
 sky130_fd_sc_hd__nand2_1 _7417_ (.A(net489),
    .B(_3684_),
    .Y(_3685_));
 sky130_fd_sc_hd__o21ai_1 _7418_ (.A1(_3509_),
    .A2(_3457_),
    .B1(_3685_),
    .Y(_0517_));
 sky130_fd_sc_hd__nor2_1 _7419_ (.A(net505),
    .B(_1113_),
    .Y(_3686_));
 sky130_fd_sc_hd__a21oi_1 _7420_ (.A1(\ks1.next_ready_o ),
    .A2(_3466_),
    .B1(_3686_),
    .Y(_0518_));
 sky130_fd_sc_hd__buf_4 _7421_ (.A(_1112_),
    .X(_3687_));
 sky130_fd_sc_hd__mux2_1 _7422_ (.A0(net692),
    .A1(_3474_),
    .S(_3687_),
    .X(_3688_));
 sky130_fd_sc_hd__clkbuf_1 _7423_ (.A(_3688_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _7424_ (.A0(net636),
    .A1(_3482_),
    .S(_3687_),
    .X(_3689_));
 sky130_fd_sc_hd__clkbuf_1 _7425_ (.A(_3689_),
    .X(_0520_));
 sky130_fd_sc_hd__nor2_1 _7426_ (.A(net494),
    .B(_1113_),
    .Y(_3690_));
 sky130_fd_sc_hd__a21oi_1 _7427_ (.A1(\ks1.next_ready_o ),
    .A2(_3490_),
    .B1(_3690_),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _7428_ (.A(_3498_),
    .Y(_3691_));
 sky130_fd_sc_hd__mux2_1 _7429_ (.A0(net666),
    .A1(_3691_),
    .S(_3687_),
    .X(_3692_));
 sky130_fd_sc_hd__clkbuf_1 _7430_ (.A(_3692_),
    .X(_0522_));
 sky130_fd_sc_hd__nor2_1 _7431_ (.A(net491),
    .B(_1113_),
    .Y(_3693_));
 sky130_fd_sc_hd__a21oi_1 _7432_ (.A1(\ks1.next_ready_o ),
    .A2(_3506_),
    .B1(_3693_),
    .Y(_0523_));
 sky130_fd_sc_hd__mux2_1 _7433_ (.A0(net645),
    .A1(_3515_),
    .S(_3687_),
    .X(_3694_));
 sky130_fd_sc_hd__clkbuf_1 _7434_ (.A(_3694_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _7435_ (.A0(net607),
    .A1(_3523_),
    .S(_3687_),
    .X(_3695_));
 sky130_fd_sc_hd__clkbuf_1 _7436_ (.A(_3695_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _7437_ (.A0(net647),
    .A1(_3531_),
    .S(_3687_),
    .X(_3696_));
 sky130_fd_sc_hd__clkbuf_1 _7438_ (.A(_3696_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _7439_ (.A0(net641),
    .A1(_3539_),
    .S(_3687_),
    .X(_3697_));
 sky130_fd_sc_hd__clkbuf_1 _7440_ (.A(_3697_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _7441_ (.A0(net617),
    .A1(_3547_),
    .S(_3687_),
    .X(_3698_));
 sky130_fd_sc_hd__clkbuf_1 _7442_ (.A(_3698_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _7443_ (.A0(net683),
    .A1(_3555_),
    .S(_3687_),
    .X(_3699_));
 sky130_fd_sc_hd__clkbuf_1 _7444_ (.A(_3699_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _7445_ (.A0(net638),
    .A1(_3563_),
    .S(_3687_),
    .X(_3700_));
 sky130_fd_sc_hd__clkbuf_1 _7446_ (.A(_3700_),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_8 _7447_ (.A(_1112_),
    .X(_3701_));
 sky130_fd_sc_hd__mux2_1 _7448_ (.A0(net653),
    .A1(_3571_),
    .S(_3701_),
    .X(_3702_));
 sky130_fd_sc_hd__clkbuf_1 _7449_ (.A(_3702_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _7450_ (.A0(net697),
    .A1(_3579_),
    .S(_3701_),
    .X(_3703_));
 sky130_fd_sc_hd__clkbuf_1 _7451_ (.A(_3703_),
    .X(_0532_));
 sky130_fd_sc_hd__nand2_1 _7452_ (.A(net514),
    .B(_3390_),
    .Y(_3704_));
 sky130_fd_sc_hd__o21ai_1 _7453_ (.A1(_3684_),
    .A2(_3595_),
    .B1(_3704_),
    .Y(_0533_));
 sky130_fd_sc_hd__nand2_1 _7454_ (.A(net490),
    .B(_3390_),
    .Y(_3705_));
 sky130_fd_sc_hd__o21ai_1 _7455_ (.A1(_3684_),
    .A2(_3608_),
    .B1(_3705_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _7456_ (.A(net484),
    .B(_3390_),
    .Y(_3706_));
 sky130_fd_sc_hd__o21ai_1 _7457_ (.A1(_3684_),
    .A2(_3621_),
    .B1(_3706_),
    .Y(_0535_));
 sky130_fd_sc_hd__nor2_1 _7458_ (.A(net501),
    .B(_1113_),
    .Y(_3707_));
 sky130_fd_sc_hd__a21oi_1 _7459_ (.A1(\ks1.next_ready_o ),
    .A2(_3632_),
    .B1(_3707_),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_1 _7460_ (.A(net486),
    .B(_3390_),
    .Y(_3708_));
 sky130_fd_sc_hd__o21ai_1 _7461_ (.A1(_3684_),
    .A2(_3642_),
    .B1(_3708_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _7462_ (.A(net487),
    .B(_3390_),
    .Y(_3709_));
 sky130_fd_sc_hd__o21ai_1 _7463_ (.A1(_3684_),
    .A2(_3652_),
    .B1(_3709_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_1 _7464_ (.A(net485),
    .B(_3390_),
    .Y(_3710_));
 sky130_fd_sc_hd__o21ai_1 _7465_ (.A1(_3684_),
    .A2(_3662_),
    .B1(_3710_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _7466_ (.A(net493),
    .B(_3390_),
    .Y(_3711_));
 sky130_fd_sc_hd__o21ai_1 _7467_ (.A1(_3684_),
    .A2(_3673_),
    .B1(_3711_),
    .Y(_0540_));
 sky130_fd_sc_hd__mux2_1 _7468_ (.A0(net628),
    .A1(_3384_),
    .S(_3701_),
    .X(_3712_));
 sky130_fd_sc_hd__clkbuf_1 _7469_ (.A(_3712_),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_1 _7470_ (.A0(net667),
    .A1(_3395_),
    .S(_3701_),
    .X(_3713_));
 sky130_fd_sc_hd__clkbuf_1 _7471_ (.A(_3713_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _7472_ (.A0(net632),
    .A1(_3404_),
    .S(_3701_),
    .X(_3714_));
 sky130_fd_sc_hd__clkbuf_1 _7473_ (.A(_3714_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _7474_ (.A0(net684),
    .A1(_3412_),
    .S(_3701_),
    .X(_3715_));
 sky130_fd_sc_hd__clkbuf_1 _7475_ (.A(_3715_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _7476_ (.A0(net634),
    .A1(_3421_),
    .S(_3701_),
    .X(_3716_));
 sky130_fd_sc_hd__clkbuf_1 _7477_ (.A(_3716_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _7478_ (.A0(net656),
    .A1(_3429_),
    .S(_3701_),
    .X(_3717_));
 sky130_fd_sc_hd__clkbuf_1 _7479_ (.A(_3717_),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _7480_ (.A0(net620),
    .A1(_3437_),
    .S(_3701_),
    .X(_3718_));
 sky130_fd_sc_hd__clkbuf_1 _7481_ (.A(_3718_),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _7482_ (.A0(net626),
    .A1(_3445_),
    .S(_3701_),
    .X(_3719_));
 sky130_fd_sc_hd__clkbuf_1 _7483_ (.A(_3719_),
    .X(_0548_));
 sky130_fd_sc_hd__buf_4 _7484_ (.A(_1112_),
    .X(_3720_));
 sky130_fd_sc_hd__mux2_1 _7485_ (.A0(net652),
    .A1(_3454_),
    .S(_3720_),
    .X(_3721_));
 sky130_fd_sc_hd__clkbuf_1 _7486_ (.A(_3721_),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _7487_ (.A0(net614),
    .A1(_3464_),
    .S(_3720_),
    .X(_3722_));
 sky130_fd_sc_hd__clkbuf_1 _7488_ (.A(_3722_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _7489_ (.A0(net688),
    .A1(_3473_),
    .S(_3720_),
    .X(_3723_));
 sky130_fd_sc_hd__clkbuf_1 _7490_ (.A(_3723_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _7491_ (.A0(net651),
    .A1(_3481_),
    .S(_3720_),
    .X(_3724_));
 sky130_fd_sc_hd__clkbuf_1 _7492_ (.A(_3724_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _7493_ (.A0(net655),
    .A1(_3488_),
    .S(_3720_),
    .X(_3725_));
 sky130_fd_sc_hd__clkbuf_1 _7494_ (.A(_3725_),
    .X(_0553_));
 sky130_fd_sc_hd__inv_2 _7495_ (.A(_3497_),
    .Y(_3726_));
 sky130_fd_sc_hd__mux2_1 _7496_ (.A0(\ks1.key_reg[77] ),
    .A1(_3726_),
    .S(_3720_),
    .X(_3727_));
 sky130_fd_sc_hd__clkbuf_1 _7497_ (.A(_3727_),
    .X(_0554_));
 sky130_fd_sc_hd__inv_2 _7498_ (.A(_3504_),
    .Y(_3728_));
 sky130_fd_sc_hd__mux2_1 _7499_ (.A0(net671),
    .A1(_3728_),
    .S(_3720_),
    .X(_3729_));
 sky130_fd_sc_hd__clkbuf_1 _7500_ (.A(_3729_),
    .X(_0555_));
 sky130_fd_sc_hd__nor2_1 _7501_ (.A(net492),
    .B(_1113_),
    .Y(_3730_));
 sky130_fd_sc_hd__a21oi_1 _7502_ (.A1(\ks1.next_ready_o ),
    .A2(_3514_),
    .B1(_3730_),
    .Y(_0556_));
 sky130_fd_sc_hd__mux2_1 _7503_ (.A0(net676),
    .A1(_3521_),
    .S(_3720_),
    .X(_3731_));
 sky130_fd_sc_hd__clkbuf_1 _7504_ (.A(_3731_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _7505_ (.A0(net635),
    .A1(_3529_),
    .S(_3720_),
    .X(_3732_));
 sky130_fd_sc_hd__clkbuf_1 _7506_ (.A(_3732_),
    .X(_0558_));
 sky130_fd_sc_hd__mux2_1 _7507_ (.A0(net705),
    .A1(_3537_),
    .S(_3720_),
    .X(_3733_));
 sky130_fd_sc_hd__clkbuf_1 _7508_ (.A(_3733_),
    .X(_0559_));
 sky130_fd_sc_hd__clkbuf_8 _7509_ (.A(_1112_),
    .X(_3734_));
 sky130_fd_sc_hd__mux2_1 _7510_ (.A0(net642),
    .A1(_3545_),
    .S(_3734_),
    .X(_3735_));
 sky130_fd_sc_hd__clkbuf_1 _7511_ (.A(_3735_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_1 _7512_ (.A0(net664),
    .A1(_3553_),
    .S(_3734_),
    .X(_3736_));
 sky130_fd_sc_hd__clkbuf_1 _7513_ (.A(_3736_),
    .X(_0561_));
 sky130_fd_sc_hd__mux2_1 _7514_ (.A0(net646),
    .A1(_3561_),
    .S(_3734_),
    .X(_3737_));
 sky130_fd_sc_hd__clkbuf_1 _7515_ (.A(_3737_),
    .X(_0562_));
 sky130_fd_sc_hd__mux2_1 _7516_ (.A0(net700),
    .A1(_3569_),
    .S(_3734_),
    .X(_3738_));
 sky130_fd_sc_hd__clkbuf_1 _7517_ (.A(_3738_),
    .X(_0563_));
 sky130_fd_sc_hd__mux2_1 _7518_ (.A0(net640),
    .A1(_3577_),
    .S(_3734_),
    .X(_3739_));
 sky130_fd_sc_hd__clkbuf_1 _7519_ (.A(_3739_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _7520_ (.A0(net631),
    .A1(_3593_),
    .S(_3734_),
    .X(_3740_));
 sky130_fd_sc_hd__clkbuf_1 _7521_ (.A(_3740_),
    .X(_0565_));
 sky130_fd_sc_hd__inv_2 _7522_ (.A(_3606_),
    .Y(_3741_));
 sky130_fd_sc_hd__mux2_1 _7523_ (.A0(net689),
    .A1(_3741_),
    .S(_3734_),
    .X(_3742_));
 sky130_fd_sc_hd__clkbuf_1 _7524_ (.A(_3742_),
    .X(_0566_));
 sky130_fd_sc_hd__inv_2 _7525_ (.A(_3619_),
    .Y(_3743_));
 sky130_fd_sc_hd__mux2_1 _7526_ (.A0(net665),
    .A1(_3743_),
    .S(_3734_),
    .X(_3744_));
 sky130_fd_sc_hd__clkbuf_1 _7527_ (.A(_3744_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_1 _7528_ (.A0(net621),
    .A1(_3630_),
    .S(_3734_),
    .X(_3745_));
 sky130_fd_sc_hd__clkbuf_1 _7529_ (.A(_3745_),
    .X(_0568_));
 sky130_fd_sc_hd__inv_2 _7530_ (.A(_3640_),
    .Y(_3746_));
 sky130_fd_sc_hd__mux2_1 _7531_ (.A0(net644),
    .A1(_3746_),
    .S(_3734_),
    .X(_3747_));
 sky130_fd_sc_hd__clkbuf_1 _7532_ (.A(_3747_),
    .X(_0569_));
 sky130_fd_sc_hd__inv_2 _7533_ (.A(_3650_),
    .Y(_3748_));
 sky130_fd_sc_hd__clkbuf_8 _7534_ (.A(_1112_),
    .X(_3749_));
 sky130_fd_sc_hd__mux2_1 _7535_ (.A0(net630),
    .A1(_3748_),
    .S(_3749_),
    .X(_3750_));
 sky130_fd_sc_hd__clkbuf_1 _7536_ (.A(_3750_),
    .X(_0570_));
 sky130_fd_sc_hd__inv_2 _7537_ (.A(_3660_),
    .Y(_3751_));
 sky130_fd_sc_hd__mux2_1 _7538_ (.A0(net662),
    .A1(_3751_),
    .S(_3749_),
    .X(_3752_));
 sky130_fd_sc_hd__clkbuf_1 _7539_ (.A(_3752_),
    .X(_0571_));
 sky130_fd_sc_hd__inv_2 _7540_ (.A(_3671_),
    .Y(_3753_));
 sky130_fd_sc_hd__mux2_1 _7541_ (.A0(net615),
    .A1(_3753_),
    .S(_3749_),
    .X(_3754_));
 sky130_fd_sc_hd__clkbuf_1 _7542_ (.A(_3754_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _7543_ (.A0(\ks1.key_reg[96] ),
    .A1(_3379_),
    .S(_3749_),
    .X(_3755_));
 sky130_fd_sc_hd__clkbuf_1 _7544_ (.A(_3755_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _7545_ (.A0(net678),
    .A1(_3393_),
    .S(_3749_),
    .X(_3756_));
 sky130_fd_sc_hd__clkbuf_1 _7546_ (.A(_3756_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _7547_ (.A0(net703),
    .A1(_3402_),
    .S(_3749_),
    .X(_3757_));
 sky130_fd_sc_hd__clkbuf_1 _7548_ (.A(_3757_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _7549_ (.A0(net672),
    .A1(_3410_),
    .S(_3749_),
    .X(_3758_));
 sky130_fd_sc_hd__clkbuf_1 _7550_ (.A(_3758_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _7551_ (.A0(net680),
    .A1(_3418_),
    .S(_3749_),
    .X(_3759_));
 sky130_fd_sc_hd__clkbuf_1 _7552_ (.A(_3759_),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _7553_ (.A0(net696),
    .A1(_3427_),
    .S(_3749_),
    .X(_3760_));
 sky130_fd_sc_hd__clkbuf_1 _7554_ (.A(_3760_),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _7555_ (.A0(net637),
    .A1(_3435_),
    .S(_3749_),
    .X(_3761_));
 sky130_fd_sc_hd__clkbuf_1 _7556_ (.A(_3761_),
    .X(_0579_));
 sky130_fd_sc_hd__clkbuf_8 _7557_ (.A(_1112_),
    .X(_3762_));
 sky130_fd_sc_hd__mux2_1 _7558_ (.A0(net669),
    .A1(_3443_),
    .S(_3762_),
    .X(_3763_));
 sky130_fd_sc_hd__clkbuf_1 _7559_ (.A(_3763_),
    .X(_0580_));
 sky130_fd_sc_hd__nand2_1 _7560_ (.A(net488),
    .B(_3390_),
    .Y(_3764_));
 sky130_fd_sc_hd__o21ai_1 _7561_ (.A1(_3684_),
    .A2(_3451_),
    .B1(_3764_),
    .Y(_0581_));
 sky130_fd_sc_hd__mux2_1 _7562_ (.A0(net658),
    .A1(_3462_),
    .S(_3762_),
    .X(_3765_));
 sky130_fd_sc_hd__clkbuf_1 _7563_ (.A(_3765_),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _7564_ (.A0(net687),
    .A1(_3472_),
    .S(_3762_),
    .X(_3766_));
 sky130_fd_sc_hd__clkbuf_1 _7565_ (.A(_3766_),
    .X(_0583_));
 sky130_fd_sc_hd__nor2_1 _7566_ (.A(net519),
    .B(_1113_),
    .Y(_3767_));
 sky130_fd_sc_hd__a21oi_1 _7567_ (.A1(\ks1.next_ready_o ),
    .A2(_3480_),
    .B1(_3767_),
    .Y(_0584_));
 sky130_fd_sc_hd__nor2_1 _7568_ (.A(net508),
    .B(_1113_),
    .Y(_3768_));
 sky130_fd_sc_hd__a21oi_1 _7569_ (.A1(\ks1.next_ready_o ),
    .A2(_3486_),
    .B1(_3768_),
    .Y(_0585_));
 sky130_fd_sc_hd__mux2_1 _7570_ (.A0(net695),
    .A1(_3496_),
    .S(_3762_),
    .X(_3769_));
 sky130_fd_sc_hd__clkbuf_1 _7571_ (.A(_3769_),
    .X(_0586_));
 sky130_fd_sc_hd__inv_2 _7572_ (.A(_3502_),
    .Y(_3770_));
 sky130_fd_sc_hd__mux2_1 _7573_ (.A0(net629),
    .A1(_3770_),
    .S(_3762_),
    .X(_3771_));
 sky130_fd_sc_hd__clkbuf_1 _7574_ (.A(_3771_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_1 _7575_ (.A0(net679),
    .A1(_3512_),
    .S(_3762_),
    .X(_3772_));
 sky130_fd_sc_hd__clkbuf_1 _7576_ (.A(_3772_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_1 _7577_ (.A0(net660),
    .A1(_3519_),
    .S(_3762_),
    .X(_3773_));
 sky130_fd_sc_hd__clkbuf_1 _7578_ (.A(_3773_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_1 _7579_ (.A0(net673),
    .A1(_3527_),
    .S(_3762_),
    .X(_3774_));
 sky130_fd_sc_hd__clkbuf_1 _7580_ (.A(_3774_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _7581_ (.A0(net668),
    .A1(_3535_),
    .S(_3762_),
    .X(_3775_));
 sky130_fd_sc_hd__clkbuf_1 _7582_ (.A(_3775_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _7583_ (.A0(\ks1.key_reg[115] ),
    .A1(_3543_),
    .S(_3762_),
    .X(_3776_));
 sky130_fd_sc_hd__clkbuf_1 _7584_ (.A(_3776_),
    .X(_0592_));
 sky130_fd_sc_hd__clkbuf_8 _7585_ (.A(_1112_),
    .X(_3777_));
 sky130_fd_sc_hd__mux2_1 _7586_ (.A0(\ks1.key_reg[116] ),
    .A1(_3551_),
    .S(_3777_),
    .X(_3778_));
 sky130_fd_sc_hd__clkbuf_1 _7587_ (.A(_3778_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _7588_ (.A0(net690),
    .A1(_3559_),
    .S(_3777_),
    .X(_3779_));
 sky130_fd_sc_hd__clkbuf_1 _7589_ (.A(_3779_),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _7590_ (.A0(net670),
    .A1(_3567_),
    .S(_3777_),
    .X(_3780_));
 sky130_fd_sc_hd__clkbuf_1 _7591_ (.A(_3780_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _7592_ (.A0(net659),
    .A1(_3575_),
    .S(_3777_),
    .X(_3781_));
 sky130_fd_sc_hd__clkbuf_1 _7593_ (.A(_3781_),
    .X(_0596_));
 sky130_fd_sc_hd__nand2_1 _7594_ (.A(net520),
    .B(_3390_),
    .Y(_3782_));
 sky130_fd_sc_hd__o21ai_1 _7595_ (.A1(_3684_),
    .A2(_3591_),
    .B1(_3782_),
    .Y(_0597_));
 sky130_fd_sc_hd__inv_2 _7596_ (.A(_3604_),
    .Y(_3783_));
 sky130_fd_sc_hd__mux2_1 _7597_ (.A0(net681),
    .A1(_3783_),
    .S(_3777_),
    .X(_3784_));
 sky130_fd_sc_hd__clkbuf_1 _7598_ (.A(_3784_),
    .X(_0598_));
 sky130_fd_sc_hd__inv_2 _7599_ (.A(_3617_),
    .Y(_3785_));
 sky130_fd_sc_hd__mux2_1 _7600_ (.A0(net685),
    .A1(_3785_),
    .S(_3777_),
    .X(_3786_));
 sky130_fd_sc_hd__clkbuf_1 _7601_ (.A(_3786_),
    .X(_0599_));
 sky130_fd_sc_hd__nor2_1 _7602_ (.A(net507),
    .B(_1113_),
    .Y(_3787_));
 sky130_fd_sc_hd__a21oi_1 _7603_ (.A1(\ks1.next_ready_o ),
    .A2(_3628_),
    .B1(_3787_),
    .Y(_0600_));
 sky130_fd_sc_hd__inv_2 _7604_ (.A(_3638_),
    .Y(_3788_));
 sky130_fd_sc_hd__mux2_1 _7605_ (.A0(\ks1.key_reg[124] ),
    .A1(_3788_),
    .S(_3777_),
    .X(_3789_));
 sky130_fd_sc_hd__clkbuf_1 _7606_ (.A(_3789_),
    .X(_0601_));
 sky130_fd_sc_hd__inv_2 _7607_ (.A(_3648_),
    .Y(_3790_));
 sky130_fd_sc_hd__mux2_1 _7608_ (.A0(net704),
    .A1(_3790_),
    .S(_3777_),
    .X(_3791_));
 sky130_fd_sc_hd__clkbuf_1 _7609_ (.A(_3791_),
    .X(_0602_));
 sky130_fd_sc_hd__inv_2 _7610_ (.A(_3658_),
    .Y(_3792_));
 sky130_fd_sc_hd__mux2_1 _7611_ (.A0(net691),
    .A1(_3792_),
    .S(_3777_),
    .X(_3793_));
 sky130_fd_sc_hd__clkbuf_1 _7612_ (.A(_3793_),
    .X(_0603_));
 sky130_fd_sc_hd__inv_2 _7613_ (.A(_3669_),
    .Y(_3794_));
 sky130_fd_sc_hd__mux2_1 _7614_ (.A0(\ks1.key_reg[127] ),
    .A1(_3794_),
    .S(_3777_),
    .X(_3795_));
 sky130_fd_sc_hd__clkbuf_1 _7615_ (.A(_3795_),
    .X(_0604_));
 sky130_fd_sc_hd__a21oi_1 _7616_ (.A1(_0679_),
    .A2(_1127_),
    .B1(_2527_),
    .Y(_3796_));
 sky130_fd_sc_hd__o21ba_1 _7617_ (.A1(\mix1.state[1] ),
    .A2(_3796_),
    .B1_N(\mix1.state[0] ),
    .X(_0605_));
 sky130_fd_sc_hd__or2_1 _7618_ (.A(_2642_),
    .B(_3010_),
    .X(_3797_));
 sky130_fd_sc_hd__clkbuf_1 _7619_ (.A(_3797_),
    .X(_0606_));
 sky130_fd_sc_hd__buf_4 _7620_ (.A(_2613_),
    .X(_3798_));
 sky130_fd_sc_hd__mux2_1 _7621_ (.A0(net538),
    .A1(_2641_),
    .S(_3798_),
    .X(_3799_));
 sky130_fd_sc_hd__clkbuf_1 _7622_ (.A(_3799_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_1 _7623_ (.A0(net542),
    .A1(_2709_),
    .S(_3798_),
    .X(_3800_));
 sky130_fd_sc_hd__clkbuf_1 _7624_ (.A(_3800_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _7625_ (.A0(net543),
    .A1(_2755_),
    .S(_3798_),
    .X(_3801_));
 sky130_fd_sc_hd__clkbuf_1 _7626_ (.A(_3801_),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _7627_ (.A0(net541),
    .A1(_2796_),
    .S(_3798_),
    .X(_3802_));
 sky130_fd_sc_hd__clkbuf_1 _7628_ (.A(_3802_),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _7629_ (.A0(net562),
    .A1(_2835_),
    .S(_3798_),
    .X(_3803_));
 sky130_fd_sc_hd__clkbuf_1 _7630_ (.A(_3803_),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _7631_ (.A0(net561),
    .A1(_2854_),
    .S(_3798_),
    .X(_3804_));
 sky130_fd_sc_hd__clkbuf_1 _7632_ (.A(_3804_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _7633_ (.A0(net551),
    .A1(_2864_),
    .S(_3798_),
    .X(_3805_));
 sky130_fd_sc_hd__clkbuf_1 _7634_ (.A(_3805_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _7635_ (.A0(net563),
    .A1(_2874_),
    .S(_3798_),
    .X(_3806_));
 sky130_fd_sc_hd__clkbuf_1 _7636_ (.A(_3806_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _7637_ (.A0(net539),
    .A1(_2883_),
    .S(_3798_),
    .X(_3807_));
 sky130_fd_sc_hd__clkbuf_1 _7638_ (.A(_3807_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _7639_ (.A0(net537),
    .A1(_2896_),
    .S(_3798_),
    .X(_3808_));
 sky130_fd_sc_hd__clkbuf_1 _7640_ (.A(_3808_),
    .X(_0616_));
 sky130_fd_sc_hd__buf_4 _7641_ (.A(_2613_),
    .X(_3809_));
 sky130_fd_sc_hd__mux2_1 _7642_ (.A0(net564),
    .A1(_2907_),
    .S(_3809_),
    .X(_3810_));
 sky130_fd_sc_hd__clkbuf_1 _7643_ (.A(_3810_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _7644_ (.A0(net574),
    .A1(_2918_),
    .S(_3809_),
    .X(_3811_));
 sky130_fd_sc_hd__clkbuf_1 _7645_ (.A(_3811_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _7646_ (.A0(net598),
    .A1(_2928_),
    .S(_3809_),
    .X(_3812_));
 sky130_fd_sc_hd__clkbuf_1 _7647_ (.A(_3812_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_1 _7648_ (.A0(net590),
    .A1(_2939_),
    .S(_3809_),
    .X(_3813_));
 sky130_fd_sc_hd__clkbuf_1 _7649_ (.A(_3813_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _7650_ (.A0(net706),
    .A1(_2948_),
    .S(_3809_),
    .X(_3814_));
 sky130_fd_sc_hd__clkbuf_1 _7651_ (.A(_3814_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_1 _7652_ (.A0(net627),
    .A1(_2954_),
    .S(_3809_),
    .X(_3815_));
 sky130_fd_sc_hd__clkbuf_1 _7653_ (.A(_3815_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_1 _7654_ (.A0(net569),
    .A1(_2958_),
    .S(_3809_),
    .X(_3816_));
 sky130_fd_sc_hd__clkbuf_1 _7655_ (.A(_3816_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_1 _7656_ (.A0(net571),
    .A1(_2962_),
    .S(_3809_),
    .X(_3817_));
 sky130_fd_sc_hd__clkbuf_1 _7657_ (.A(_3817_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_1 _7658_ (.A0(net592),
    .A1(_2964_),
    .S(_3809_),
    .X(_3818_));
 sky130_fd_sc_hd__clkbuf_1 _7659_ (.A(_3818_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_1 _7660_ (.A0(net622),
    .A1(_2968_),
    .S(_3809_),
    .X(_3819_));
 sky130_fd_sc_hd__clkbuf_1 _7661_ (.A(_3819_),
    .X(_0626_));
 sky130_fd_sc_hd__buf_4 _7662_ (.A(_2613_),
    .X(_3820_));
 sky130_fd_sc_hd__mux2_1 _7663_ (.A0(net570),
    .A1(_2973_),
    .S(_3820_),
    .X(_3821_));
 sky130_fd_sc_hd__clkbuf_1 _7664_ (.A(_3821_),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _7665_ (.A0(net526),
    .A1(_2976_),
    .S(_3820_),
    .X(_3822_));
 sky130_fd_sc_hd__clkbuf_1 _7666_ (.A(_3822_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _7667_ (.A0(net610),
    .A1(_2978_),
    .S(_3820_),
    .X(_3823_));
 sky130_fd_sc_hd__clkbuf_1 _7668_ (.A(_3823_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _7669_ (.A0(net616),
    .A1(_2981_),
    .S(_3820_),
    .X(_3824_));
 sky130_fd_sc_hd__clkbuf_1 _7670_ (.A(_3824_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _7671_ (.A0(net575),
    .A1(_2985_),
    .S(_3820_),
    .X(_3825_));
 sky130_fd_sc_hd__clkbuf_1 _7672_ (.A(_3825_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _7673_ (.A0(net595),
    .A1(_2987_),
    .S(_3820_),
    .X(_3826_));
 sky130_fd_sc_hd__clkbuf_1 _7674_ (.A(_3826_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _7675_ (.A0(net580),
    .A1(_2992_),
    .S(_3820_),
    .X(_3827_));
 sky130_fd_sc_hd__clkbuf_1 _7676_ (.A(_3827_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _7677_ (.A0(net567),
    .A1(_2996_),
    .S(_3820_),
    .X(_3828_));
 sky130_fd_sc_hd__clkbuf_1 _7678_ (.A(_3828_),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _7679_ (.A0(net593),
    .A1(_2998_),
    .S(_3820_),
    .X(_3829_));
 sky130_fd_sc_hd__clkbuf_1 _7680_ (.A(_3829_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _7681_ (.A0(net586),
    .A1(_3000_),
    .S(_3820_),
    .X(_3830_));
 sky130_fd_sc_hd__clkbuf_1 _7682_ (.A(_3830_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _7683_ (.A0(net540),
    .A1(_3004_),
    .S(_2613_),
    .X(_3831_));
 sky130_fd_sc_hd__clkbuf_1 _7684_ (.A(_3831_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _7685_ (.A0(net581),
    .A1(_3008_),
    .S(_2613_),
    .X(_3832_));
 sky130_fd_sc_hd__clkbuf_1 _7686_ (.A(_3832_),
    .X(_0638_));
 sky130_fd_sc_hd__nor2_2 _7687_ (.A(_2491_),
    .B(_0958_),
    .Y(_3833_));
 sky130_fd_sc_hd__a22o_1 _7688_ (.A1(\sub1.data_o[40] ),
    .A2(_3127_),
    .B1(_3833_),
    .B2(\sub1.data_o[104] ),
    .X(_3834_));
 sky130_fd_sc_hd__a31o_1 _7689_ (.A1(_3339_),
    .A2(_0958_),
    .A3(_1213_),
    .B1(_3834_),
    .X(_0639_));
 sky130_fd_sc_hd__a22o_1 _7690_ (.A1(\sub1.data_o[41] ),
    .A2(_3127_),
    .B1(_3833_),
    .B2(\sub1.data_o[105] ),
    .X(_3835_));
 sky130_fd_sc_hd__a31o_1 _7691_ (.A1(_3339_),
    .A2(_0958_),
    .A3(_1247_),
    .B1(_3835_),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _7692_ (.A1(\sub1.data_o[42] ),
    .A2(_3055_),
    .B1(_3833_),
    .B2(\sub1.data_o[106] ),
    .X(_3836_));
 sky130_fd_sc_hd__a31o_1 _7693_ (.A1(_3339_),
    .A2(_0958_),
    .A3(_1257_),
    .B1(_3836_),
    .X(_0641_));
 sky130_fd_sc_hd__a22o_1 _7694_ (.A1(\sub1.data_o[43] ),
    .A2(_3055_),
    .B1(_3833_),
    .B2(\sub1.data_o[107] ),
    .X(_3837_));
 sky130_fd_sc_hd__a31o_1 _7695_ (.A1(_3339_),
    .A2(_0958_),
    .A3(_1272_),
    .B1(_3837_),
    .X(_0642_));
 sky130_fd_sc_hd__a22o_1 _7696_ (.A1(\sub1.data_o[44] ),
    .A2(_3055_),
    .B1(_3833_),
    .B2(\sub1.data_o[108] ),
    .X(_3838_));
 sky130_fd_sc_hd__a31o_1 _7697_ (.A1(_3339_),
    .A2(_0958_),
    .A3(_1278_),
    .B1(_3838_),
    .X(_0643_));
 sky130_fd_sc_hd__a22o_1 _7698_ (.A1(\sub1.data_o[45] ),
    .A2(_3055_),
    .B1(_3833_),
    .B2(\sub1.data_o[109] ),
    .X(_3839_));
 sky130_fd_sc_hd__a31o_1 _7699_ (.A1(_3339_),
    .A2(_0958_),
    .A3(_1286_),
    .B1(_3839_),
    .X(_0644_));
 sky130_fd_sc_hd__a22o_1 _7700_ (.A1(\sub1.data_o[46] ),
    .A2(_3055_),
    .B1(_3833_),
    .B2(\sub1.data_o[110] ),
    .X(_3840_));
 sky130_fd_sc_hd__a31o_1 _7701_ (.A1(_1139_),
    .A2(_0958_),
    .A3(_1293_),
    .B1(_3840_),
    .X(_0645_));
 sky130_fd_sc_hd__a22o_1 _7702_ (.A1(\sub1.data_o[47] ),
    .A2(_3055_),
    .B1(_3833_),
    .B2(\sub1.data_o[111] ),
    .X(_3841_));
 sky130_fd_sc_hd__a31o_1 _7703_ (.A1(_1139_),
    .A2(_0958_),
    .A3(_1300_),
    .B1(_3841_),
    .X(_0646_));
 sky130_fd_sc_hd__nor2_1 _7704_ (.A(\ks1.state[2] ),
    .B(\ks1.state[0] ),
    .Y(_3842_));
 sky130_fd_sc_hd__o21a_1 _7705_ (.A1(net528),
    .A2(_0751_),
    .B1(_3842_),
    .X(_0647_));
 sky130_fd_sc_hd__or2_1 _7706_ (.A(_0850_),
    .B(_0974_),
    .X(_3843_));
 sky130_fd_sc_hd__clkbuf_1 _7707_ (.A(_3843_),
    .X(_0648_));
 sky130_fd_sc_hd__dfrtp_4 _7708_ (.CLK(clknet_leaf_72_clk),
    .D(_0000_),
    .RESET_B(net412),
    .Q(\addroundkey_round[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7709_ (.CLK(clknet_leaf_71_clk),
    .D(_0001_),
    .RESET_B(net412),
    .Q(\addroundkey_round[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7710_ (.CLK(clknet_leaf_72_clk),
    .D(_0002_),
    .RESET_B(net412),
    .Q(\addroundkey_round[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7711_ (.CLK(clknet_leaf_70_clk),
    .D(_0003_),
    .RESET_B(net413),
    .Q(\addroundkey_round[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7712_ (.CLK(clknet_leaf_19_clk),
    .D(next_ready_o),
    .RESET_B(net449),
    .Q(net388));
 sky130_fd_sc_hd__dfrtp_4 _7713_ (.CLK(clknet_leaf_82_clk),
    .D(next_state),
    .RESET_B(net391),
    .Q(state));
 sky130_fd_sc_hd__dfrtp_4 _7714_ (.CLK(clknet_leaf_23_clk),
    .D(_0004_),
    .RESET_B(net452),
    .Q(\sub1.data_o[112] ));
 sky130_fd_sc_hd__dfrtp_4 _7715_ (.CLK(clknet_leaf_35_clk),
    .D(_0005_),
    .RESET_B(net473),
    .Q(\sub1.data_o[113] ));
 sky130_fd_sc_hd__dfrtp_4 _7716_ (.CLK(clknet_leaf_35_clk),
    .D(_0006_),
    .RESET_B(net473),
    .Q(\sub1.data_o[114] ));
 sky130_fd_sc_hd__dfrtp_4 _7717_ (.CLK(clknet_leaf_23_clk),
    .D(_0007_),
    .RESET_B(net452),
    .Q(\sub1.data_o[115] ));
 sky130_fd_sc_hd__dfrtp_4 _7718_ (.CLK(clknet_leaf_36_clk),
    .D(_0008_),
    .RESET_B(net474),
    .Q(\sub1.data_o[116] ));
 sky130_fd_sc_hd__dfrtp_4 _7719_ (.CLK(clknet_leaf_36_clk),
    .D(_0009_),
    .RESET_B(net473),
    .Q(\sub1.data_o[117] ));
 sky130_fd_sc_hd__dfrtp_4 _7720_ (.CLK(clknet_leaf_24_clk),
    .D(_0010_),
    .RESET_B(net474),
    .Q(\sub1.data_o[118] ));
 sky130_fd_sc_hd__dfrtp_4 _7721_ (.CLK(clknet_leaf_34_clk),
    .D(_0011_),
    .RESET_B(net474),
    .Q(\sub1.data_o[119] ));
 sky130_fd_sc_hd__dfrtp_1 _7722_ (.CLK(clknet_leaf_84_clk),
    .D(_0012_),
    .RESET_B(net391),
    .Q(\round[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7723_ (.CLK(clknet_leaf_84_clk),
    .D(_0013_),
    .RESET_B(net391),
    .Q(\round[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7724_ (.CLK(clknet_leaf_82_clk),
    .D(_0014_),
    .RESET_B(net391),
    .Q(\round[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7725_ (.CLK(clknet_leaf_81_clk),
    .D(_0015_),
    .RESET_B(net390),
    .Q(\round[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7726_ (.CLK(clknet_leaf_82_clk),
    .D(next_addroundkey_ready_o),
    .RESET_B(net391),
    .Q(addroundkey_ready_o));
 sky130_fd_sc_hd__dfrtp_4 _7727_ (.CLK(clknet_leaf_84_clk),
    .D(next_addroundkey_start_i),
    .RESET_B(net391),
    .Q(addroundkey_start_i));
 sky130_fd_sc_hd__dfrtp_4 _7728_ (.CLK(clknet_leaf_57_clk),
    .D(_0016_),
    .RESET_B(net428),
    .Q(net260));
 sky130_fd_sc_hd__dfrtp_4 _7729_ (.CLK(clknet_leaf_54_clk),
    .D(_0017_),
    .RESET_B(net458),
    .Q(net299));
 sky130_fd_sc_hd__dfrtp_4 _7730_ (.CLK(clknet_leaf_8_clk),
    .D(_0018_),
    .RESET_B(net410),
    .Q(net310));
 sky130_fd_sc_hd__dfrtp_4 _7731_ (.CLK(clknet_leaf_8_clk),
    .D(_0019_),
    .RESET_B(net410),
    .Q(net321));
 sky130_fd_sc_hd__dfrtp_4 _7732_ (.CLK(clknet_leaf_81_clk),
    .D(_0020_),
    .RESET_B(net390),
    .Q(net332));
 sky130_fd_sc_hd__dfrtp_4 _7733_ (.CLK(clknet_leaf_53_clk),
    .D(_0021_),
    .RESET_B(net458),
    .Q(net343));
 sky130_fd_sc_hd__dfrtp_4 _7734_ (.CLK(clknet_leaf_9_clk),
    .D(_0022_),
    .RESET_B(net443),
    .Q(net354));
 sky130_fd_sc_hd__dfrtp_4 _7735_ (.CLK(clknet_leaf_5_clk),
    .D(_0023_),
    .RESET_B(net410),
    .Q(net365));
 sky130_fd_sc_hd__dfrtp_4 _7736_ (.CLK(clknet_leaf_8_clk),
    .D(_0024_),
    .RESET_B(net443),
    .Q(net376));
 sky130_fd_sc_hd__dfrtp_4 _7737_ (.CLK(clknet_leaf_50_clk),
    .D(_0025_),
    .RESET_B(net459),
    .Q(net387));
 sky130_fd_sc_hd__dfrtp_4 _7738_ (.CLK(clknet_leaf_51_clk),
    .D(_0026_),
    .RESET_B(net463),
    .Q(net271));
 sky130_fd_sc_hd__dfrtp_4 _7739_ (.CLK(clknet_leaf_48_clk),
    .D(_0027_),
    .RESET_B(net461),
    .Q(net282));
 sky130_fd_sc_hd__dfrtp_4 _7740_ (.CLK(clknet_leaf_50_clk),
    .D(_0028_),
    .RESET_B(net459),
    .Q(net291));
 sky130_fd_sc_hd__dfrtp_4 _7741_ (.CLK(clknet_leaf_47_clk),
    .D(_0029_),
    .RESET_B(net461),
    .Q(net292));
 sky130_fd_sc_hd__dfrtp_4 _7742_ (.CLK(clknet_leaf_48_clk),
    .D(_0030_),
    .RESET_B(net461),
    .Q(net293));
 sky130_fd_sc_hd__dfrtp_4 _7743_ (.CLK(clknet_leaf_47_clk),
    .D(_0031_),
    .RESET_B(net462),
    .Q(net294));
 sky130_fd_sc_hd__dfrtp_4 _7744_ (.CLK(clknet_leaf_51_clk),
    .D(_0032_),
    .RESET_B(net463),
    .Q(net295));
 sky130_fd_sc_hd__dfrtp_4 _7745_ (.CLK(clknet_leaf_52_clk),
    .D(_0033_),
    .RESET_B(net463),
    .Q(net296));
 sky130_fd_sc_hd__dfrtp_4 _7746_ (.CLK(clknet_leaf_52_clk),
    .D(_0034_),
    .RESET_B(net463),
    .Q(net297));
 sky130_fd_sc_hd__dfrtp_4 _7747_ (.CLK(clknet_leaf_47_clk),
    .D(_0035_),
    .RESET_B(net465),
    .Q(net298));
 sky130_fd_sc_hd__dfrtp_4 _7748_ (.CLK(clknet_leaf_52_clk),
    .D(_0036_),
    .RESET_B(net456),
    .Q(net300));
 sky130_fd_sc_hd__dfrtp_4 _7749_ (.CLK(clknet_leaf_52_clk),
    .D(_0037_),
    .RESET_B(net463),
    .Q(net301));
 sky130_fd_sc_hd__dfrtp_4 _7750_ (.CLK(clknet_leaf_46_clk),
    .D(_0038_),
    .RESET_B(net465),
    .Q(net302));
 sky130_fd_sc_hd__dfrtp_4 _7751_ (.CLK(clknet_leaf_52_clk),
    .D(_0039_),
    .RESET_B(net456),
    .Q(net303));
 sky130_fd_sc_hd__dfrtp_4 _7752_ (.CLK(clknet_leaf_61_clk),
    .D(_0040_),
    .RESET_B(net428),
    .Q(net304));
 sky130_fd_sc_hd__dfrtp_4 _7753_ (.CLK(clknet_leaf_61_clk),
    .D(_0041_),
    .RESET_B(net428),
    .Q(net305));
 sky130_fd_sc_hd__dfrtp_4 _7754_ (.CLK(clknet_leaf_62_clk),
    .D(_0042_),
    .RESET_B(net430),
    .Q(net306));
 sky130_fd_sc_hd__dfrtp_4 _7755_ (.CLK(clknet_leaf_51_clk),
    .D(_0043_),
    .RESET_B(net459),
    .Q(net307));
 sky130_fd_sc_hd__dfrtp_4 _7756_ (.CLK(clknet_leaf_62_clk),
    .D(_0044_),
    .RESET_B(net430),
    .Q(net308));
 sky130_fd_sc_hd__dfrtp_4 _7757_ (.CLK(clknet_leaf_51_clk),
    .D(_0045_),
    .RESET_B(net459),
    .Q(net309));
 sky130_fd_sc_hd__dfrtp_4 _7758_ (.CLK(clknet_leaf_48_clk),
    .D(_0046_),
    .RESET_B(net461),
    .Q(net311));
 sky130_fd_sc_hd__dfrtp_4 _7759_ (.CLK(clknet_leaf_63_clk),
    .D(_0047_),
    .RESET_B(net426),
    .Q(net312));
 sky130_fd_sc_hd__dfrtp_4 _7760_ (.CLK(clknet_leaf_7_clk),
    .D(_0048_),
    .RESET_B(net408),
    .Q(net313));
 sky130_fd_sc_hd__dfrtp_4 _7761_ (.CLK(clknet_leaf_63_clk),
    .D(_0049_),
    .RESET_B(net426),
    .Q(net314));
 sky130_fd_sc_hd__dfrtp_2 _7762_ (.CLK(clknet_leaf_8_clk),
    .D(_0050_),
    .RESET_B(net410),
    .Q(net315));
 sky130_fd_sc_hd__dfrtp_4 _7763_ (.CLK(clknet_leaf_10_clk),
    .D(_0051_),
    .RESET_B(net443),
    .Q(net316));
 sky130_fd_sc_hd__dfrtp_4 _7764_ (.CLK(clknet_leaf_80_clk),
    .D(_0052_),
    .RESET_B(net408),
    .Q(net317));
 sky130_fd_sc_hd__dfrtp_4 _7765_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0053_),
    .RESET_B(net457),
    .Q(net318));
 sky130_fd_sc_hd__dfrtp_4 _7766_ (.CLK(clknet_leaf_29_clk),
    .D(_0054_),
    .RESET_B(net457),
    .Q(net319));
 sky130_fd_sc_hd__dfrtp_4 _7767_ (.CLK(clknet_leaf_52_clk),
    .D(_0055_),
    .RESET_B(net464),
    .Q(net320));
 sky130_fd_sc_hd__dfrtp_4 _7768_ (.CLK(clknet_leaf_50_clk),
    .D(_0056_),
    .RESET_B(net459),
    .Q(net322));
 sky130_fd_sc_hd__dfrtp_4 _7769_ (.CLK(clknet_leaf_50_clk),
    .D(_0057_),
    .RESET_B(net460),
    .Q(net323));
 sky130_fd_sc_hd__dfrtp_4 _7770_ (.CLK(clknet_leaf_51_clk),
    .D(_0058_),
    .RESET_B(net460),
    .Q(net324));
 sky130_fd_sc_hd__dfrtp_4 _7771_ (.CLK(clknet_leaf_50_clk),
    .D(_0059_),
    .RESET_B(net459),
    .Q(net325));
 sky130_fd_sc_hd__dfrtp_4 _7772_ (.CLK(clknet_leaf_61_clk),
    .D(_0060_),
    .RESET_B(net429),
    .Q(net326));
 sky130_fd_sc_hd__dfrtp_4 _7773_ (.CLK(clknet_leaf_53_clk),
    .D(_0061_),
    .RESET_B(net458),
    .Q(net327));
 sky130_fd_sc_hd__dfrtp_4 _7774_ (.CLK(clknet_leaf_57_clk),
    .D(_0062_),
    .RESET_B(net423),
    .Q(net328));
 sky130_fd_sc_hd__dfrtp_4 _7775_ (.CLK(clknet_leaf_51_clk),
    .D(_0063_),
    .RESET_B(net460),
    .Q(net329));
 sky130_fd_sc_hd__dfrtp_4 _7776_ (.CLK(clknet_leaf_30_clk),
    .D(_0064_),
    .RESET_B(net456),
    .Q(net330));
 sky130_fd_sc_hd__dfrtp_4 _7777_ (.CLK(clknet_leaf_31_clk),
    .D(_0065_),
    .RESET_B(net470),
    .Q(net331));
 sky130_fd_sc_hd__dfrtp_4 _7778_ (.CLK(clknet_leaf_47_clk),
    .D(_0066_),
    .RESET_B(net465),
    .Q(net333));
 sky130_fd_sc_hd__dfrtp_4 _7779_ (.CLK(clknet_leaf_43_clk),
    .D(_0067_),
    .RESET_B(net479),
    .Q(net334));
 sky130_fd_sc_hd__dfrtp_4 _7780_ (.CLK(clknet_leaf_31_clk),
    .D(_0068_),
    .RESET_B(net456),
    .Q(net335));
 sky130_fd_sc_hd__dfrtp_4 _7781_ (.CLK(clknet_leaf_39_clk),
    .D(_0069_),
    .RESET_B(net470),
    .Q(net336));
 sky130_fd_sc_hd__dfrtp_4 _7782_ (.CLK(clknet_leaf_45_clk),
    .D(_0070_),
    .RESET_B(net477),
    .Q(net337));
 sky130_fd_sc_hd__dfrtp_4 _7783_ (.CLK(clknet_leaf_39_clk),
    .D(_0071_),
    .RESET_B(net477),
    .Q(net338));
 sky130_fd_sc_hd__dfrtp_4 _7784_ (.CLK(clknet_leaf_57_clk),
    .D(_0072_),
    .RESET_B(net423),
    .Q(net339));
 sky130_fd_sc_hd__dfrtp_4 _7785_ (.CLK(clknet_leaf_60_clk),
    .D(_0073_),
    .RESET_B(net424),
    .Q(net340));
 sky130_fd_sc_hd__dfrtp_4 _7786_ (.CLK(clknet_leaf_63_clk),
    .D(_0074_),
    .RESET_B(net427),
    .Q(net341));
 sky130_fd_sc_hd__dfrtp_4 _7787_ (.CLK(clknet_leaf_57_clk),
    .D(_0075_),
    .RESET_B(net423),
    .Q(net342));
 sky130_fd_sc_hd__dfrtp_4 _7788_ (.CLK(clknet_leaf_75_clk),
    .D(_0076_),
    .RESET_B(net421),
    .Q(net344));
 sky130_fd_sc_hd__dfrtp_4 _7789_ (.CLK(clknet_leaf_60_clk),
    .D(_0077_),
    .RESET_B(net428),
    .Q(net345));
 sky130_fd_sc_hd__dfrtp_4 _7790_ (.CLK(clknet_leaf_64_clk),
    .D(_0078_),
    .RESET_B(net426),
    .Q(net346));
 sky130_fd_sc_hd__dfrtp_4 _7791_ (.CLK(clknet_leaf_58_clk),
    .D(_0079_),
    .RESET_B(net421),
    .Q(net347));
 sky130_fd_sc_hd__dfrtp_4 _7792_ (.CLK(clknet_leaf_75_clk),
    .D(_0080_),
    .RESET_B(net421),
    .Q(net348));
 sky130_fd_sc_hd__dfrtp_4 _7793_ (.CLK(clknet_leaf_58_clk),
    .D(_0081_),
    .RESET_B(net423),
    .Q(net349));
 sky130_fd_sc_hd__dfrtp_4 _7794_ (.CLK(clknet_leaf_48_clk),
    .D(_0082_),
    .RESET_B(net461),
    .Q(net350));
 sky130_fd_sc_hd__dfrtp_4 _7795_ (.CLK(clknet_leaf_53_clk),
    .D(_0083_),
    .RESET_B(net459),
    .Q(net351));
 sky130_fd_sc_hd__dfrtp_4 _7796_ (.CLK(clknet_leaf_64_clk),
    .D(_0084_),
    .RESET_B(net426),
    .Q(net352));
 sky130_fd_sc_hd__dfrtp_4 _7797_ (.CLK(clknet_leaf_74_clk),
    .D(_0085_),
    .RESET_B(net414),
    .Q(net353));
 sky130_fd_sc_hd__dfrtp_4 _7798_ (.CLK(clknet_leaf_51_clk),
    .D(_0086_),
    .RESET_B(net463),
    .Q(net355));
 sky130_fd_sc_hd__dfrtp_4 _7799_ (.CLK(clknet_leaf_62_clk),
    .D(_0087_),
    .RESET_B(net430),
    .Q(net356));
 sky130_fd_sc_hd__dfrtp_4 _7800_ (.CLK(clknet_leaf_62_clk),
    .D(_0088_),
    .RESET_B(net430),
    .Q(net357));
 sky130_fd_sc_hd__dfrtp_4 _7801_ (.CLK(clknet_leaf_62_clk),
    .D(_0089_),
    .RESET_B(net431),
    .Q(net358));
 sky130_fd_sc_hd__dfrtp_4 _7802_ (.CLK(clknet_leaf_52_clk),
    .D(_0090_),
    .RESET_B(net463),
    .Q(net359));
 sky130_fd_sc_hd__dfrtp_4 _7803_ (.CLK(clknet_leaf_61_clk),
    .D(_0091_),
    .RESET_B(net429),
    .Q(net360));
 sky130_fd_sc_hd__dfrtp_4 _7804_ (.CLK(clknet_leaf_76_clk),
    .D(_0092_),
    .RESET_B(net421),
    .Q(net361));
 sky130_fd_sc_hd__dfrtp_4 _7805_ (.CLK(clknet_leaf_64_clk),
    .D(_0093_),
    .RESET_B(net427),
    .Q(net362));
 sky130_fd_sc_hd__dfrtp_4 _7806_ (.CLK(clknet_leaf_66_clk),
    .D(_0094_),
    .RESET_B(net418),
    .Q(net363));
 sky130_fd_sc_hd__dfrtp_4 _7807_ (.CLK(clknet_leaf_59_clk),
    .D(_0095_),
    .RESET_B(net424),
    .Q(net364));
 sky130_fd_sc_hd__dfrtp_4 _7808_ (.CLK(clknet_leaf_23_clk),
    .D(_0096_),
    .RESET_B(net452),
    .Q(net366));
 sky130_fd_sc_hd__dfrtp_4 _7809_ (.CLK(clknet_leaf_40_clk),
    .D(_0097_),
    .RESET_B(net478),
    .Q(net367));
 sky130_fd_sc_hd__dfrtp_4 _7810_ (.CLK(clknet_leaf_39_clk),
    .D(_0098_),
    .RESET_B(net478),
    .Q(net368));
 sky130_fd_sc_hd__dfrtp_4 _7811_ (.CLK(clknet_leaf_40_clk),
    .D(_0099_),
    .RESET_B(net478),
    .Q(net369));
 sky130_fd_sc_hd__dfrtp_4 _7812_ (.CLK(clknet_leaf_79_clk),
    .D(_0100_),
    .RESET_B(net409),
    .Q(net370));
 sky130_fd_sc_hd__dfrtp_4 _7813_ (.CLK(clknet_leaf_39_clk),
    .D(_0101_),
    .RESET_B(net477),
    .Q(net371));
 sky130_fd_sc_hd__dfrtp_4 _7814_ (.CLK(clknet_leaf_34_clk),
    .D(_0102_),
    .RESET_B(net469),
    .Q(net372));
 sky130_fd_sc_hd__dfrtp_4 _7815_ (.CLK(clknet_leaf_35_clk),
    .D(_0103_),
    .RESET_B(net473),
    .Q(net373));
 sky130_fd_sc_hd__dfrtp_4 _7816_ (.CLK(clknet_leaf_79_clk),
    .D(_0104_),
    .RESET_B(net409),
    .Q(net374));
 sky130_fd_sc_hd__dfrtp_4 _7817_ (.CLK(clknet_leaf_73_clk),
    .D(_0105_),
    .RESET_B(net414),
    .Q(net375));
 sky130_fd_sc_hd__dfrtp_2 _7818_ (.CLK(clknet_leaf_84_clk),
    .D(_0106_),
    .RESET_B(net391),
    .Q(net377));
 sky130_fd_sc_hd__dfrtp_4 _7819_ (.CLK(clknet_leaf_74_clk),
    .D(_0107_),
    .RESET_B(net414),
    .Q(net378));
 sky130_fd_sc_hd__dfrtp_4 _7820_ (.CLK(clknet_leaf_74_clk),
    .D(_0108_),
    .RESET_B(net414),
    .Q(net379));
 sky130_fd_sc_hd__dfrtp_4 _7821_ (.CLK(clknet_leaf_72_clk),
    .D(_0109_),
    .RESET_B(net414),
    .Q(net380));
 sky130_fd_sc_hd__dfrtp_4 _7822_ (.CLK(clknet_leaf_79_clk),
    .D(_0110_),
    .RESET_B(net409),
    .Q(net381));
 sky130_fd_sc_hd__dfrtp_4 _7823_ (.CLK(clknet_leaf_84_clk),
    .D(_0111_),
    .RESET_B(net391),
    .Q(net382));
 sky130_fd_sc_hd__dfrtp_4 _7824_ (.CLK(clknet_leaf_22_clk),
    .D(_0112_),
    .RESET_B(net452),
    .Q(net383));
 sky130_fd_sc_hd__dfrtp_4 _7825_ (.CLK(clknet_leaf_22_clk),
    .D(_0113_),
    .RESET_B(net452),
    .Q(net384));
 sky130_fd_sc_hd__dfrtp_4 _7826_ (.CLK(clknet_leaf_36_clk),
    .D(_0114_),
    .RESET_B(net476),
    .Q(net385));
 sky130_fd_sc_hd__dfrtp_4 _7827_ (.CLK(clknet_leaf_21_clk),
    .D(_0115_),
    .RESET_B(net453),
    .Q(net386));
 sky130_fd_sc_hd__dfrtp_4 _7828_ (.CLK(clknet_leaf_86_clk),
    .D(_0116_),
    .RESET_B(net390),
    .Q(net261));
 sky130_fd_sc_hd__dfrtp_4 _7829_ (.CLK(clknet_leaf_86_clk),
    .D(_0117_),
    .RESET_B(net390),
    .Q(net262));
 sky130_fd_sc_hd__dfrtp_4 _7830_ (.CLK(clknet_leaf_22_clk),
    .D(_0118_),
    .RESET_B(net453),
    .Q(net263));
 sky130_fd_sc_hd__dfrtp_4 _7831_ (.CLK(clknet_leaf_21_clk),
    .D(_0119_),
    .RESET_B(net453),
    .Q(net264));
 sky130_fd_sc_hd__dfrtp_4 _7832_ (.CLK(clknet_leaf_58_clk),
    .D(_0120_),
    .RESET_B(net422),
    .Q(net265));
 sky130_fd_sc_hd__dfrtp_4 _7833_ (.CLK(clknet_leaf_58_clk),
    .D(_0121_),
    .RESET_B(net421),
    .Q(net266));
 sky130_fd_sc_hd__dfrtp_4 _7834_ (.CLK(clknet_leaf_7_clk),
    .D(_0122_),
    .RESET_B(net408),
    .Q(net267));
 sky130_fd_sc_hd__dfrtp_4 _7835_ (.CLK(clknet_leaf_7_clk),
    .D(_0123_),
    .RESET_B(net408),
    .Q(net268));
 sky130_fd_sc_hd__dfrtp_4 _7836_ (.CLK(clknet_leaf_80_clk),
    .D(_0124_),
    .RESET_B(net408),
    .Q(net269));
 sky130_fd_sc_hd__dfrtp_4 _7837_ (.CLK(clknet_leaf_76_clk),
    .D(_0125_),
    .RESET_B(net422),
    .Q(net270));
 sky130_fd_sc_hd__dfrtp_4 _7838_ (.CLK(clknet_leaf_65_clk),
    .D(_0126_),
    .RESET_B(net424),
    .Q(net272));
 sky130_fd_sc_hd__dfrtp_4 _7839_ (.CLK(clknet_leaf_80_clk),
    .D(_0127_),
    .RESET_B(net408),
    .Q(net273));
 sky130_fd_sc_hd__dfrtp_4 _7840_ (.CLK(clknet_leaf_80_clk),
    .D(_0128_),
    .RESET_B(net409),
    .Q(net274));
 sky130_fd_sc_hd__dfrtp_4 _7841_ (.CLK(clknet_leaf_23_clk),
    .D(_0129_),
    .RESET_B(net452),
    .Q(net275));
 sky130_fd_sc_hd__dfrtp_4 _7842_ (.CLK(clknet_leaf_22_clk),
    .D(_0130_),
    .RESET_B(net453),
    .Q(net276));
 sky130_fd_sc_hd__dfrtp_4 _7843_ (.CLK(clknet_leaf_40_clk),
    .D(_0131_),
    .RESET_B(net480),
    .Q(net277));
 sky130_fd_sc_hd__dfrtp_4 _7844_ (.CLK(clknet_leaf_22_clk),
    .D(_0132_),
    .RESET_B(net452),
    .Q(net278));
 sky130_fd_sc_hd__dfrtp_4 _7845_ (.CLK(clknet_leaf_44_clk),
    .D(_0133_),
    .RESET_B(net477),
    .Q(net279));
 sky130_fd_sc_hd__dfrtp_4 _7846_ (.CLK(clknet_leaf_22_clk),
    .D(_0134_),
    .RESET_B(net453),
    .Q(net280));
 sky130_fd_sc_hd__dfrtp_4 _7847_ (.CLK(clknet_leaf_51_clk),
    .D(_0135_),
    .RESET_B(net463),
    .Q(net281));
 sky130_fd_sc_hd__dfrtp_4 _7848_ (.CLK(clknet_leaf_81_clk),
    .D(_0136_),
    .RESET_B(net390),
    .Q(net283));
 sky130_fd_sc_hd__dfrtp_4 _7849_ (.CLK(clknet_leaf_74_clk),
    .D(_0137_),
    .RESET_B(net414),
    .Q(net284));
 sky130_fd_sc_hd__dfrtp_4 _7850_ (.CLK(clknet_leaf_86_clk),
    .D(_0138_),
    .RESET_B(net390),
    .Q(net285));
 sky130_fd_sc_hd__dfrtp_4 _7851_ (.CLK(clknet_leaf_83_clk),
    .D(_0139_),
    .RESET_B(net391),
    .Q(net286));
 sky130_fd_sc_hd__dfrtp_4 _7852_ (.CLK(clknet_leaf_83_clk),
    .D(_0140_),
    .RESET_B(net392),
    .Q(net287));
 sky130_fd_sc_hd__dfrtp_4 _7853_ (.CLK(clknet_leaf_75_clk),
    .D(_0141_),
    .RESET_B(net418),
    .Q(net288));
 sky130_fd_sc_hd__dfrtp_4 _7854_ (.CLK(clknet_leaf_83_clk),
    .D(_0142_),
    .RESET_B(net392),
    .Q(net289));
 sky130_fd_sc_hd__dfrtp_4 _7855_ (.CLK(clknet_leaf_81_clk),
    .D(_0143_),
    .RESET_B(net390),
    .Q(net290));
 sky130_fd_sc_hd__dfrtp_1 _7856_ (.CLK(clknet_leaf_82_clk),
    .D(next_first_round_reg),
    .RESET_B(net392),
    .Q(first_round_reg));
 sky130_fd_sc_hd__dfrtp_4 _7857_ (.CLK(clknet_leaf_32_clk),
    .D(_0144_),
    .RESET_B(net470),
    .Q(\sub1.data_o[72] ));
 sky130_fd_sc_hd__dfrtp_4 _7858_ (.CLK(clknet_leaf_36_clk),
    .D(_0145_),
    .RESET_B(net475),
    .Q(\sub1.data_o[73] ));
 sky130_fd_sc_hd__dfrtp_4 _7859_ (.CLK(clknet_leaf_32_clk),
    .D(_0146_),
    .RESET_B(net470),
    .Q(\sub1.data_o[74] ));
 sky130_fd_sc_hd__dfrtp_4 _7860_ (.CLK(clknet_leaf_32_clk),
    .D(_0147_),
    .RESET_B(net470),
    .Q(\sub1.data_o[75] ));
 sky130_fd_sc_hd__dfrtp_4 _7861_ (.CLK(clknet_leaf_32_clk),
    .D(_0148_),
    .RESET_B(net471),
    .Q(\sub1.data_o[76] ));
 sky130_fd_sc_hd__dfrtp_4 _7862_ (.CLK(clknet_leaf_38_clk),
    .D(_0149_),
    .RESET_B(net475),
    .Q(\sub1.data_o[77] ));
 sky130_fd_sc_hd__dfrtp_4 _7863_ (.CLK(clknet_leaf_31_clk),
    .D(_0150_),
    .RESET_B(net470),
    .Q(\sub1.data_o[78] ));
 sky130_fd_sc_hd__dfrtp_4 _7864_ (.CLK(clknet_leaf_32_clk),
    .D(_0151_),
    .RESET_B(net470),
    .Q(\sub1.data_o[79] ));
 sky130_fd_sc_hd__dfrtp_4 _7865_ (.CLK(clknet_leaf_72_clk),
    .D(\sbox1.intermediate_to_invert_var[0] ),
    .RESET_B(net413),
    .Q(\sbox1.inversion_to_invert_var[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7866_ (.CLK(clknet_leaf_71_clk),
    .D(\sbox1.intermediate_to_invert_var[1] ),
    .RESET_B(net412),
    .Q(\sbox1.inversion_to_invert_var[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7867_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sbox1.intermediate_to_invert_var[2] ),
    .RESET_B(net394),
    .Q(\sbox1.inversion_to_invert_var[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7868_ (.CLK(clknet_leaf_71_clk),
    .D(\sbox1.intermediate_to_invert_var[3] ),
    .RESET_B(net412),
    .Q(\sbox1.inversion_to_invert_var[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7869_ (.CLK(clknet_leaf_72_clk),
    .D(\sbox1.next_alph[0] ),
    .RESET_B(net413),
    .Q(\sbox1.alph[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7870_ (.CLK(clknet_leaf_71_clk),
    .D(\sbox1.next_alph[1] ),
    .RESET_B(net412),
    .Q(\sbox1.alph[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7871_ (.CLK(clknet_leaf_72_clk),
    .D(\sbox1.next_alph[2] ),
    .RESET_B(net413),
    .Q(\sbox1.alph[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7872_ (.CLK(clknet_leaf_71_clk),
    .D(\sbox1.next_alph[3] ),
    .RESET_B(net413),
    .Q(\sbox1.alph[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7873_ (.CLK(clknet_leaf_71_clk),
    .D(\sbox1.ah[0] ),
    .RESET_B(net412),
    .Q(\sbox1.ah_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7874_ (.CLK(clknet_leaf_71_clk),
    .D(\sbox1.ah[1] ),
    .RESET_B(net412),
    .Q(\sbox1.ah_reg[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7875_ (.CLK(clknet_leaf_71_clk),
    .D(\sbox1.ah[2] ),
    .RESET_B(net412),
    .Q(\sbox1.ah_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7876_ (.CLK(clknet_leaf_71_clk),
    .D(\sbox1.ah[3] ),
    .RESET_B(net412),
    .Q(\sbox1.ah_reg[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7877_ (.CLK(clknet_leaf_37_clk),
    .D(_0152_),
    .RESET_B(net476),
    .Q(\ks1.col[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7878_ (.CLK(clknet_leaf_37_clk),
    .D(_0153_),
    .RESET_B(net476),
    .Q(\ks1.col[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7879_ (.CLK(clknet_leaf_36_clk),
    .D(_0154_),
    .RESET_B(net476),
    .Q(\ks1.col[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7880_ (.CLK(clknet_leaf_37_clk),
    .D(_0155_),
    .RESET_B(net480),
    .Q(\ks1.col[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7881_ (.CLK(clknet_leaf_68_clk),
    .D(_0156_),
    .RESET_B(net420),
    .Q(\ks1.col[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7882_ (.CLK(clknet_leaf_68_clk),
    .D(_0157_),
    .RESET_B(net420),
    .Q(\ks1.col[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7883_ (.CLK(clknet_leaf_38_clk),
    .D(_0158_),
    .RESET_B(net475),
    .Q(\ks1.col[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7884_ (.CLK(clknet_leaf_40_clk),
    .D(_0159_),
    .RESET_B(net480),
    .Q(\ks1.col[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7885_ (.CLK(clknet_leaf_70_clk),
    .D(_0160_),
    .RESET_B(net417),
    .Q(\ks1.col[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7886_ (.CLK(clknet_leaf_70_clk),
    .D(_0161_),
    .RESET_B(net415),
    .Q(\ks1.col[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7887_ (.CLK(clknet_leaf_68_clk),
    .D(_0162_),
    .RESET_B(net420),
    .Q(\ks1.col[26] ));
 sky130_fd_sc_hd__dfrtp_2 _7888_ (.CLK(clknet_leaf_68_clk),
    .D(_0163_),
    .RESET_B(net415),
    .Q(\ks1.col[27] ));
 sky130_fd_sc_hd__dfrtp_2 _7889_ (.CLK(clknet_leaf_74_clk),
    .D(_0164_),
    .RESET_B(net414),
    .Q(\ks1.col[28] ));
 sky130_fd_sc_hd__dfrtp_1 _7890_ (.CLK(clknet_leaf_74_clk),
    .D(_0165_),
    .RESET_B(net415),
    .Q(\ks1.col[29] ));
 sky130_fd_sc_hd__dfrtp_1 _7891_ (.CLK(clknet_leaf_70_clk),
    .D(_0166_),
    .RESET_B(net417),
    .Q(\ks1.col[30] ));
 sky130_fd_sc_hd__dfrtp_4 _7892_ (.CLK(clknet_leaf_70_clk),
    .D(_0167_),
    .RESET_B(net413),
    .Q(\ks1.col[31] ));
 sky130_fd_sc_hd__dfrtp_4 _7893_ (.CLK(clknet_leaf_74_clk),
    .D(_0168_),
    .RESET_B(net415),
    .Q(\ks1.col[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7894_ (.CLK(clknet_leaf_40_clk),
    .D(_0169_),
    .RESET_B(net478),
    .Q(\ks1.col[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7895_ (.CLK(clknet_leaf_38_clk),
    .D(_0170_),
    .RESET_B(net475),
    .Q(\ks1.col[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7896_ (.CLK(clknet_leaf_40_clk),
    .D(_0171_),
    .RESET_B(net480),
    .Q(\ks1.col[19] ));
 sky130_fd_sc_hd__dfrtp_4 _7897_ (.CLK(clknet_leaf_75_clk),
    .D(_0172_),
    .RESET_B(net421),
    .Q(\ks1.col[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7898_ (.CLK(clknet_leaf_44_clk),
    .D(_0173_),
    .RESET_B(net477),
    .Q(\ks1.col[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7899_ (.CLK(clknet_leaf_39_clk),
    .D(_0174_),
    .RESET_B(net471),
    .Q(\ks1.col[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7900_ (.CLK(clknet_leaf_40_clk),
    .D(_0175_),
    .RESET_B(net478),
    .Q(\ks1.col[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7901_ (.CLK(clknet_leaf_1_clk),
    .D(_0176_),
    .RESET_B(net395),
    .Q(\mix1.data_reg[64] ));
 sky130_fd_sc_hd__dfrtp_1 _7902_ (.CLK(clknet_leaf_1_clk),
    .D(_0177_),
    .RESET_B(net395),
    .Q(\mix1.data_reg[65] ));
 sky130_fd_sc_hd__dfrtp_1 _7903_ (.CLK(clknet_leaf_2_clk),
    .D(_0178_),
    .RESET_B(net402),
    .Q(\mix1.data_reg[66] ));
 sky130_fd_sc_hd__dfrtp_1 _7904_ (.CLK(clknet_leaf_2_clk),
    .D(_0179_),
    .RESET_B(net434),
    .Q(\mix1.data_reg[67] ));
 sky130_fd_sc_hd__dfrtp_1 _7905_ (.CLK(clknet_leaf_2_clk),
    .D(_0180_),
    .RESET_B(net401),
    .Q(\mix1.data_reg[68] ));
 sky130_fd_sc_hd__dfrtp_1 _7906_ (.CLK(clknet_leaf_2_clk),
    .D(_0181_),
    .RESET_B(net402),
    .Q(\mix1.data_reg[69] ));
 sky130_fd_sc_hd__dfrtp_1 _7907_ (.CLK(clknet_leaf_12_clk),
    .D(_0182_),
    .RESET_B(net434),
    .Q(\mix1.data_reg[70] ));
 sky130_fd_sc_hd__dfrtp_1 _7908_ (.CLK(clknet_leaf_2_clk),
    .D(_0183_),
    .RESET_B(net402),
    .Q(\mix1.data_reg[71] ));
 sky130_fd_sc_hd__dfrtp_1 _7909_ (.CLK(clknet_leaf_2_clk),
    .D(_0184_),
    .RESET_B(net402),
    .Q(\mix1.data_reg[72] ));
 sky130_fd_sc_hd__dfrtp_1 _7910_ (.CLK(clknet_leaf_3_clk),
    .D(_0185_),
    .RESET_B(net401),
    .Q(\mix1.data_reg[73] ));
 sky130_fd_sc_hd__dfrtp_1 _7911_ (.CLK(clknet_leaf_2_clk),
    .D(_0186_),
    .RESET_B(net402),
    .Q(\mix1.data_reg[74] ));
 sky130_fd_sc_hd__dfrtp_1 _7912_ (.CLK(clknet_leaf_3_clk),
    .D(_0187_),
    .RESET_B(net402),
    .Q(\mix1.data_reg[75] ));
 sky130_fd_sc_hd__dfrtp_1 _7913_ (.CLK(clknet_leaf_1_clk),
    .D(_0188_),
    .RESET_B(net395),
    .Q(\mix1.data_reg[76] ));
 sky130_fd_sc_hd__dfrtp_1 _7914_ (.CLK(clknet_leaf_3_clk),
    .D(_0189_),
    .RESET_B(net406),
    .Q(\mix1.data_reg[77] ));
 sky130_fd_sc_hd__dfrtp_1 _7915_ (.CLK(clknet_leaf_1_clk),
    .D(_0190_),
    .RESET_B(net401),
    .Q(\mix1.data_reg[78] ));
 sky130_fd_sc_hd__dfrtp_1 _7916_ (.CLK(clknet_leaf_6_clk),
    .D(_0191_),
    .RESET_B(net398),
    .Q(\mix1.data_reg[79] ));
 sky130_fd_sc_hd__dfrtp_1 _7917_ (.CLK(clknet_leaf_18_clk),
    .D(_0192_),
    .RESET_B(net444),
    .Q(\mix1.data_reg[80] ));
 sky130_fd_sc_hd__dfrtp_1 _7918_ (.CLK(clknet_leaf_17_clk),
    .D(_0193_),
    .RESET_B(net445),
    .Q(\mix1.data_reg[81] ));
 sky130_fd_sc_hd__dfrtp_1 _7919_ (.CLK(clknet_leaf_17_clk),
    .D(_0194_),
    .RESET_B(net445),
    .Q(\mix1.data_reg[82] ));
 sky130_fd_sc_hd__dfrtp_1 _7920_ (.CLK(clknet_leaf_20_clk),
    .D(_0195_),
    .RESET_B(net447),
    .Q(\mix1.data_reg[83] ));
 sky130_fd_sc_hd__dfrtp_1 _7921_ (.CLK(clknet_leaf_19_clk),
    .D(_0196_),
    .RESET_B(net447),
    .Q(\mix1.data_reg[84] ));
 sky130_fd_sc_hd__dfrtp_1 _7922_ (.CLK(clknet_leaf_17_clk),
    .D(_0197_),
    .RESET_B(net447),
    .Q(\mix1.data_reg[85] ));
 sky130_fd_sc_hd__dfrtp_1 _7923_ (.CLK(clknet_leaf_19_clk),
    .D(_0198_),
    .RESET_B(net447),
    .Q(\mix1.data_reg[86] ));
 sky130_fd_sc_hd__dfrtp_1 _7924_ (.CLK(clknet_leaf_17_clk),
    .D(_0199_),
    .RESET_B(net446),
    .Q(\mix1.data_reg[87] ));
 sky130_fd_sc_hd__dfrtp_1 _7925_ (.CLK(clknet_leaf_6_clk),
    .D(_0200_),
    .RESET_B(net397),
    .Q(\mix1.data_reg[88] ));
 sky130_fd_sc_hd__dfrtp_1 _7926_ (.CLK(clknet_leaf_87_clk),
    .D(_0201_),
    .RESET_B(net394),
    .Q(\mix1.data_reg[89] ));
 sky130_fd_sc_hd__dfrtp_1 _7927_ (.CLK(clknet_leaf_87_clk),
    .D(_0202_),
    .RESET_B(net390),
    .Q(\mix1.data_reg[90] ));
 sky130_fd_sc_hd__dfrtp_1 _7928_ (.CLK(clknet_leaf_87_clk),
    .D(_0203_),
    .RESET_B(net394),
    .Q(\mix1.data_reg[91] ));
 sky130_fd_sc_hd__dfrtp_1 _7929_ (.CLK(clknet_leaf_87_clk),
    .D(_0204_),
    .RESET_B(net394),
    .Q(\mix1.data_reg[92] ));
 sky130_fd_sc_hd__dfrtp_1 _7930_ (.CLK(clknet_leaf_0_clk),
    .D(_0205_),
    .RESET_B(net397),
    .Q(\mix1.data_reg[93] ));
 sky130_fd_sc_hd__dfrtp_1 _7931_ (.CLK(clknet_leaf_0_clk),
    .D(_0206_),
    .RESET_B(net396),
    .Q(\mix1.data_reg[94] ));
 sky130_fd_sc_hd__dfrtp_1 _7932_ (.CLK(clknet_leaf_0_clk),
    .D(_0207_),
    .RESET_B(net396),
    .Q(\mix1.data_reg[95] ));
 sky130_fd_sc_hd__dfrtp_1 _7933_ (.CLK(clknet_leaf_1_clk),
    .D(_0208_),
    .RESET_B(net395),
    .Q(\mix1.data_reg[32] ));
 sky130_fd_sc_hd__dfrtp_1 _7934_ (.CLK(clknet_leaf_1_clk),
    .D(_0209_),
    .RESET_B(net395),
    .Q(\mix1.data_reg[33] ));
 sky130_fd_sc_hd__dfrtp_1 _7935_ (.CLK(clknet_leaf_12_clk),
    .D(_0210_),
    .RESET_B(net434),
    .Q(\mix1.data_reg[34] ));
 sky130_fd_sc_hd__dfrtp_1 _7936_ (.CLK(clknet_leaf_14_clk),
    .D(_0211_),
    .RESET_B(net440),
    .Q(\mix1.data_reg[35] ));
 sky130_fd_sc_hd__dfrtp_1 _7937_ (.CLK(clknet_leaf_14_clk),
    .D(_0212_),
    .RESET_B(net439),
    .Q(\mix1.data_reg[36] ));
 sky130_fd_sc_hd__dfrtp_1 _7938_ (.CLK(clknet_leaf_14_clk),
    .D(_0213_),
    .RESET_B(net439),
    .Q(\mix1.data_reg[37] ));
 sky130_fd_sc_hd__dfrtp_1 _7939_ (.CLK(clknet_leaf_15_clk),
    .D(_0214_),
    .RESET_B(net440),
    .Q(\mix1.data_reg[38] ));
 sky130_fd_sc_hd__dfrtp_1 _7940_ (.CLK(clknet_leaf_14_clk),
    .D(_0215_),
    .RESET_B(net439),
    .Q(\mix1.data_reg[39] ));
 sky130_fd_sc_hd__dfrtp_1 _7941_ (.CLK(clknet_leaf_13_clk),
    .D(_0216_),
    .RESET_B(net434),
    .Q(\mix1.data_reg[40] ));
 sky130_fd_sc_hd__dfrtp_1 _7942_ (.CLK(clknet_leaf_12_clk),
    .D(_0217_),
    .RESET_B(net434),
    .Q(\mix1.data_reg[41] ));
 sky130_fd_sc_hd__dfrtp_1 _7943_ (.CLK(clknet_leaf_13_clk),
    .D(_0218_),
    .RESET_B(net436),
    .Q(\mix1.data_reg[42] ));
 sky130_fd_sc_hd__dfrtp_1 _7944_ (.CLK(clknet_leaf_12_clk),
    .D(_0219_),
    .RESET_B(net434),
    .Q(\mix1.data_reg[43] ));
 sky130_fd_sc_hd__dfrtp_1 _7945_ (.CLK(clknet_leaf_12_clk),
    .D(_0220_),
    .RESET_B(net434),
    .Q(\mix1.data_reg[44] ));
 sky130_fd_sc_hd__dfrtp_1 _7946_ (.CLK(clknet_leaf_12_clk),
    .D(_0221_),
    .RESET_B(net436),
    .Q(\mix1.data_reg[45] ));
 sky130_fd_sc_hd__dfrtp_1 _7947_ (.CLK(clknet_leaf_12_clk),
    .D(_0222_),
    .RESET_B(net435),
    .Q(\mix1.data_reg[46] ));
 sky130_fd_sc_hd__dfrtp_1 _7948_ (.CLK(clknet_leaf_13_clk),
    .D(_0223_),
    .RESET_B(net436),
    .Q(\mix1.data_reg[47] ));
 sky130_fd_sc_hd__dfrtp_1 _7949_ (.CLK(clknet_leaf_14_clk),
    .D(_0224_),
    .RESET_B(net439),
    .Q(\mix1.data_reg[48] ));
 sky130_fd_sc_hd__dfrtp_1 _7950_ (.CLK(clknet_leaf_17_clk),
    .D(_0225_),
    .RESET_B(net444),
    .Q(\mix1.data_reg[49] ));
 sky130_fd_sc_hd__dfrtp_1 _7951_ (.CLK(clknet_leaf_15_clk),
    .D(_0226_),
    .RESET_B(net440),
    .Q(\mix1.data_reg[50] ));
 sky130_fd_sc_hd__dfrtp_1 _7952_ (.CLK(clknet_leaf_16_clk),
    .D(_0227_),
    .RESET_B(net446),
    .Q(\mix1.data_reg[51] ));
 sky130_fd_sc_hd__dfrtp_1 _7953_ (.CLK(clknet_leaf_20_clk),
    .D(_0228_),
    .RESET_B(net446),
    .Q(\mix1.data_reg[52] ));
 sky130_fd_sc_hd__dfrtp_1 _7954_ (.CLK(clknet_leaf_16_clk),
    .D(_0229_),
    .RESET_B(net446),
    .Q(\mix1.data_reg[53] ));
 sky130_fd_sc_hd__dfrtp_1 _7955_ (.CLK(clknet_leaf_16_clk),
    .D(_0230_),
    .RESET_B(net446),
    .Q(\mix1.data_reg[54] ));
 sky130_fd_sc_hd__dfrtp_1 _7956_ (.CLK(clknet_leaf_17_clk),
    .D(_0231_),
    .RESET_B(net444),
    .Q(\mix1.data_reg[55] ));
 sky130_fd_sc_hd__dfrtp_1 _7957_ (.CLK(clknet_leaf_6_clk),
    .D(_0232_),
    .RESET_B(net398),
    .Q(\mix1.data_reg[56] ));
 sky130_fd_sc_hd__dfrtp_1 _7958_ (.CLK(clknet_leaf_5_clk),
    .D(_0233_),
    .RESET_B(net404),
    .Q(\mix1.data_reg[57] ));
 sky130_fd_sc_hd__dfrtp_1 _7959_ (.CLK(clknet_leaf_6_clk),
    .D(_0234_),
    .RESET_B(net398),
    .Q(\mix1.data_reg[58] ));
 sky130_fd_sc_hd__dfrtp_1 _7960_ (.CLK(clknet_leaf_6_clk),
    .D(_0235_),
    .RESET_B(net398),
    .Q(\mix1.data_reg[59] ));
 sky130_fd_sc_hd__dfrtp_1 _7961_ (.CLK(clknet_leaf_6_clk),
    .D(_0236_),
    .RESET_B(net399),
    .Q(\mix1.data_reg[60] ));
 sky130_fd_sc_hd__dfrtp_1 _7962_ (.CLK(clknet_leaf_0_clk),
    .D(_0237_),
    .RESET_B(net398),
    .Q(\mix1.data_reg[61] ));
 sky130_fd_sc_hd__dfrtp_1 _7963_ (.CLK(clknet_leaf_1_clk),
    .D(_0238_),
    .RESET_B(net395),
    .Q(\mix1.data_reg[62] ));
 sky130_fd_sc_hd__dfrtp_1 _7964_ (.CLK(clknet_leaf_0_clk),
    .D(_0239_),
    .RESET_B(net398),
    .Q(\mix1.data_reg[63] ));
 sky130_fd_sc_hd__dfrtp_2 _7965_ (.CLK(clknet_leaf_81_clk),
    .D(_0240_),
    .RESET_B(net390),
    .Q(\sub1.data_o[120] ));
 sky130_fd_sc_hd__dfrtp_2 _7966_ (.CLK(clknet_leaf_73_clk),
    .D(_0241_),
    .RESET_B(net414),
    .Q(\sub1.data_o[121] ));
 sky130_fd_sc_hd__dfrtp_1 _7967_ (.CLK(clknet_leaf_81_clk),
    .D(_0242_),
    .RESET_B(net390),
    .Q(\sub1.data_o[122] ));
 sky130_fd_sc_hd__dfrtp_2 _7968_ (.CLK(clknet_leaf_79_clk),
    .D(_0243_),
    .RESET_B(net392),
    .Q(\sub1.data_o[123] ));
 sky130_fd_sc_hd__dfrtp_2 _7969_ (.CLK(clknet_leaf_81_clk),
    .D(_0244_),
    .RESET_B(net393),
    .Q(\sub1.data_o[124] ));
 sky130_fd_sc_hd__dfrtp_4 _7970_ (.CLK(clknet_leaf_77_clk),
    .D(_0245_),
    .RESET_B(net422),
    .Q(\sub1.data_o[125] ));
 sky130_fd_sc_hd__dfrtp_4 _7971_ (.CLK(clknet_leaf_83_clk),
    .D(_0246_),
    .RESET_B(net392),
    .Q(\sub1.data_o[126] ));
 sky130_fd_sc_hd__dfrtp_2 _7972_ (.CLK(clknet_leaf_81_clk),
    .D(_0247_),
    .RESET_B(net393),
    .Q(\sub1.data_o[127] ));
 sky130_fd_sc_hd__dfrtp_1 _7973_ (.CLK(clknet_leaf_26_clk),
    .D(_0248_),
    .RESET_B(net443),
    .Q(\sub1.data_o[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7974_ (.CLK(clknet_leaf_10_clk),
    .D(_0249_),
    .RESET_B(net443),
    .Q(\sub1.data_o[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7975_ (.CLK(clknet_leaf_10_clk),
    .D(_0250_),
    .RESET_B(net443),
    .Q(\sub1.data_o[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7976_ (.CLK(clknet_leaf_26_clk),
    .D(_0251_),
    .RESET_B(net443),
    .Q(\sub1.data_o[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7977_ (.CLK(clknet_leaf_20_clk),
    .D(_0252_),
    .RESET_B(net450),
    .Q(\sub1.data_o[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7978_ (.CLK(clknet_leaf_26_clk),
    .D(_0253_),
    .RESET_B(net443),
    .Q(\sub1.data_o[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7979_ (.CLK(clknet_leaf_26_clk),
    .D(_0254_),
    .RESET_B(net455),
    .Q(\sub1.data_o[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7980_ (.CLK(clknet_leaf_20_clk),
    .D(_0255_),
    .RESET_B(net450),
    .Q(\sub1.data_o[7] ));
 sky130_fd_sc_hd__dfrtp_4 _7981_ (.CLK(clknet_leaf_32_clk),
    .D(_0256_),
    .RESET_B(net471),
    .Q(\sub1.data_o[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7982_ (.CLK(clknet_leaf_38_clk),
    .D(_0257_),
    .RESET_B(net471),
    .Q(\sub1.data_o[9] ));
 sky130_fd_sc_hd__dfrtp_4 _7983_ (.CLK(clknet_leaf_38_clk),
    .D(_0258_),
    .RESET_B(net471),
    .Q(\sub1.data_o[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7984_ (.CLK(clknet_leaf_31_clk),
    .D(_0259_),
    .RESET_B(net470),
    .Q(\sub1.data_o[11] ));
 sky130_fd_sc_hd__dfrtp_4 _7985_ (.CLK(clknet_leaf_32_clk),
    .D(_0260_),
    .RESET_B(net469),
    .Q(\sub1.data_o[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7986_ (.CLK(clknet_leaf_38_clk),
    .D(_0261_),
    .RESET_B(net475),
    .Q(\sub1.data_o[13] ));
 sky130_fd_sc_hd__dfrtp_4 _7987_ (.CLK(clknet_leaf_39_clk),
    .D(_0262_),
    .RESET_B(net470),
    .Q(\sub1.data_o[14] ));
 sky130_fd_sc_hd__dfrtp_2 _7988_ (.CLK(clknet_leaf_39_clk),
    .D(_0263_),
    .RESET_B(net470),
    .Q(\sub1.data_o[15] ));
 sky130_fd_sc_hd__dfrtp_4 _7989_ (.CLK(clknet_leaf_36_clk),
    .D(_0264_),
    .RESET_B(net476),
    .Q(\sub1.data_o[16] ));
 sky130_fd_sc_hd__dfrtp_4 _7990_ (.CLK(clknet_leaf_36_clk),
    .D(_0265_),
    .RESET_B(net473),
    .Q(\sub1.data_o[17] ));
 sky130_fd_sc_hd__dfrtp_4 _7991_ (.CLK(clknet_leaf_36_clk),
    .D(_0266_),
    .RESET_B(net473),
    .Q(\sub1.data_o[18] ));
 sky130_fd_sc_hd__dfrtp_4 _7992_ (.CLK(clknet_leaf_36_clk),
    .D(_0267_),
    .RESET_B(net476),
    .Q(\sub1.data_o[19] ));
 sky130_fd_sc_hd__dfrtp_4 _7993_ (.CLK(clknet_leaf_36_clk),
    .D(_0268_),
    .RESET_B(net475),
    .Q(\sub1.data_o[20] ));
 sky130_fd_sc_hd__dfrtp_4 _7994_ (.CLK(clknet_leaf_36_clk),
    .D(_0269_),
    .RESET_B(net476),
    .Q(\sub1.data_o[21] ));
 sky130_fd_sc_hd__dfrtp_4 _7995_ (.CLK(clknet_leaf_36_clk),
    .D(_0270_),
    .RESET_B(net475),
    .Q(\sub1.data_o[22] ));
 sky130_fd_sc_hd__dfrtp_4 _7996_ (.CLK(clknet_leaf_36_clk),
    .D(_0271_),
    .RESET_B(net475),
    .Q(\sub1.data_o[23] ));
 sky130_fd_sc_hd__dfrtp_2 _7997_ (.CLK(clknet_leaf_57_clk),
    .D(_0272_),
    .RESET_B(net458),
    .Q(\sub1.data_o[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7998_ (.CLK(clknet_leaf_57_clk),
    .D(_0273_),
    .RESET_B(net423),
    .Q(\sub1.data_o[25] ));
 sky130_fd_sc_hd__dfrtp_2 _7999_ (.CLK(clknet_leaf_56_clk),
    .D(_0274_),
    .RESET_B(net423),
    .Q(\sub1.data_o[26] ));
 sky130_fd_sc_hd__dfrtp_2 _8000_ (.CLK(clknet_leaf_53_clk),
    .D(_0275_),
    .RESET_B(net458),
    .Q(\sub1.data_o[27] ));
 sky130_fd_sc_hd__dfrtp_2 _8001_ (.CLK(clknet_leaf_57_clk),
    .D(_0276_),
    .RESET_B(net423),
    .Q(\sub1.data_o[28] ));
 sky130_fd_sc_hd__dfrtp_2 _8002_ (.CLK(clknet_leaf_53_clk),
    .D(_0277_),
    .RESET_B(net458),
    .Q(\sub1.data_o[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8003_ (.CLK(clknet_leaf_57_clk),
    .D(_0278_),
    .RESET_B(net423),
    .Q(\sub1.data_o[30] ));
 sky130_fd_sc_hd__dfrtp_2 _8004_ (.CLK(clknet_leaf_56_clk),
    .D(_0279_),
    .RESET_B(net433),
    .Q(\sub1.data_o[31] ));
 sky130_fd_sc_hd__dfrtp_4 _8005_ (.CLK(clknet_leaf_20_clk),
    .D(_0280_),
    .RESET_B(net450),
    .Q(\sub1.data_o[32] ));
 sky130_fd_sc_hd__dfrtp_4 _8006_ (.CLK(clknet_leaf_25_clk),
    .D(_0281_),
    .RESET_B(net454),
    .Q(\sub1.data_o[33] ));
 sky130_fd_sc_hd__dfrtp_4 _8007_ (.CLK(clknet_leaf_20_clk),
    .D(_0282_),
    .RESET_B(net450),
    .Q(\sub1.data_o[34] ));
 sky130_fd_sc_hd__dfrtp_4 _8008_ (.CLK(clknet_leaf_20_clk),
    .D(_0283_),
    .RESET_B(net450),
    .Q(\sub1.data_o[35] ));
 sky130_fd_sc_hd__dfrtp_4 _8009_ (.CLK(clknet_leaf_20_clk),
    .D(_0284_),
    .RESET_B(net450),
    .Q(\sub1.data_o[36] ));
 sky130_fd_sc_hd__dfrtp_4 _8010_ (.CLK(clknet_leaf_25_clk),
    .D(_0285_),
    .RESET_B(net450),
    .Q(\sub1.data_o[37] ));
 sky130_fd_sc_hd__dfrtp_4 _8011_ (.CLK(clknet_leaf_25_clk),
    .D(_0286_),
    .RESET_B(net450),
    .Q(\sub1.data_o[38] ));
 sky130_fd_sc_hd__dfrtp_4 _8012_ (.CLK(clknet_leaf_20_clk),
    .D(_0287_),
    .RESET_B(net451),
    .Q(\sub1.data_o[39] ));
 sky130_fd_sc_hd__dfrtp_4 _8013_ (.CLK(clknet_leaf_30_clk),
    .D(_0288_),
    .RESET_B(net456),
    .Q(\sub1.data_o[40] ));
 sky130_fd_sc_hd__dfrtp_2 _8014_ (.CLK(clknet_leaf_30_clk),
    .D(_0289_),
    .RESET_B(net456),
    .Q(\sub1.data_o[41] ));
 sky130_fd_sc_hd__dfrtp_4 _8015_ (.CLK(clknet_leaf_30_clk),
    .D(_0290_),
    .RESET_B(net456),
    .Q(\sub1.data_o[42] ));
 sky130_fd_sc_hd__dfrtp_2 _8016_ (.CLK(clknet_leaf_30_clk),
    .D(_0291_),
    .RESET_B(net456),
    .Q(\sub1.data_o[43] ));
 sky130_fd_sc_hd__dfrtp_4 _8017_ (.CLK(clknet_leaf_30_clk),
    .D(_0292_),
    .RESET_B(net456),
    .Q(\sub1.data_o[44] ));
 sky130_fd_sc_hd__dfrtp_2 _8018_ (.CLK(clknet_leaf_30_clk),
    .D(_0293_),
    .RESET_B(net456),
    .Q(\sub1.data_o[45] ));
 sky130_fd_sc_hd__dfrtp_4 _8019_ (.CLK(clknet_leaf_30_clk),
    .D(_0294_),
    .RESET_B(net468),
    .Q(\sub1.data_o[46] ));
 sky130_fd_sc_hd__dfrtp_4 _8020_ (.CLK(clknet_leaf_30_clk),
    .D(_0295_),
    .RESET_B(net468),
    .Q(\sub1.data_o[47] ));
 sky130_fd_sc_hd__dfrtp_4 _8021_ (.CLK(clknet_leaf_23_clk),
    .D(_0296_),
    .RESET_B(net453),
    .Q(\sub1.data_o[48] ));
 sky130_fd_sc_hd__dfrtp_4 _8022_ (.CLK(clknet_leaf_35_clk),
    .D(_0297_),
    .RESET_B(net473),
    .Q(\sub1.data_o[49] ));
 sky130_fd_sc_hd__dfrtp_4 _8023_ (.CLK(clknet_leaf_35_clk),
    .D(_0298_),
    .RESET_B(net473),
    .Q(\sub1.data_o[50] ));
 sky130_fd_sc_hd__dfrtp_4 _8024_ (.CLK(clknet_leaf_23_clk),
    .D(_0299_),
    .RESET_B(net453),
    .Q(\sub1.data_o[51] ));
 sky130_fd_sc_hd__dfrtp_4 _8025_ (.CLK(clknet_leaf_34_clk),
    .D(_0300_),
    .RESET_B(net474),
    .Q(\sub1.data_o[52] ));
 sky130_fd_sc_hd__dfrtp_4 _8026_ (.CLK(clknet_leaf_36_clk),
    .D(_0301_),
    .RESET_B(net474),
    .Q(\sub1.data_o[53] ));
 sky130_fd_sc_hd__dfrtp_4 _8027_ (.CLK(clknet_leaf_24_clk),
    .D(_0302_),
    .RESET_B(net452),
    .Q(\sub1.data_o[54] ));
 sky130_fd_sc_hd__dfrtp_4 _8028_ (.CLK(clknet_leaf_34_clk),
    .D(_0303_),
    .RESET_B(net474),
    .Q(\sub1.data_o[55] ));
 sky130_fd_sc_hd__dfrtp_1 _8029_ (.CLK(clknet_leaf_78_clk),
    .D(_0304_),
    .RESET_B(net423),
    .Q(\sub1.data_o[56] ));
 sky130_fd_sc_hd__dfrtp_1 _8030_ (.CLK(clknet_leaf_78_clk),
    .D(_0305_),
    .RESET_B(net422),
    .Q(\sub1.data_o[57] ));
 sky130_fd_sc_hd__dfrtp_1 _8031_ (.CLK(clknet_leaf_79_clk),
    .D(_0306_),
    .RESET_B(net409),
    .Q(\sub1.data_o[58] ));
 sky130_fd_sc_hd__dfrtp_1 _8032_ (.CLK(clknet_leaf_78_clk),
    .D(_0307_),
    .RESET_B(net423),
    .Q(\sub1.data_o[59] ));
 sky130_fd_sc_hd__dfrtp_2 _8033_ (.CLK(clknet_leaf_76_clk),
    .D(_0308_),
    .RESET_B(net421),
    .Q(\sub1.data_o[60] ));
 sky130_fd_sc_hd__dfrtp_2 _8034_ (.CLK(clknet_leaf_76_clk),
    .D(_0309_),
    .RESET_B(net422),
    .Q(\sub1.data_o[61] ));
 sky130_fd_sc_hd__dfrtp_1 _8035_ (.CLK(clknet_leaf_76_clk),
    .D(_0310_),
    .RESET_B(net422),
    .Q(\sub1.data_o[62] ));
 sky130_fd_sc_hd__dfrtp_2 _8036_ (.CLK(clknet_leaf_80_clk),
    .D(_0311_),
    .RESET_B(net409),
    .Q(\sub1.data_o[63] ));
 sky130_fd_sc_hd__dfrtp_4 _8037_ (.CLK(clknet_leaf_34_clk),
    .D(_0312_),
    .RESET_B(net469),
    .Q(\sub1.data_o[64] ));
 sky130_fd_sc_hd__dfrtp_4 _8038_ (.CLK(clknet_leaf_34_clk),
    .D(_0313_),
    .RESET_B(net469),
    .Q(\sub1.data_o[65] ));
 sky130_fd_sc_hd__dfrtp_4 _8039_ (.CLK(clknet_leaf_33_clk),
    .D(_0314_),
    .RESET_B(net472),
    .Q(\sub1.data_o[66] ));
 sky130_fd_sc_hd__dfrtp_4 _8040_ (.CLK(clknet_leaf_33_clk),
    .D(_0315_),
    .RESET_B(net469),
    .Q(\sub1.data_o[67] ));
 sky130_fd_sc_hd__dfrtp_4 _8041_ (.CLK(clknet_leaf_32_clk),
    .D(_0316_),
    .RESET_B(net469),
    .Q(\sub1.data_o[68] ));
 sky130_fd_sc_hd__dfrtp_4 _8042_ (.CLK(clknet_leaf_33_clk),
    .D(_0317_),
    .RESET_B(net469),
    .Q(\sub1.data_o[69] ));
 sky130_fd_sc_hd__dfrtp_4 _8043_ (.CLK(clknet_leaf_33_clk),
    .D(_0318_),
    .RESET_B(net469),
    .Q(\sub1.data_o[70] ));
 sky130_fd_sc_hd__dfrtp_4 _8044_ (.CLK(clknet_leaf_32_clk),
    .D(_0319_),
    .RESET_B(net472),
    .Q(\sub1.data_o[71] ));
 sky130_fd_sc_hd__dfrtp_2 _8045_ (.CLK(clknet_leaf_77_clk),
    .D(\sub1.next_ready_o ),
    .RESET_B(net422),
    .Q(\sub1.ready_o ));
 sky130_fd_sc_hd__dfrtp_2 _8046_ (.CLK(clknet_leaf_5_clk),
    .D(_0320_),
    .RESET_B(net404),
    .Q(\mix1.data_o[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8047_ (.CLK(clknet_leaf_9_clk),
    .D(_0321_),
    .RESET_B(net443),
    .Q(\mix1.data_o[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8048_ (.CLK(clknet_leaf_8_clk),
    .D(_0322_),
    .RESET_B(net410),
    .Q(\mix1.data_o[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8049_ (.CLK(clknet_leaf_4_clk),
    .D(_0323_),
    .RESET_B(net406),
    .Q(\mix1.data_o[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8050_ (.CLK(clknet_leaf_5_clk),
    .D(_0324_),
    .RESET_B(net404),
    .Q(\mix1.data_o[4] ));
 sky130_fd_sc_hd__dfrtp_4 _8051_ (.CLK(clknet_leaf_12_clk),
    .D(_0325_),
    .RESET_B(net438),
    .Q(\mix1.data_o[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8052_ (.CLK(clknet_leaf_4_clk),
    .D(_0326_),
    .RESET_B(net438),
    .Q(\mix1.data_o[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8053_ (.CLK(clknet_leaf_3_clk),
    .D(_0327_),
    .RESET_B(net404),
    .Q(\mix1.data_o[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8054_ (.CLK(clknet_leaf_8_clk),
    .D(_0328_),
    .RESET_B(net443),
    .Q(\mix1.data_o[8] ));
 sky130_fd_sc_hd__dfrtp_2 _8055_ (.CLK(clknet_leaf_4_clk),
    .D(_0329_),
    .RESET_B(net406),
    .Q(\mix1.data_o[9] ));
 sky130_fd_sc_hd__dfrtp_4 _8056_ (.CLK(clknet_leaf_13_clk),
    .D(_0330_),
    .RESET_B(net436),
    .Q(\mix1.data_o[10] ));
 sky130_fd_sc_hd__dfrtp_4 _8057_ (.CLK(clknet_leaf_4_clk),
    .D(_0331_),
    .RESET_B(net406),
    .Q(\mix1.data_o[11] ));
 sky130_fd_sc_hd__dfrtp_4 _8058_ (.CLK(clknet_leaf_11_clk),
    .D(_0332_),
    .RESET_B(net438),
    .Q(\mix1.data_o[12] ));
 sky130_fd_sc_hd__dfrtp_4 _8059_ (.CLK(clknet_leaf_13_clk),
    .D(_0333_),
    .RESET_B(net436),
    .Q(\mix1.data_o[13] ));
 sky130_fd_sc_hd__dfrtp_4 _8060_ (.CLK(clknet_leaf_12_clk),
    .D(_0334_),
    .RESET_B(net435),
    .Q(\mix1.data_o[14] ));
 sky130_fd_sc_hd__dfrtp_4 _8061_ (.CLK(clknet_leaf_13_clk),
    .D(_0335_),
    .RESET_B(net437),
    .Q(\mix1.data_o[15] ));
 sky130_fd_sc_hd__dfrtp_4 _8062_ (.CLK(clknet_leaf_16_clk),
    .D(_0336_),
    .RESET_B(net442),
    .Q(\mix1.data_o[16] ));
 sky130_fd_sc_hd__dfrtp_4 _8063_ (.CLK(clknet_leaf_16_clk),
    .D(_0337_),
    .RESET_B(net442),
    .Q(\mix1.data_o[17] ));
 sky130_fd_sc_hd__dfrtp_4 _8064_ (.CLK(clknet_leaf_10_clk),
    .D(_0338_),
    .RESET_B(net442),
    .Q(\mix1.data_o[18] ));
 sky130_fd_sc_hd__dfrtp_4 _8065_ (.CLK(clknet_leaf_16_clk),
    .D(_0339_),
    .RESET_B(net442),
    .Q(\mix1.data_o[19] ));
 sky130_fd_sc_hd__dfrtp_4 _8066_ (.CLK(clknet_leaf_16_clk),
    .D(_0340_),
    .RESET_B(net442),
    .Q(\mix1.data_o[20] ));
 sky130_fd_sc_hd__dfrtp_4 _8067_ (.CLK(clknet_leaf_16_clk),
    .D(_0341_),
    .RESET_B(net446),
    .Q(\mix1.data_o[21] ));
 sky130_fd_sc_hd__dfrtp_4 _8068_ (.CLK(clknet_leaf_16_clk),
    .D(_0342_),
    .RESET_B(net442),
    .Q(\mix1.data_o[22] ));
 sky130_fd_sc_hd__dfrtp_4 _8069_ (.CLK(clknet_leaf_16_clk),
    .D(_0343_),
    .RESET_B(net446),
    .Q(\mix1.data_o[23] ));
 sky130_fd_sc_hd__dfrtp_4 _8070_ (.CLK(clknet_leaf_4_clk),
    .D(_0344_),
    .RESET_B(net406),
    .Q(\mix1.data_o[24] ));
 sky130_fd_sc_hd__dfrtp_4 _8071_ (.CLK(clknet_leaf_4_clk),
    .D(_0345_),
    .RESET_B(net406),
    .Q(\mix1.data_o[25] ));
 sky130_fd_sc_hd__dfrtp_4 _8072_ (.CLK(clknet_leaf_5_clk),
    .D(_0346_),
    .RESET_B(net405),
    .Q(\mix1.data_o[26] ));
 sky130_fd_sc_hd__dfrtp_4 _8073_ (.CLK(clknet_leaf_4_clk),
    .D(_0347_),
    .RESET_B(net407),
    .Q(\mix1.data_o[27] ));
 sky130_fd_sc_hd__dfrtp_4 _8074_ (.CLK(clknet_leaf_5_clk),
    .D(_0348_),
    .RESET_B(net405),
    .Q(\mix1.data_o[28] ));
 sky130_fd_sc_hd__dfrtp_4 _8075_ (.CLK(clknet_leaf_3_clk),
    .D(_0349_),
    .RESET_B(net404),
    .Q(\mix1.data_o[29] ));
 sky130_fd_sc_hd__dfrtp_4 _8076_ (.CLK(clknet_leaf_3_clk),
    .D(_0350_),
    .RESET_B(net406),
    .Q(\mix1.data_o[30] ));
 sky130_fd_sc_hd__dfrtp_4 _8077_ (.CLK(clknet_leaf_5_clk),
    .D(_0351_),
    .RESET_B(net404),
    .Q(\mix1.data_o[31] ));
 sky130_fd_sc_hd__dfrtp_2 _8078_ (.CLK(clknet_leaf_1_clk),
    .D(_0352_),
    .RESET_B(net395),
    .Q(\mix1.data_o[32] ));
 sky130_fd_sc_hd__dfrtp_4 _8079_ (.CLK(clknet_leaf_1_clk),
    .D(_0353_),
    .RESET_B(net401),
    .Q(\mix1.data_o[33] ));
 sky130_fd_sc_hd__dfrtp_4 _8080_ (.CLK(clknet_leaf_12_clk),
    .D(_0354_),
    .RESET_B(net434),
    .Q(\mix1.data_o[34] ));
 sky130_fd_sc_hd__dfrtp_4 _8081_ (.CLK(clknet_leaf_14_clk),
    .D(_0355_),
    .RESET_B(net440),
    .Q(\mix1.data_o[35] ));
 sky130_fd_sc_hd__dfrtp_4 _8082_ (.CLK(clknet_leaf_14_clk),
    .D(_0356_),
    .RESET_B(net440),
    .Q(\mix1.data_o[36] ));
 sky130_fd_sc_hd__dfrtp_4 _8083_ (.CLK(clknet_leaf_14_clk),
    .D(_0357_),
    .RESET_B(net439),
    .Q(\mix1.data_o[37] ));
 sky130_fd_sc_hd__dfrtp_4 _8084_ (.CLK(clknet_leaf_15_clk),
    .D(_0358_),
    .RESET_B(net440),
    .Q(\mix1.data_o[38] ));
 sky130_fd_sc_hd__dfrtp_4 _8085_ (.CLK(clknet_leaf_14_clk),
    .D(_0359_),
    .RESET_B(net439),
    .Q(\mix1.data_o[39] ));
 sky130_fd_sc_hd__dfrtp_4 _8086_ (.CLK(clknet_leaf_13_clk),
    .D(_0360_),
    .RESET_B(net436),
    .Q(\mix1.data_o[40] ));
 sky130_fd_sc_hd__dfrtp_4 _8087_ (.CLK(clknet_leaf_13_clk),
    .D(_0361_),
    .RESET_B(net434),
    .Q(\mix1.data_o[41] ));
 sky130_fd_sc_hd__dfrtp_4 _8088_ (.CLK(clknet_leaf_13_clk),
    .D(_0362_),
    .RESET_B(net436),
    .Q(\mix1.data_o[42] ));
 sky130_fd_sc_hd__dfrtp_4 _8089_ (.CLK(clknet_leaf_11_clk),
    .D(_0363_),
    .RESET_B(net438),
    .Q(\mix1.data_o[43] ));
 sky130_fd_sc_hd__dfrtp_4 _8090_ (.CLK(clknet_leaf_12_clk),
    .D(_0364_),
    .RESET_B(net435),
    .Q(\mix1.data_o[44] ));
 sky130_fd_sc_hd__dfrtp_4 _8091_ (.CLK(clknet_leaf_13_clk),
    .D(_0365_),
    .RESET_B(net437),
    .Q(\mix1.data_o[45] ));
 sky130_fd_sc_hd__dfrtp_4 _8092_ (.CLK(clknet_leaf_12_clk),
    .D(_0366_),
    .RESET_B(net435),
    .Q(\mix1.data_o[46] ));
 sky130_fd_sc_hd__dfrtp_4 _8093_ (.CLK(clknet_leaf_13_clk),
    .D(_0367_),
    .RESET_B(net436),
    .Q(\mix1.data_o[47] ));
 sky130_fd_sc_hd__dfrtp_4 _8094_ (.CLK(clknet_leaf_14_clk),
    .D(_0368_),
    .RESET_B(net441),
    .Q(\mix1.data_o[48] ));
 sky130_fd_sc_hd__dfrtp_4 _8095_ (.CLK(clknet_leaf_17_clk),
    .D(_0369_),
    .RESET_B(net444),
    .Q(\mix1.data_o[49] ));
 sky130_fd_sc_hd__dfrtp_4 _8096_ (.CLK(clknet_leaf_15_clk),
    .D(_0370_),
    .RESET_B(net441),
    .Q(\mix1.data_o[50] ));
 sky130_fd_sc_hd__dfrtp_4 _8097_ (.CLK(clknet_leaf_20_clk),
    .D(_0371_),
    .RESET_B(net448),
    .Q(\mix1.data_o[51] ));
 sky130_fd_sc_hd__dfrtp_4 _8098_ (.CLK(clknet_leaf_20_clk),
    .D(_0372_),
    .RESET_B(net448),
    .Q(\mix1.data_o[52] ));
 sky130_fd_sc_hd__dfrtp_4 _8099_ (.CLK(clknet_leaf_17_clk),
    .D(_0373_),
    .RESET_B(net446),
    .Q(\mix1.data_o[53] ));
 sky130_fd_sc_hd__dfrtp_4 _8100_ (.CLK(clknet_leaf_16_clk),
    .D(_0374_),
    .RESET_B(net448),
    .Q(\mix1.data_o[54] ));
 sky130_fd_sc_hd__dfrtp_4 _8101_ (.CLK(clknet_leaf_17_clk),
    .D(_0375_),
    .RESET_B(net444),
    .Q(\mix1.data_o[55] ));
 sky130_fd_sc_hd__dfrtp_4 _8102_ (.CLK(clknet_leaf_6_clk),
    .D(_0376_),
    .RESET_B(net399),
    .Q(\mix1.data_o[56] ));
 sky130_fd_sc_hd__dfrtp_4 _8103_ (.CLK(clknet_leaf_5_clk),
    .D(_0377_),
    .RESET_B(net405),
    .Q(\mix1.data_o[57] ));
 sky130_fd_sc_hd__dfrtp_4 _8104_ (.CLK(clknet_leaf_6_clk),
    .D(_0378_),
    .RESET_B(net399),
    .Q(\mix1.data_o[58] ));
 sky130_fd_sc_hd__dfrtp_4 _8105_ (.CLK(clknet_leaf_5_clk),
    .D(_0379_),
    .RESET_B(net405),
    .Q(\mix1.data_o[59] ));
 sky130_fd_sc_hd__dfrtp_4 _8106_ (.CLK(clknet_leaf_6_clk),
    .D(_0380_),
    .RESET_B(net399),
    .Q(\mix1.data_o[60] ));
 sky130_fd_sc_hd__dfrtp_4 _8107_ (.CLK(clknet_leaf_0_clk),
    .D(_0381_),
    .RESET_B(net398),
    .Q(\mix1.data_o[61] ));
 sky130_fd_sc_hd__dfrtp_4 _8108_ (.CLK(clknet_leaf_0_clk),
    .D(_0382_),
    .RESET_B(net395),
    .Q(\mix1.data_o[62] ));
 sky130_fd_sc_hd__dfrtp_4 _8109_ (.CLK(clknet_leaf_0_clk),
    .D(_0383_),
    .RESET_B(net398),
    .Q(\mix1.data_o[63] ));
 sky130_fd_sc_hd__dfrtp_4 _8110_ (.CLK(clknet_leaf_1_clk),
    .D(_0384_),
    .RESET_B(net395),
    .Q(\mix1.data_o[64] ));
 sky130_fd_sc_hd__dfrtp_4 _8111_ (.CLK(clknet_leaf_1_clk),
    .D(_0385_),
    .RESET_B(net395),
    .Q(\mix1.data_o[65] ));
 sky130_fd_sc_hd__dfrtp_4 _8112_ (.CLK(clknet_leaf_2_clk),
    .D(_0386_),
    .RESET_B(net402),
    .Q(\mix1.data_o[66] ));
 sky130_fd_sc_hd__dfrtp_4 _8113_ (.CLK(clknet_leaf_12_clk),
    .D(_0387_),
    .RESET_B(net434),
    .Q(\mix1.data_o[67] ));
 sky130_fd_sc_hd__dfrtp_4 _8114_ (.CLK(clknet_leaf_1_clk),
    .D(_0388_),
    .RESET_B(net401),
    .Q(\mix1.data_o[68] ));
 sky130_fd_sc_hd__dfrtp_4 _8115_ (.CLK(clknet_leaf_2_clk),
    .D(_0389_),
    .RESET_B(net402),
    .Q(\mix1.data_o[69] ));
 sky130_fd_sc_hd__dfrtp_4 _8116_ (.CLK(clknet_leaf_12_clk),
    .D(_0390_),
    .RESET_B(net435),
    .Q(\mix1.data_o[70] ));
 sky130_fd_sc_hd__dfrtp_4 _8117_ (.CLK(clknet_leaf_2_clk),
    .D(_0391_),
    .RESET_B(net401),
    .Q(\mix1.data_o[71] ));
 sky130_fd_sc_hd__dfrtp_4 _8118_ (.CLK(clknet_leaf_2_clk),
    .D(_0392_),
    .RESET_B(net402),
    .Q(\mix1.data_o[72] ));
 sky130_fd_sc_hd__dfrtp_4 _8119_ (.CLK(clknet_leaf_2_clk),
    .D(_0393_),
    .RESET_B(net402),
    .Q(\mix1.data_o[73] ));
 sky130_fd_sc_hd__dfrtp_4 _8120_ (.CLK(clknet_leaf_2_clk),
    .D(_0394_),
    .RESET_B(net403),
    .Q(\mix1.data_o[74] ));
 sky130_fd_sc_hd__dfrtp_4 _8121_ (.CLK(clknet_leaf_4_clk),
    .D(_0395_),
    .RESET_B(net406),
    .Q(\mix1.data_o[75] ));
 sky130_fd_sc_hd__dfrtp_4 _8122_ (.CLK(clknet_leaf_0_clk),
    .D(_0396_),
    .RESET_B(net398),
    .Q(\mix1.data_o[76] ));
 sky130_fd_sc_hd__dfrtp_4 _8123_ (.CLK(clknet_leaf_3_clk),
    .D(_0397_),
    .RESET_B(net404),
    .Q(\mix1.data_o[77] ));
 sky130_fd_sc_hd__dfrtp_4 _8124_ (.CLK(clknet_leaf_1_clk),
    .D(_0398_),
    .RESET_B(net396),
    .Q(\mix1.data_o[78] ));
 sky130_fd_sc_hd__dfrtp_4 _8125_ (.CLK(clknet_leaf_6_clk),
    .D(_0399_),
    .RESET_B(net398),
    .Q(\mix1.data_o[79] ));
 sky130_fd_sc_hd__dfrtp_4 _8126_ (.CLK(clknet_leaf_17_clk),
    .D(_0400_),
    .RESET_B(net444),
    .Q(\mix1.data_o[80] ));
 sky130_fd_sc_hd__dfrtp_4 _8127_ (.CLK(clknet_leaf_17_clk),
    .D(_0401_),
    .RESET_B(net445),
    .Q(\mix1.data_o[81] ));
 sky130_fd_sc_hd__dfrtp_4 _8128_ (.CLK(clknet_leaf_17_clk),
    .D(_0402_),
    .RESET_B(net445),
    .Q(\mix1.data_o[82] ));
 sky130_fd_sc_hd__dfrtp_4 _8129_ (.CLK(clknet_leaf_20_clk),
    .D(_0403_),
    .RESET_B(net447),
    .Q(\mix1.data_o[83] ));
 sky130_fd_sc_hd__dfrtp_4 _8130_ (.CLK(clknet_leaf_19_clk),
    .D(_0404_),
    .RESET_B(net448),
    .Q(\mix1.data_o[84] ));
 sky130_fd_sc_hd__dfrtp_4 _8131_ (.CLK(clknet_leaf_19_clk),
    .D(_0405_),
    .RESET_B(net447),
    .Q(\mix1.data_o[85] ));
 sky130_fd_sc_hd__dfrtp_4 _8132_ (.CLK(clknet_leaf_19_clk),
    .D(_0406_),
    .RESET_B(net448),
    .Q(\mix1.data_o[86] ));
 sky130_fd_sc_hd__dfrtp_4 _8133_ (.CLK(clknet_leaf_17_clk),
    .D(_0407_),
    .RESET_B(net447),
    .Q(\mix1.data_o[87] ));
 sky130_fd_sc_hd__dfrtp_2 _8134_ (.CLK(clknet_leaf_6_clk),
    .D(_0408_),
    .RESET_B(net399),
    .Q(\mix1.data_o[88] ));
 sky130_fd_sc_hd__dfrtp_4 _8135_ (.CLK(clknet_leaf_86_clk),
    .D(_0409_),
    .RESET_B(net393),
    .Q(\mix1.data_o[89] ));
 sky130_fd_sc_hd__dfrtp_2 _8136_ (.CLK(clknet_leaf_81_clk),
    .D(_0410_),
    .RESET_B(net393),
    .Q(\mix1.data_o[90] ));
 sky130_fd_sc_hd__dfrtp_4 _8137_ (.CLK(clknet_leaf_87_clk),
    .D(_0411_),
    .RESET_B(net394),
    .Q(\mix1.data_o[91] ));
 sky130_fd_sc_hd__dfrtp_4 _8138_ (.CLK(clknet_leaf_87_clk),
    .D(_0412_),
    .RESET_B(net394),
    .Q(\mix1.data_o[92] ));
 sky130_fd_sc_hd__dfrtp_4 _8139_ (.CLK(clknet_leaf_87_clk),
    .D(_0413_),
    .RESET_B(net394),
    .Q(\mix1.data_o[93] ));
 sky130_fd_sc_hd__dfrtp_4 _8140_ (.CLK(clknet_leaf_0_clk),
    .D(_0414_),
    .RESET_B(net396),
    .Q(\mix1.data_o[94] ));
 sky130_fd_sc_hd__dfrtp_2 _8141_ (.CLK(clknet_leaf_0_clk),
    .D(_0415_),
    .RESET_B(net397),
    .Q(\mix1.data_o[95] ));
 sky130_fd_sc_hd__dfrtp_4 _8142_ (.CLK(clknet_leaf_18_clk),
    .D(_0416_),
    .RESET_B(net444),
    .Q(\mix1.data_o[96] ));
 sky130_fd_sc_hd__dfrtp_4 _8143_ (.CLK(clknet_leaf_18_clk),
    .D(_0417_),
    .RESET_B(net444),
    .Q(\mix1.data_o[97] ));
 sky130_fd_sc_hd__dfrtp_4 _8144_ (.CLK(clknet_leaf_18_clk),
    .D(_0418_),
    .RESET_B(net444),
    .Q(\mix1.data_o[98] ));
 sky130_fd_sc_hd__dfrtp_4 _8145_ (.CLK(clknet_leaf_15_clk),
    .D(_0419_),
    .RESET_B(net440),
    .Q(\mix1.data_o[99] ));
 sky130_fd_sc_hd__dfrtp_4 _8146_ (.CLK(clknet_leaf_14_clk),
    .D(_0420_),
    .RESET_B(net439),
    .Q(\mix1.data_o[100] ));
 sky130_fd_sc_hd__dfrtp_4 _8147_ (.CLK(clknet_leaf_14_clk),
    .D(_0421_),
    .RESET_B(net439),
    .Q(\mix1.data_o[101] ));
 sky130_fd_sc_hd__dfrtp_4 _8148_ (.CLK(clknet_leaf_15_clk),
    .D(_0422_),
    .RESET_B(net441),
    .Q(\mix1.data_o[102] ));
 sky130_fd_sc_hd__dfrtp_4 _8149_ (.CLK(clknet_leaf_13_clk),
    .D(_0423_),
    .RESET_B(net436),
    .Q(\mix1.data_o[103] ));
 sky130_fd_sc_hd__dfrtp_4 _8150_ (.CLK(clknet_leaf_1_clk),
    .D(_0424_),
    .RESET_B(net401),
    .Q(\mix1.data_o[104] ));
 sky130_fd_sc_hd__dfrtp_4 _8151_ (.CLK(clknet_leaf_1_clk),
    .D(_0425_),
    .RESET_B(net401),
    .Q(\mix1.data_o[105] ));
 sky130_fd_sc_hd__dfrtp_4 _8152_ (.CLK(clknet_leaf_3_clk),
    .D(_0426_),
    .RESET_B(net403),
    .Q(\mix1.data_o[106] ));
 sky130_fd_sc_hd__dfrtp_2 _8153_ (.CLK(clknet_leaf_3_clk),
    .D(_0427_),
    .RESET_B(net403),
    .Q(\mix1.data_o[107] ));
 sky130_fd_sc_hd__dfrtp_2 _8154_ (.CLK(clknet_leaf_3_clk),
    .D(_0428_),
    .RESET_B(net404),
    .Q(\mix1.data_o[108] ));
 sky130_fd_sc_hd__dfrtp_4 _8155_ (.CLK(clknet_leaf_4_clk),
    .D(_0429_),
    .RESET_B(net406),
    .Q(\mix1.data_o[109] ));
 sky130_fd_sc_hd__dfrtp_4 _8156_ (.CLK(clknet_leaf_5_clk),
    .D(_0430_),
    .RESET_B(net404),
    .Q(\mix1.data_o[110] ));
 sky130_fd_sc_hd__dfrtp_2 _8157_ (.CLK(clknet_leaf_5_clk),
    .D(_0431_),
    .RESET_B(net405),
    .Q(\mix1.data_o[111] ));
 sky130_fd_sc_hd__dfrtp_4 _8158_ (.CLK(clknet_leaf_19_clk),
    .D(_0432_),
    .RESET_B(net449),
    .Q(\mix1.data_o[112] ));
 sky130_fd_sc_hd__dfrtp_4 _8159_ (.CLK(clknet_leaf_19_clk),
    .D(_0433_),
    .RESET_B(net449),
    .Q(\mix1.data_o[113] ));
 sky130_fd_sc_hd__dfrtp_2 _8160_ (.CLK(clknet_leaf_21_clk),
    .D(_0434_),
    .RESET_B(net453),
    .Q(\mix1.data_o[114] ));
 sky130_fd_sc_hd__dfrtp_4 _8161_ (.CLK(clknet_leaf_19_clk),
    .D(_0435_),
    .RESET_B(net449),
    .Q(\mix1.data_o[115] ));
 sky130_fd_sc_hd__dfrtp_4 _8162_ (.CLK(clknet_leaf_19_clk),
    .D(_0436_),
    .RESET_B(net448),
    .Q(\mix1.data_o[116] ));
 sky130_fd_sc_hd__dfrtp_4 _8163_ (.CLK(clknet_leaf_19_clk),
    .D(_0437_),
    .RESET_B(net447),
    .Q(\mix1.data_o[117] ));
 sky130_fd_sc_hd__dfrtp_4 _8164_ (.CLK(clknet_leaf_19_clk),
    .D(_0438_),
    .RESET_B(net449),
    .Q(\mix1.data_o[118] ));
 sky130_fd_sc_hd__dfrtp_4 _8165_ (.CLK(clknet_leaf_16_clk),
    .D(_0439_),
    .RESET_B(net446),
    .Q(\mix1.data_o[119] ));
 sky130_fd_sc_hd__dfrtp_1 _8166_ (.CLK(clknet_leaf_7_clk),
    .D(_0440_),
    .RESET_B(net408),
    .Q(\mix1.data_o[120] ));
 sky130_fd_sc_hd__dfrtp_2 _8167_ (.CLK(clknet_leaf_7_clk),
    .D(_0441_),
    .RESET_B(net408),
    .Q(\mix1.data_o[121] ));
 sky130_fd_sc_hd__dfrtp_1 _8168_ (.CLK(clknet_leaf_7_clk),
    .D(_0442_),
    .RESET_B(net408),
    .Q(\mix1.data_o[122] ));
 sky130_fd_sc_hd__dfrtp_2 _8169_ (.CLK(clknet_leaf_87_clk),
    .D(_0443_),
    .RESET_B(net397),
    .Q(\mix1.data_o[123] ));
 sky130_fd_sc_hd__dfrtp_2 _8170_ (.CLK(clknet_leaf_87_clk),
    .D(_0444_),
    .RESET_B(net397),
    .Q(\mix1.data_o[124] ));
 sky130_fd_sc_hd__dfrtp_4 _8171_ (.CLK(clknet_leaf_87_clk),
    .D(_0445_),
    .RESET_B(net397),
    .Q(\mix1.data_o[125] ));
 sky130_fd_sc_hd__dfrtp_2 _8172_ (.CLK(clknet_leaf_87_clk),
    .D(_0446_),
    .RESET_B(net400),
    .Q(\mix1.data_o[126] ));
 sky130_fd_sc_hd__dfrtp_2 _8173_ (.CLK(clknet_leaf_0_clk),
    .D(_0447_),
    .RESET_B(net397),
    .Q(\mix1.data_o[127] ));
 sky130_fd_sc_hd__dfrtp_1 _8174_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0448_),
    .RESET_B(net458),
    .Q(\sub1.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8175_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0449_),
    .RESET_B(net458),
    .Q(\sub1.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8176_ (.CLK(clknet_leaf_54_clk),
    .D(_0450_),
    .RESET_B(net458),
    .Q(\sub1.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8177_ (.CLK(clknet_leaf_54_clk),
    .D(_0451_),
    .RESET_B(net458),
    .Q(\sub1.state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _8178_ (.CLK(clknet_leaf_29_clk),
    .D(_0452_),
    .RESET_B(net457),
    .Q(\sub1.state[4] ));
 sky130_fd_sc_hd__dfrtp_4 _8179_ (.CLK(clknet_leaf_23_clk),
    .D(_0453_),
    .RESET_B(net452),
    .Q(\sub1.data_o[80] ));
 sky130_fd_sc_hd__dfrtp_4 _8180_ (.CLK(clknet_leaf_35_clk),
    .D(_0454_),
    .RESET_B(net473),
    .Q(\sub1.data_o[81] ));
 sky130_fd_sc_hd__dfrtp_4 _8181_ (.CLK(clknet_leaf_35_clk),
    .D(_0455_),
    .RESET_B(net473),
    .Q(\sub1.data_o[82] ));
 sky130_fd_sc_hd__dfrtp_4 _8182_ (.CLK(clknet_leaf_35_clk),
    .D(_0456_),
    .RESET_B(net452),
    .Q(\sub1.data_o[83] ));
 sky130_fd_sc_hd__dfrtp_4 _8183_ (.CLK(clknet_leaf_34_clk),
    .D(_0457_),
    .RESET_B(net474),
    .Q(\sub1.data_o[84] ));
 sky130_fd_sc_hd__dfrtp_4 _8184_ (.CLK(clknet_leaf_35_clk),
    .D(_0458_),
    .RESET_B(net474),
    .Q(\sub1.data_o[85] ));
 sky130_fd_sc_hd__dfrtp_4 _8185_ (.CLK(clknet_leaf_34_clk),
    .D(_0459_),
    .RESET_B(net474),
    .Q(\sub1.data_o[86] ));
 sky130_fd_sc_hd__dfrtp_4 _8186_ (.CLK(clknet_leaf_34_clk),
    .D(_0460_),
    .RESET_B(net472),
    .Q(\sub1.data_o[87] ));
 sky130_fd_sc_hd__dfrtp_2 _8187_ (.CLK(clknet_leaf_83_clk),
    .D(_0461_),
    .RESET_B(net391),
    .Q(\sub1.data_o[88] ));
 sky130_fd_sc_hd__dfrtp_1 _8188_ (.CLK(clknet_leaf_73_clk),
    .D(_0462_),
    .RESET_B(net416),
    .Q(\sub1.data_o[89] ));
 sky130_fd_sc_hd__dfrtp_1 _8189_ (.CLK(clknet_leaf_83_clk),
    .D(_0463_),
    .RESET_B(net392),
    .Q(\sub1.data_o[90] ));
 sky130_fd_sc_hd__dfrtp_2 _8190_ (.CLK(clknet_leaf_73_clk),
    .D(_0464_),
    .RESET_B(net414),
    .Q(\sub1.data_o[91] ));
 sky130_fd_sc_hd__dfrtp_2 _8191_ (.CLK(clknet_leaf_73_clk),
    .D(_0465_),
    .RESET_B(net414),
    .Q(\sub1.data_o[92] ));
 sky130_fd_sc_hd__dfrtp_1 _8192_ (.CLK(clknet_leaf_73_clk),
    .D(_0466_),
    .RESET_B(net416),
    .Q(\sub1.data_o[93] ));
 sky130_fd_sc_hd__dfrtp_2 _8193_ (.CLK(clknet_leaf_83_clk),
    .D(_0467_),
    .RESET_B(net392),
    .Q(\sub1.data_o[94] ));
 sky130_fd_sc_hd__dfrtp_1 _8194_ (.CLK(clknet_leaf_81_clk),
    .D(_0468_),
    .RESET_B(net392),
    .Q(\sub1.data_o[95] ));
 sky130_fd_sc_hd__dfrtp_4 _8195_ (.CLK(clknet_leaf_21_clk),
    .D(_0469_),
    .RESET_B(net453),
    .Q(\sub1.data_o[96] ));
 sky130_fd_sc_hd__dfrtp_4 _8196_ (.CLK(clknet_leaf_25_clk),
    .D(_0470_),
    .RESET_B(net451),
    .Q(\sub1.data_o[97] ));
 sky130_fd_sc_hd__dfrtp_4 _8197_ (.CLK(clknet_leaf_21_clk),
    .D(_0471_),
    .RESET_B(net451),
    .Q(\sub1.data_o[98] ));
 sky130_fd_sc_hd__dfrtp_4 _8198_ (.CLK(clknet_leaf_25_clk),
    .D(_0472_),
    .RESET_B(net450),
    .Q(\sub1.data_o[99] ));
 sky130_fd_sc_hd__dfrtp_4 _8199_ (.CLK(clknet_leaf_20_clk),
    .D(_0473_),
    .RESET_B(net451),
    .Q(\sub1.data_o[100] ));
 sky130_fd_sc_hd__dfrtp_4 _8200_ (.CLK(clknet_leaf_25_clk),
    .D(_0474_),
    .RESET_B(net450),
    .Q(\sub1.data_o[101] ));
 sky130_fd_sc_hd__dfrtp_4 _8201_ (.CLK(clknet_leaf_25_clk),
    .D(_0475_),
    .RESET_B(net454),
    .Q(\sub1.data_o[102] ));
 sky130_fd_sc_hd__dfrtp_4 _8202_ (.CLK(clknet_leaf_20_clk),
    .D(_0476_),
    .RESET_B(net451),
    .Q(\sub1.data_o[103] ));
 sky130_fd_sc_hd__dfrtp_4 _8203_ (.CLK(clknet_leaf_8_clk),
    .D(\mix1.next_ready_o ),
    .RESET_B(net410),
    .Q(\mix1.ready_o ));
 sky130_fd_sc_hd__dfrtp_1 _8204_ (.CLK(clknet_leaf_62_clk),
    .D(_0477_),
    .RESET_B(net430),
    .Q(\ks1.key_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8205_ (.CLK(clknet_leaf_48_clk),
    .D(_0478_),
    .RESET_B(net462),
    .Q(\ks1.key_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8206_ (.CLK(clknet_leaf_62_clk),
    .D(_0479_),
    .RESET_B(net431),
    .Q(\ks1.key_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8207_ (.CLK(clknet_leaf_49_clk),
    .D(_0480_),
    .RESET_B(net462),
    .Q(\ks1.key_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8208_ (.CLK(clknet_leaf_62_clk),
    .D(_0481_),
    .RESET_B(net430),
    .Q(\ks1.key_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8209_ (.CLK(clknet_leaf_62_clk),
    .D(_0482_),
    .RESET_B(net431),
    .Q(\ks1.key_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8210_ (.CLK(clknet_leaf_47_clk),
    .D(_0483_),
    .RESET_B(net462),
    .Q(\ks1.key_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8211_ (.CLK(clknet_leaf_48_clk),
    .D(_0484_),
    .RESET_B(net461),
    .Q(\ks1.key_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8212_ (.CLK(clknet_leaf_49_clk),
    .D(_0485_),
    .RESET_B(net459),
    .Q(\ks1.key_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8213_ (.CLK(clknet_leaf_60_clk),
    .D(_0486_),
    .RESET_B(net428),
    .Q(\ks1.key_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8214_ (.CLK(clknet_leaf_49_clk),
    .D(_0487_),
    .RESET_B(net462),
    .Q(\ks1.key_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8215_ (.CLK(clknet_leaf_48_clk),
    .D(_0488_),
    .RESET_B(net461),
    .Q(\ks1.key_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8216_ (.CLK(clknet_leaf_60_clk),
    .D(_0489_),
    .RESET_B(net428),
    .Q(\ks1.key_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8217_ (.CLK(clknet_leaf_62_clk),
    .D(_0490_),
    .RESET_B(net431),
    .Q(\ks1.key_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8218_ (.CLK(clknet_leaf_48_clk),
    .D(_0491_),
    .RESET_B(net461),
    .Q(\ks1.key_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8219_ (.CLK(clknet_leaf_48_clk),
    .D(_0492_),
    .RESET_B(net462),
    .Q(\ks1.key_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8220_ (.CLK(clknet_leaf_46_clk),
    .D(_0493_),
    .RESET_B(net465),
    .Q(\ks1.key_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8221_ (.CLK(clknet_leaf_47_clk),
    .D(_0494_),
    .RESET_B(net465),
    .Q(\ks1.key_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8222_ (.CLK(clknet_leaf_47_clk),
    .D(_0495_),
    .RESET_B(net465),
    .Q(\ks1.key_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8223_ (.CLK(clknet_leaf_47_clk),
    .D(_0496_),
    .RESET_B(net465),
    .Q(\ks1.key_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8224_ (.CLK(clknet_leaf_46_clk),
    .D(_0497_),
    .RESET_B(net465),
    .Q(\ks1.key_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8225_ (.CLK(clknet_leaf_46_clk),
    .D(_0498_),
    .RESET_B(net463),
    .Q(\ks1.key_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8226_ (.CLK(clknet_leaf_47_clk),
    .D(_0499_),
    .RESET_B(net465),
    .Q(\ks1.key_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8227_ (.CLK(clknet_leaf_47_clk),
    .D(_0500_),
    .RESET_B(net465),
    .Q(\ks1.key_reg[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8228_ (.CLK(clknet_leaf_62_clk),
    .D(_0501_),
    .RESET_B(net431),
    .Q(\ks1.key_reg[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8229_ (.CLK(clknet_leaf_60_clk),
    .D(_0502_),
    .RESET_B(net428),
    .Q(\ks1.key_reg[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8230_ (.CLK(clknet_leaf_63_clk),
    .D(_0503_),
    .RESET_B(net430),
    .Q(\ks1.key_reg[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8231_ (.CLK(clknet_leaf_49_clk),
    .D(_0504_),
    .RESET_B(net459),
    .Q(\ks1.key_reg[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8232_ (.CLK(clknet_leaf_63_clk),
    .D(_0505_),
    .RESET_B(net430),
    .Q(\ks1.key_reg[28] ));
 sky130_fd_sc_hd__dfrtp_1 _8233_ (.CLK(clknet_leaf_49_clk),
    .D(_0506_),
    .RESET_B(net461),
    .Q(\ks1.key_reg[29] ));
 sky130_fd_sc_hd__dfrtp_1 _8234_ (.CLK(clknet_leaf_48_clk),
    .D(_0507_),
    .RESET_B(net461),
    .Q(\ks1.key_reg[30] ));
 sky130_fd_sc_hd__dfrtp_1 _8235_ (.CLK(clknet_leaf_63_clk),
    .D(_0508_),
    .RESET_B(net427),
    .Q(\ks1.key_reg[31] ));
 sky130_fd_sc_hd__dfrtp_1 _8236_ (.CLK(clknet_leaf_65_clk),
    .D(_0509_),
    .RESET_B(net425),
    .Q(\ks1.key_reg[32] ));
 sky130_fd_sc_hd__dfrtp_1 _8237_ (.CLK(clknet_leaf_63_clk),
    .D(_0510_),
    .RESET_B(net427),
    .Q(\ks1.key_reg[33] ));
 sky130_fd_sc_hd__dfrtp_1 _8238_ (.CLK(clknet_leaf_61_clk),
    .D(_0511_),
    .RESET_B(net429),
    .Q(\ks1.key_reg[34] ));
 sky130_fd_sc_hd__dfrtp_1 _8239_ (.CLK(clknet_leaf_45_clk),
    .D(_0512_),
    .RESET_B(net464),
    .Q(\ks1.key_reg[35] ));
 sky130_fd_sc_hd__dfrtp_1 _8240_ (.CLK(clknet_leaf_65_clk),
    .D(_0513_),
    .RESET_B(net426),
    .Q(\ks1.key_reg[36] ));
 sky130_fd_sc_hd__dfrtp_1 _8241_ (.CLK(clknet_leaf_64_clk),
    .D(_0514_),
    .RESET_B(net426),
    .Q(\ks1.key_reg[37] ));
 sky130_fd_sc_hd__dfrtp_1 _8242_ (.CLK(clknet_leaf_46_clk),
    .D(_0515_),
    .RESET_B(net466),
    .Q(\ks1.key_reg[38] ));
 sky130_fd_sc_hd__dfrtp_1 _8243_ (.CLK(clknet_leaf_45_clk),
    .D(_0516_),
    .RESET_B(net466),
    .Q(\ks1.key_reg[39] ));
 sky130_fd_sc_hd__dfrtp_1 _8244_ (.CLK(clknet_leaf_61_clk),
    .D(_0517_),
    .RESET_B(net429),
    .Q(\ks1.key_reg[40] ));
 sky130_fd_sc_hd__dfrtp_1 _8245_ (.CLK(clknet_leaf_64_clk),
    .D(_0518_),
    .RESET_B(net426),
    .Q(\ks1.key_reg[41] ));
 sky130_fd_sc_hd__dfrtp_1 _8246_ (.CLK(clknet_leaf_51_clk),
    .D(_0519_),
    .RESET_B(net460),
    .Q(\ks1.key_reg[42] ));
 sky130_fd_sc_hd__dfrtp_1 _8247_ (.CLK(clknet_leaf_50_clk),
    .D(_0520_),
    .RESET_B(net459),
    .Q(\ks1.key_reg[43] ));
 sky130_fd_sc_hd__dfrtp_1 _8248_ (.CLK(clknet_leaf_59_clk),
    .D(_0521_),
    .RESET_B(net425),
    .Q(\ks1.key_reg[44] ));
 sky130_fd_sc_hd__dfrtp_1 _8249_ (.CLK(clknet_leaf_62_clk),
    .D(_0522_),
    .RESET_B(net431),
    .Q(\ks1.key_reg[45] ));
 sky130_fd_sc_hd__dfrtp_1 _8250_ (.CLK(clknet_leaf_65_clk),
    .D(_0523_),
    .RESET_B(net424),
    .Q(\ks1.key_reg[46] ));
 sky130_fd_sc_hd__dfrtp_1 _8251_ (.CLK(clknet_leaf_49_clk),
    .D(_0524_),
    .RESET_B(net460),
    .Q(\ks1.key_reg[47] ));
 sky130_fd_sc_hd__dfrtp_1 _8252_ (.CLK(clknet_leaf_45_clk),
    .D(_0525_),
    .RESET_B(net464),
    .Q(\ks1.key_reg[48] ));
 sky130_fd_sc_hd__dfrtp_1 _8253_ (.CLK(clknet_leaf_45_clk),
    .D(_0526_),
    .RESET_B(net464),
    .Q(\ks1.key_reg[49] ));
 sky130_fd_sc_hd__dfrtp_1 _8254_ (.CLK(clknet_leaf_46_clk),
    .D(_0527_),
    .RESET_B(net466),
    .Q(\ks1.key_reg[50] ));
 sky130_fd_sc_hd__dfrtp_1 _8255_ (.CLK(clknet_leaf_43_clk),
    .D(_0528_),
    .RESET_B(net479),
    .Q(\ks1.key_reg[51] ));
 sky130_fd_sc_hd__dfrtp_1 _8256_ (.CLK(clknet_leaf_45_clk),
    .D(_0529_),
    .RESET_B(net464),
    .Q(\ks1.key_reg[52] ));
 sky130_fd_sc_hd__dfrtp_1 _8257_ (.CLK(clknet_leaf_45_clk),
    .D(_0530_),
    .RESET_B(net464),
    .Q(\ks1.key_reg[53] ));
 sky130_fd_sc_hd__dfrtp_1 _8258_ (.CLK(clknet_leaf_44_clk),
    .D(_0531_),
    .RESET_B(net479),
    .Q(\ks1.key_reg[54] ));
 sky130_fd_sc_hd__dfrtp_1 _8259_ (.CLK(clknet_leaf_45_clk),
    .D(_0532_),
    .RESET_B(net464),
    .Q(\ks1.key_reg[55] ));
 sky130_fd_sc_hd__dfrtp_1 _8260_ (.CLK(clknet_leaf_63_clk),
    .D(_0533_),
    .RESET_B(net430),
    .Q(\ks1.key_reg[56] ));
 sky130_fd_sc_hd__dfrtp_1 _8261_ (.CLK(clknet_leaf_60_clk),
    .D(_0534_),
    .RESET_B(net428),
    .Q(\ks1.key_reg[57] ));
 sky130_fd_sc_hd__dfrtp_1 _8262_ (.CLK(clknet_leaf_64_clk),
    .D(_0535_),
    .RESET_B(net426),
    .Q(\ks1.key_reg[58] ));
 sky130_fd_sc_hd__dfrtp_1 _8263_ (.CLK(clknet_leaf_59_clk),
    .D(_0536_),
    .RESET_B(net425),
    .Q(\ks1.key_reg[59] ));
 sky130_fd_sc_hd__dfrtp_1 _8264_ (.CLK(clknet_leaf_64_clk),
    .D(_0537_),
    .RESET_B(net426),
    .Q(\ks1.key_reg[60] ));
 sky130_fd_sc_hd__dfrtp_1 _8265_ (.CLK(clknet_leaf_60_clk),
    .D(_0538_),
    .RESET_B(net428),
    .Q(\ks1.key_reg[61] ));
 sky130_fd_sc_hd__dfrtp_1 _8266_ (.CLK(clknet_leaf_64_clk),
    .D(_0539_),
    .RESET_B(net426),
    .Q(\ks1.key_reg[62] ));
 sky130_fd_sc_hd__dfrtp_1 _8267_ (.CLK(clknet_leaf_66_clk),
    .D(_0540_),
    .RESET_B(net424),
    .Q(\ks1.key_reg[63] ));
 sky130_fd_sc_hd__dfrtp_1 _8268_ (.CLK(clknet_leaf_59_clk),
    .D(_0541_),
    .RESET_B(net425),
    .Q(\ks1.key_reg[64] ));
 sky130_fd_sc_hd__dfrtp_1 _8269_ (.CLK(clknet_leaf_63_clk),
    .D(_0542_),
    .RESET_B(net430),
    .Q(\ks1.key_reg[65] ));
 sky130_fd_sc_hd__dfrtp_1 _8270_ (.CLK(clknet_leaf_44_clk),
    .D(_0543_),
    .RESET_B(net479),
    .Q(\ks1.key_reg[66] ));
 sky130_fd_sc_hd__dfrtp_1 _8271_ (.CLK(clknet_leaf_44_clk),
    .D(_0544_),
    .RESET_B(net477),
    .Q(\ks1.key_reg[67] ));
 sky130_fd_sc_hd__dfrtp_1 _8272_ (.CLK(clknet_leaf_66_clk),
    .D(_0545_),
    .RESET_B(net419),
    .Q(\ks1.key_reg[68] ));
 sky130_fd_sc_hd__dfrtp_1 _8273_ (.CLK(clknet_leaf_66_clk),
    .D(_0546_),
    .RESET_B(net418),
    .Q(\ks1.key_reg[69] ));
 sky130_fd_sc_hd__dfrtp_1 _8274_ (.CLK(clknet_leaf_52_clk),
    .D(_0547_),
    .RESET_B(net464),
    .Q(\ks1.key_reg[70] ));
 sky130_fd_sc_hd__dfrtp_1 _8275_ (.CLK(clknet_leaf_43_clk),
    .D(_0548_),
    .RESET_B(net479),
    .Q(\ks1.key_reg[71] ));
 sky130_fd_sc_hd__dfrtp_1 _8276_ (.CLK(clknet_leaf_61_clk),
    .D(_0549_),
    .RESET_B(net429),
    .Q(\ks1.key_reg[72] ));
 sky130_fd_sc_hd__dfrtp_1 _8277_ (.CLK(clknet_leaf_67_clk),
    .D(_0550_),
    .RESET_B(net419),
    .Q(\ks1.key_reg[73] ));
 sky130_fd_sc_hd__dfrtp_1 _8278_ (.CLK(clknet_leaf_51_clk),
    .D(_0551_),
    .RESET_B(net463),
    .Q(\ks1.key_reg[74] ));
 sky130_fd_sc_hd__dfrtp_1 _8279_ (.CLK(clknet_leaf_60_clk),
    .D(_0552_),
    .RESET_B(net428),
    .Q(\ks1.key_reg[75] ));
 sky130_fd_sc_hd__dfrtp_1 _8280_ (.CLK(clknet_leaf_58_clk),
    .D(_0553_),
    .RESET_B(net425),
    .Q(\ks1.key_reg[76] ));
 sky130_fd_sc_hd__dfrtp_1 _8281_ (.CLK(clknet_leaf_67_clk),
    .D(_0554_),
    .RESET_B(net419),
    .Q(\ks1.key_reg[77] ));
 sky130_fd_sc_hd__dfrtp_1 _8282_ (.CLK(clknet_leaf_68_clk),
    .D(_0555_),
    .RESET_B(net418),
    .Q(\ks1.key_reg[78] ));
 sky130_fd_sc_hd__dfrtp_1 _8283_ (.CLK(clknet_leaf_65_clk),
    .D(_0556_),
    .RESET_B(net424),
    .Q(\ks1.key_reg[79] ));
 sky130_fd_sc_hd__dfrtp_1 _8284_ (.CLK(clknet_leaf_39_clk),
    .D(_0557_),
    .RESET_B(net477),
    .Q(\ks1.key_reg[80] ));
 sky130_fd_sc_hd__dfrtp_1 _8285_ (.CLK(clknet_leaf_44_clk),
    .D(_0558_),
    .RESET_B(net477),
    .Q(\ks1.key_reg[81] ));
 sky130_fd_sc_hd__dfrtp_1 _8286_ (.CLK(clknet_leaf_39_clk),
    .D(_0559_),
    .RESET_B(net477),
    .Q(\ks1.key_reg[82] ));
 sky130_fd_sc_hd__dfrtp_1 _8287_ (.CLK(clknet_leaf_44_clk),
    .D(_0560_),
    .RESET_B(net479),
    .Q(\ks1.key_reg[83] ));
 sky130_fd_sc_hd__dfrtp_1 _8288_ (.CLK(clknet_leaf_58_clk),
    .D(_0561_),
    .RESET_B(net421),
    .Q(\ks1.key_reg[84] ));
 sky130_fd_sc_hd__dfrtp_1 _8289_ (.CLK(clknet_leaf_39_clk),
    .D(_0562_),
    .RESET_B(net477),
    .Q(\ks1.key_reg[85] ));
 sky130_fd_sc_hd__dfrtp_1 _8290_ (.CLK(clknet_leaf_38_clk),
    .D(_0563_),
    .RESET_B(net478),
    .Q(\ks1.key_reg[86] ));
 sky130_fd_sc_hd__dfrtp_1 _8291_ (.CLK(clknet_leaf_39_clk),
    .D(_0564_),
    .RESET_B(net478),
    .Q(\ks1.key_reg[87] ));
 sky130_fd_sc_hd__dfrtp_1 _8292_ (.CLK(clknet_leaf_59_clk),
    .D(_0565_),
    .RESET_B(net424),
    .Q(\ks1.key_reg[88] ));
 sky130_fd_sc_hd__dfrtp_1 _8293_ (.CLK(clknet_leaf_68_clk),
    .D(_0566_),
    .RESET_B(net418),
    .Q(\ks1.key_reg[89] ));
 sky130_fd_sc_hd__dfrtp_1 _8294_ (.CLK(clknet_leaf_67_clk),
    .D(_0567_),
    .RESET_B(net419),
    .Q(\ks1.key_reg[90] ));
 sky130_fd_sc_hd__dfrtp_1 _8295_ (.CLK(clknet_leaf_68_clk),
    .D(_0568_),
    .RESET_B(net418),
    .Q(\ks1.key_reg[91] ));
 sky130_fd_sc_hd__dfrtp_1 _8296_ (.CLK(clknet_leaf_69_clk),
    .D(_0569_),
    .RESET_B(net415),
    .Q(\ks1.key_reg[92] ));
 sky130_fd_sc_hd__dfrtp_1 _8297_ (.CLK(clknet_leaf_69_clk),
    .D(_0570_),
    .RESET_B(net415),
    .Q(\ks1.key_reg[93] ));
 sky130_fd_sc_hd__dfrtp_1 _8298_ (.CLK(clknet_leaf_66_clk),
    .D(_0571_),
    .RESET_B(net424),
    .Q(\ks1.key_reg[94] ));
 sky130_fd_sc_hd__dfrtp_1 _8299_ (.CLK(clknet_leaf_69_clk),
    .D(_0572_),
    .RESET_B(net415),
    .Q(\ks1.key_reg[95] ));
 sky130_fd_sc_hd__dfrtp_1 _8300_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0573_),
    .RESET_B(net480),
    .Q(\ks1.key_reg[96] ));
 sky130_fd_sc_hd__dfrtp_1 _8301_ (.CLK(clknet_leaf_37_clk),
    .D(_0574_),
    .RESET_B(net476),
    .Q(\ks1.key_reg[97] ));
 sky130_fd_sc_hd__dfrtp_1 _8302_ (.CLK(clknet_leaf_36_clk),
    .D(_0575_),
    .RESET_B(net476),
    .Q(\ks1.key_reg[98] ));
 sky130_fd_sc_hd__dfrtp_1 _8303_ (.CLK(clknet_leaf_37_clk),
    .D(_0576_),
    .RESET_B(net480),
    .Q(\ks1.key_reg[99] ));
 sky130_fd_sc_hd__dfrtp_1 _8304_ (.CLK(clknet_leaf_68_clk),
    .D(_0577_),
    .RESET_B(net418),
    .Q(\ks1.key_reg[100] ));
 sky130_fd_sc_hd__dfrtp_1 _8305_ (.CLK(clknet_leaf_68_clk),
    .D(_0578_),
    .RESET_B(net418),
    .Q(\ks1.key_reg[101] ));
 sky130_fd_sc_hd__dfrtp_1 _8306_ (.CLK(clknet_leaf_37_clk),
    .D(_0579_),
    .RESET_B(net475),
    .Q(\ks1.key_reg[102] ));
 sky130_fd_sc_hd__dfrtp_1 _8307_ (.CLK(clknet_leaf_40_clk),
    .D(_0580_),
    .RESET_B(net480),
    .Q(\ks1.key_reg[103] ));
 sky130_fd_sc_hd__dfrtp_1 _8308_ (.CLK(clknet_leaf_59_clk),
    .D(_0581_),
    .RESET_B(net425),
    .Q(\ks1.key_reg[104] ));
 sky130_fd_sc_hd__dfrtp_1 _8309_ (.CLK(clknet_leaf_66_clk),
    .D(_0582_),
    .RESET_B(net419),
    .Q(\ks1.key_reg[105] ));
 sky130_fd_sc_hd__dfrtp_1 _8310_ (.CLK(clknet_leaf_59_clk),
    .D(_0583_),
    .RESET_B(net425),
    .Q(\ks1.key_reg[106] ));
 sky130_fd_sc_hd__dfrtp_1 _8311_ (.CLK(clknet_leaf_59_clk),
    .D(_0584_),
    .RESET_B(net425),
    .Q(\ks1.key_reg[107] ));
 sky130_fd_sc_hd__dfrtp_1 _8312_ (.CLK(clknet_leaf_58_clk),
    .D(_0585_),
    .RESET_B(net424),
    .Q(\ks1.key_reg[108] ));
 sky130_fd_sc_hd__dfrtp_1 _8313_ (.CLK(clknet_leaf_66_clk),
    .D(_0586_),
    .RESET_B(net419),
    .Q(\ks1.key_reg[109] ));
 sky130_fd_sc_hd__dfrtp_1 _8314_ (.CLK(clknet_leaf_66_clk),
    .D(_0587_),
    .RESET_B(net419),
    .Q(\ks1.key_reg[110] ));
 sky130_fd_sc_hd__dfrtp_1 _8315_ (.CLK(clknet_leaf_75_clk),
    .D(_0588_),
    .RESET_B(net421),
    .Q(\ks1.key_reg[111] ));
 sky130_fd_sc_hd__dfrtp_1 _8316_ (.CLK(clknet_leaf_75_clk),
    .D(_0589_),
    .RESET_B(net415),
    .Q(\ks1.key_reg[112] ));
 sky130_fd_sc_hd__dfrtp_1 _8317_ (.CLK(clknet_leaf_40_clk),
    .D(_0590_),
    .RESET_B(net478),
    .Q(\ks1.key_reg[113] ));
 sky130_fd_sc_hd__dfrtp_1 _8318_ (.CLK(clknet_leaf_38_clk),
    .D(_0591_),
    .RESET_B(net475),
    .Q(\ks1.key_reg[114] ));
 sky130_fd_sc_hd__dfrtp_1 _8319_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0592_),
    .RESET_B(net480),
    .Q(\ks1.key_reg[115] ));
 sky130_fd_sc_hd__dfrtp_1 _8320_ (.CLK(clknet_leaf_75_clk),
    .D(_0593_),
    .RESET_B(net421),
    .Q(\ks1.key_reg[116] ));
 sky130_fd_sc_hd__dfrtp_1 _8321_ (.CLK(clknet_leaf_44_clk),
    .D(_0594_),
    .RESET_B(net478),
    .Q(\ks1.key_reg[117] ));
 sky130_fd_sc_hd__dfrtp_1 _8322_ (.CLK(clknet_leaf_38_clk),
    .D(_0595_),
    .RESET_B(net471),
    .Q(\ks1.key_reg[118] ));
 sky130_fd_sc_hd__dfrtp_1 _8323_ (.CLK(clknet_leaf_40_clk),
    .D(_0596_),
    .RESET_B(net479),
    .Q(\ks1.key_reg[119] ));
 sky130_fd_sc_hd__dfrtp_1 _8324_ (.CLK(clknet_leaf_66_clk),
    .D(_0597_),
    .RESET_B(net424),
    .Q(\ks1.key_reg[120] ));
 sky130_fd_sc_hd__dfrtp_1 _8325_ (.CLK(clknet_leaf_74_clk),
    .D(_0598_),
    .RESET_B(net416),
    .Q(\ks1.key_reg[121] ));
 sky130_fd_sc_hd__dfrtp_1 _8326_ (.CLK(clknet_leaf_68_clk),
    .D(_0599_),
    .RESET_B(net418),
    .Q(\ks1.key_reg[122] ));
 sky130_fd_sc_hd__dfrtp_1 _8327_ (.CLK(clknet_leaf_68_clk),
    .D(_0600_),
    .RESET_B(net419),
    .Q(\ks1.key_reg[123] ));
 sky130_fd_sc_hd__dfrtp_1 _8328_ (.CLK(clknet_leaf_74_clk),
    .D(_0601_),
    .RESET_B(net416),
    .Q(\ks1.key_reg[124] ));
 sky130_fd_sc_hd__dfrtp_1 _8329_ (.CLK(clknet_leaf_69_clk),
    .D(_0602_),
    .RESET_B(net415),
    .Q(\ks1.key_reg[125] ));
 sky130_fd_sc_hd__dfrtp_1 _8330_ (.CLK(clknet_leaf_74_clk),
    .D(_0603_),
    .RESET_B(net416),
    .Q(\ks1.key_reg[126] ));
 sky130_fd_sc_hd__dfrtp_1 _8331_ (.CLK(clknet_leaf_74_clk),
    .D(_0604_),
    .RESET_B(net415),
    .Q(\ks1.key_reg[127] ));
 sky130_fd_sc_hd__dfrtp_2 _8332_ (.CLK(clknet_leaf_80_clk),
    .D(_0605_),
    .RESET_B(net408),
    .Q(\mix1.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8333_ (.CLK(clknet_leaf_0_clk),
    .D(_0606_),
    .RESET_B(net396),
    .Q(\mix1.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8334_ (.CLK(clknet_leaf_18_clk),
    .D(_0607_),
    .RESET_B(net445),
    .Q(\mix1.data_reg[96] ));
 sky130_fd_sc_hd__dfrtp_1 _8335_ (.CLK(clknet_leaf_18_clk),
    .D(_0608_),
    .RESET_B(net440),
    .Q(\mix1.data_reg[97] ));
 sky130_fd_sc_hd__dfrtp_1 _8336_ (.CLK(clknet_leaf_18_clk),
    .D(_0609_),
    .RESET_B(net444),
    .Q(\mix1.data_reg[98] ));
 sky130_fd_sc_hd__dfrtp_1 _8337_ (.CLK(clknet_leaf_15_clk),
    .D(_0610_),
    .RESET_B(net440),
    .Q(\mix1.data_reg[99] ));
 sky130_fd_sc_hd__dfrtp_1 _8338_ (.CLK(clknet_leaf_14_clk),
    .D(_0611_),
    .RESET_B(net439),
    .Q(\mix1.data_reg[100] ));
 sky130_fd_sc_hd__dfrtp_1 _8339_ (.CLK(clknet_leaf_14_clk),
    .D(_0612_),
    .RESET_B(net439),
    .Q(\mix1.data_reg[101] ));
 sky130_fd_sc_hd__dfrtp_1 _8340_ (.CLK(clknet_leaf_15_clk),
    .D(_0613_),
    .RESET_B(net440),
    .Q(\mix1.data_reg[102] ));
 sky130_fd_sc_hd__dfrtp_1 _8341_ (.CLK(clknet_leaf_13_clk),
    .D(_0614_),
    .RESET_B(net436),
    .Q(\mix1.data_reg[103] ));
 sky130_fd_sc_hd__dfrtp_1 _8342_ (.CLK(clknet_leaf_2_clk),
    .D(_0615_),
    .RESET_B(net401),
    .Q(\mix1.data_reg[104] ));
 sky130_fd_sc_hd__dfrtp_1 _8343_ (.CLK(clknet_leaf_2_clk),
    .D(_0616_),
    .RESET_B(net401),
    .Q(\mix1.data_reg[105] ));
 sky130_fd_sc_hd__dfrtp_1 _8344_ (.CLK(clknet_leaf_3_clk),
    .D(_0617_),
    .RESET_B(net403),
    .Q(\mix1.data_reg[106] ));
 sky130_fd_sc_hd__dfrtp_1 _8345_ (.CLK(clknet_leaf_3_clk),
    .D(_0618_),
    .RESET_B(net403),
    .Q(\mix1.data_reg[107] ));
 sky130_fd_sc_hd__dfrtp_1 _8346_ (.CLK(clknet_leaf_3_clk),
    .D(_0619_),
    .RESET_B(net403),
    .Q(\mix1.data_reg[108] ));
 sky130_fd_sc_hd__dfrtp_1 _8347_ (.CLK(clknet_leaf_3_clk),
    .D(_0620_),
    .RESET_B(net406),
    .Q(\mix1.data_reg[109] ));
 sky130_fd_sc_hd__dfrtp_1 _8348_ (.CLK(clknet_leaf_3_clk),
    .D(_0621_),
    .RESET_B(net403),
    .Q(\mix1.data_reg[110] ));
 sky130_fd_sc_hd__dfrtp_1 _8349_ (.CLK(clknet_leaf_3_clk),
    .D(_0622_),
    .RESET_B(net404),
    .Q(\mix1.data_reg[111] ));
 sky130_fd_sc_hd__dfrtp_1 _8350_ (.CLK(clknet_leaf_19_clk),
    .D(_0623_),
    .RESET_B(net449),
    .Q(\mix1.data_reg[112] ));
 sky130_fd_sc_hd__dfrtp_1 _8351_ (.CLK(clknet_leaf_19_clk),
    .D(_0624_),
    .RESET_B(net449),
    .Q(\mix1.data_reg[113] ));
 sky130_fd_sc_hd__dfrtp_1 _8352_ (.CLK(clknet_leaf_19_clk),
    .D(_0625_),
    .RESET_B(net449),
    .Q(\mix1.data_reg[114] ));
 sky130_fd_sc_hd__dfrtp_1 _8353_ (.CLK(clknet_leaf_19_clk),
    .D(_0626_),
    .RESET_B(net455),
    .Q(\mix1.data_reg[115] ));
 sky130_fd_sc_hd__dfrtp_1 _8354_ (.CLK(clknet_leaf_19_clk),
    .D(_0627_),
    .RESET_B(net448),
    .Q(\mix1.data_reg[116] ));
 sky130_fd_sc_hd__dfrtp_1 _8355_ (.CLK(clknet_leaf_17_clk),
    .D(_0628_),
    .RESET_B(net447),
    .Q(\mix1.data_reg[117] ));
 sky130_fd_sc_hd__dfrtp_1 _8356_ (.CLK(clknet_leaf_19_clk),
    .D(_0629_),
    .RESET_B(net447),
    .Q(\mix1.data_reg[118] ));
 sky130_fd_sc_hd__dfrtp_1 _8357_ (.CLK(clknet_leaf_16_clk),
    .D(_0630_),
    .RESET_B(net446),
    .Q(\mix1.data_reg[119] ));
 sky130_fd_sc_hd__dfrtp_1 _8358_ (.CLK(clknet_leaf_7_clk),
    .D(_0631_),
    .RESET_B(net400),
    .Q(\mix1.data_reg[120] ));
 sky130_fd_sc_hd__dfrtp_1 _8359_ (.CLK(clknet_leaf_87_clk),
    .D(_0632_),
    .RESET_B(net400),
    .Q(\mix1.data_reg[121] ));
 sky130_fd_sc_hd__dfrtp_1 _8360_ (.CLK(clknet_leaf_87_clk),
    .D(_0633_),
    .RESET_B(net394),
    .Q(\mix1.data_reg[122] ));
 sky130_fd_sc_hd__dfrtp_1 _8361_ (.CLK(clknet_leaf_87_clk),
    .D(_0634_),
    .RESET_B(net394),
    .Q(\mix1.data_reg[123] ));
 sky130_fd_sc_hd__dfrtp_1 _8362_ (.CLK(clknet_leaf_87_clk),
    .D(_0635_),
    .RESET_B(net400),
    .Q(\mix1.data_reg[124] ));
 sky130_fd_sc_hd__dfrtp_1 _8363_ (.CLK(clknet_leaf_87_clk),
    .D(_0636_),
    .RESET_B(net397),
    .Q(\mix1.data_reg[125] ));
 sky130_fd_sc_hd__dfrtp_1 _8364_ (.CLK(clknet_leaf_0_clk),
    .D(_0637_),
    .RESET_B(net397),
    .Q(\mix1.data_reg[126] ));
 sky130_fd_sc_hd__dfrtp_1 _8365_ (.CLK(clknet_leaf_0_clk),
    .D(_0638_),
    .RESET_B(net397),
    .Q(\mix1.data_reg[127] ));
 sky130_fd_sc_hd__dfrtp_4 _8366_ (.CLK(clknet_leaf_29_clk),
    .D(_0639_),
    .RESET_B(net457),
    .Q(\sub1.data_o[104] ));
 sky130_fd_sc_hd__dfrtp_4 _8367_ (.CLK(clknet_leaf_29_clk),
    .D(_0640_),
    .RESET_B(net457),
    .Q(\sub1.data_o[105] ));
 sky130_fd_sc_hd__dfrtp_4 _8368_ (.CLK(clknet_leaf_32_clk),
    .D(_0641_),
    .RESET_B(net457),
    .Q(\sub1.data_o[106] ));
 sky130_fd_sc_hd__dfrtp_4 _8369_ (.CLK(clknet_leaf_29_clk),
    .D(_0642_),
    .RESET_B(net457),
    .Q(\sub1.data_o[107] ));
 sky130_fd_sc_hd__dfrtp_4 _8370_ (.CLK(clknet_leaf_29_clk),
    .D(_0643_),
    .RESET_B(net457),
    .Q(\sub1.data_o[108] ));
 sky130_fd_sc_hd__dfrtp_4 _8371_ (.CLK(clknet_leaf_29_clk),
    .D(_0644_),
    .RESET_B(net457),
    .Q(\sub1.data_o[109] ));
 sky130_fd_sc_hd__dfrtp_4 _8372_ (.CLK(clknet_leaf_33_clk),
    .D(_0645_),
    .RESET_B(net469),
    .Q(\sub1.data_o[110] ));
 sky130_fd_sc_hd__dfrtp_4 _8373_ (.CLK(clknet_leaf_32_clk),
    .D(_0646_),
    .RESET_B(net469),
    .Q(\sub1.data_o[111] ));
 sky130_fd_sc_hd__dfrtp_4 _8374_ (.CLK(clknet_leaf_64_clk),
    .D(_0647_),
    .RESET_B(net427),
    .Q(\ks1.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8375_ (.CLK(clknet_leaf_65_clk),
    .D(_0648_),
    .RESET_B(net427),
    .Q(\ks1.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8376_ (.CLK(clknet_leaf_65_clk),
    .D(_0649_),
    .RESET_B(net427),
    .Q(\ks1.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8377_ (.CLK(clknet_leaf_68_clk),
    .D(\ks1.next_ready_o ),
    .RESET_B(net418),
    .Q(\ks1.ready_o ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout390 (.A(net393),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_4 fanout391 (.A(net393),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_4 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_2 fanout393 (.A(net394),
    .X(net393));
 sky130_fd_sc_hd__buf_4 fanout394 (.A(net411),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_4 fanout395 (.A(net396),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_2 fanout396 (.A(net411),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_4 fanout397 (.A(net400),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_4 fanout398 (.A(net400),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_2 fanout399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__buf_2 fanout400 (.A(net411),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_4 fanout401 (.A(net403),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_4 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_4 fanout403 (.A(net407),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_4 fanout404 (.A(net407),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_2 fanout405 (.A(net407),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_4 fanout406 (.A(net407),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 fanout407 (.A(net411),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_4 fanout408 (.A(net410),
    .X(net408));
 sky130_fd_sc_hd__buf_2 fanout409 (.A(net410),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_4 fanout410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__buf_2 fanout411 (.A(net482),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_4 fanout412 (.A(net417),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_2 fanout413 (.A(net417),
    .X(net413));
 sky130_fd_sc_hd__buf_4 fanout414 (.A(net416),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_4 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_4 fanout416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_2 fanout417 (.A(net420),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_4 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_4 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__buf_2 fanout420 (.A(net433),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_4 fanout421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_4 fanout422 (.A(net433),
    .X(net422));
 sky130_fd_sc_hd__buf_4 fanout423 (.A(net433),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_4 fanout424 (.A(net432),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_4 fanout425 (.A(net432),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_4 fanout426 (.A(net432),
    .X(net426));
 sky130_fd_sc_hd__buf_2 fanout427 (.A(net432),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_4 fanout428 (.A(net432),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 fanout429 (.A(net432),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_4 fanout430 (.A(net432),
    .X(net430));
 sky130_fd_sc_hd__buf_2 fanout431 (.A(net432),
    .X(net431));
 sky130_fd_sc_hd__buf_2 fanout432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_2 fanout433 (.A(net482),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_4 fanout434 (.A(net437),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_2 fanout435 (.A(net437),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_4 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_2 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 fanout438 (.A(net455),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_4 fanout439 (.A(net441),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_4 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_2 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_2 fanout442 (.A(net455),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_4 fanout443 (.A(net455),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_4 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__buf_2 fanout445 (.A(net449),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_4 fanout446 (.A(net448),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_4 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_4 fanout449 (.A(net455),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_4 fanout450 (.A(net454),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 fanout451 (.A(net454),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_4 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__buf_4 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_2 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_4 fanout455 (.A(net482),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_4 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_4 fanout457 (.A(net468),
    .X(net457));
 sky130_fd_sc_hd__buf_4 fanout458 (.A(net468),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 fanout459 (.A(net467),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_2 fanout460 (.A(net467),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_4 fanout461 (.A(net467),
    .X(net461));
 sky130_fd_sc_hd__buf_2 fanout462 (.A(net467),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_4 fanout463 (.A(net466),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_4 fanout464 (.A(net466),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_2 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_2 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__buf_2 fanout468 (.A(net482),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_4 fanout469 (.A(net472),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_4 fanout470 (.A(net472),
    .X(net470));
 sky130_fd_sc_hd__buf_2 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_2 fanout472 (.A(net481),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_4 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_4 fanout474 (.A(net481),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_4 fanout475 (.A(net481),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_4 fanout476 (.A(net481),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_4 fanout477 (.A(net478),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_4 fanout478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_4 fanout479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_4 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_2 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_4 fanout482 (.A(net259),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(first_round_reg),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\ks1.key_reg[79] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\mix1.data_reg[69] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\mix1.data_reg[37] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\mix1.data_reg[65] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\mix1.data_reg[66] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\mix1.data_reg[125] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\mix1.data_reg[36] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\mix1.data_reg[84] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\mix1.data_reg[54] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\mix1.data_reg[109] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\mix1.data_reg[92] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\ks1.key_reg[63] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\mix1.data_reg[114] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\mix1.data_reg[124] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\mix1.data_reg[50] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\mix1.data_reg[121] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\mix1.data_reg[72] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\mix1.data_reg[79] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\mix1.data_reg[108] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\mix1.data_reg[63] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\mix1.data_reg[48] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\mix1.data_reg[91] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\ks1.key_reg[44] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\mix1.data_reg[78] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\mix1.data_reg[61] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\mix1.data_reg[60] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\mix1.data_reg[33] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\mix1.data_reg[71] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\ks1.key_reg[48] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\mix1.data_reg[32] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\mix1.data_reg[44] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\mix1.data_reg[118] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\mix1.data_reg[87] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\ks1.key_reg[10] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\ks1.key_reg[25] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\mix1.data_reg[77] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\ks1.key_reg[73] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\ks1.key_reg[95] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\mix1.data_reg[119] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\ks1.key_reg[51] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\mix1.data_reg[47] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\mix1.data_reg[46] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\ks1.key_reg[70] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\ks1.key_reg[91] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\ks1.key_reg[20] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\mix1.data_reg[115] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\mix1.data_reg[55] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\ks1.key_reg[27] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\ks1.key_reg[12] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\ks1.key_reg[71] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\mix1.data_reg[111] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\ks1.key_reg[64] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\ks1.key_reg[110] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\ks1.key_reg[93] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\ks1.key_reg[88] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\sub1.state[4] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\ks1.key_reg[66] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\mix1.data_reg[89] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\ks1.key_reg[68] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\ks1.key_reg[81] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\ks1.key_reg[43] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\ks1.key_reg[102] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\ks1.key_reg[53] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\ks1.key_reg[38] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\ks1.key_reg[87] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\ks1.key_reg[50] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\ks1.key_reg[21] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\ks1.key_reg[83] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\ks1.key_reg[30] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\ks1.key_reg[92] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\ks1.key_reg[47] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\ks1.key_reg[85] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\ks1.key_reg[49] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\ks1.key_reg[39] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\ks1.key_reg[14] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\ks1.key_reg[8] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\ks1.key_reg[75] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\ks1.key_reg[19] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\ks1.key_reg[72] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\ks1.key_reg[54] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\ks1.key_reg[32] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\ks1.key_reg[76] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\ks1.key_reg[69] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\ks1.key_reg[33] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\ks1.key_reg[105] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\ks1.key_reg[119] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\ks1.key_reg[112] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\ks1.key_reg[26] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\ks1.key_reg[13] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\ks1.key_reg[94] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\ks1.key_reg[34] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\ks1.key_reg[84] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\ks1.key_reg[90] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\ks1.key_reg[45] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\ks1.key_reg[65] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\ks1.key_reg[114] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\ks1.key_reg[103] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\ks1.key_reg[118] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\ks1.key_reg[78] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\ks1.key_reg[59] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\ks1.key_reg[99] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\ks1.key_reg[113] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\ks1.key_reg[9] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\ks1.key_reg[29] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\ks1.key_reg[80] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\ks1.key_reg[36] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\ks1.key_reg[97] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\ks1.key_reg[111] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\ks1.key_reg[100] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\ks1.key_reg[121] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\ks1.key_reg[58] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\ks1.key_reg[3] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\ks1.col[25] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\ks1.key_reg[52] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\ks1.key_reg[67] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\ks1.key_reg[122] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\ks1.col[27] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\ks1.key_reg[106] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\ks1.key_reg[74] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\ks1.key_reg[89] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\ks1.key_reg[117] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\ks1.key_reg[126] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\ks1.key_reg[23] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\ks1.key_reg[42] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\ks1.key_reg[31] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\ks1.col[17] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\ks1.key_reg[109] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\ks1.key_reg[101] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\ks1.key_reg[55] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\ks1.key_reg[37] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\ks1.key_reg[28] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\ks1.key_reg[86] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\mix1.data_reg[110] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\ks1.key_reg[22] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\ks1.key_reg[35] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\ks1.key_reg[98] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\ks1.key_reg[125] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\ks1.key_reg[82] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\mix1.data_reg[110] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\ks1.key_reg[41] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\ks1.key_reg[11] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\ks1.key_reg[123] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\ks1.key_reg[108] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\ks1.key_reg[7] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\ks1.key_reg[15] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\ks1.key_reg[5] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\ks1.key_reg[62] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\ks1.key_reg[0] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\ks1.key_reg[6] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\ks1.key_reg[56] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\ks1.key_reg[16] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\ks1.key_reg[4] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\ks1.key_reg[17] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\ks1.key_reg[1] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\ks1.key_reg[107] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\ks1.key_reg[120] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\mix1.data_reg[67] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\ks1.key_reg[60] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\ks1.key_reg[2] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\ks1.key_reg[18] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\mix1.data_reg[80] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\mix1.data_reg[85] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\mix1.data_reg[117] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\mix1.data_reg[93] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\ks1.state[1] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\mix1.data_reg[68] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\mix1.data_reg[59] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\mix1.data_reg[41] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\ks1.key_reg[61] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\mix1.data_reg[76] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\mix1.data_reg[45] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\mix1.data_reg[73] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\mix1.data_reg[62] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\mix1.data_reg[51] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\mix1.data_reg[105] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\mix1.data_reg[96] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\mix1.data_reg[104] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\mix1.data_reg[126] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\mix1.data_reg[99] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\ks1.key_reg[104] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\mix1.data_reg[97] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\mix1.data_reg[98] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\mix1.data_reg[38] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\mix1.data_reg[53] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\mix1.data_reg[40] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\mix1.data_reg[94] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\mix1.data_reg[81] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\mix1.data_reg[82] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\mix1.data_reg[35] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\mix1.data_reg[102] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\ks1.key_reg[40] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\mix1.data_reg[56] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\mix1.data_reg[75] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\mix1.data_reg[95] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\mix1.data_reg[74] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\mix1.data_reg[88] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\mix1.data_reg[42] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\mix1.data_reg[58] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\mix1.data_reg[34] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\mix1.data_reg[57] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\mix1.data_reg[101] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\ks1.key_reg[57] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\mix1.data_reg[100] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\mix1.data_reg[103] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\mix1.data_reg[106] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\mix1.data_reg[86] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\mix1.data_reg[70] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\mix1.data_reg[123] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\mix1.data_reg[64] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\mix1.data_reg[112] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\mix1.data_reg[116] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\mix1.data_reg[113] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\ks1.key_reg[46] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\mix1.data_reg[83] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\mix1.data_reg[52] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\mix1.data_reg[107] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\mix1.data_reg[120] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\mix1.data_reg[90] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\mix1.data_reg[39] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\mix1.data_reg[43] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\mix1.data_reg[49] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\mix1.data_reg[122] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\mix1.data_reg[127] ),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(data_i[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(data_i[108]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(data_i[74]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 input101 (.A(data_i[75]),
    .X(net101));
 sky130_fd_sc_hd__buf_2 input102 (.A(data_i[76]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(data_i[77]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(data_i[78]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 input105 (.A(data_i[79]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(data_i[7]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(data_i[80]),
    .X(net107));
 sky130_fd_sc_hd__buf_1 input108 (.A(data_i[81]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(data_i[82]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(data_i[109]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(data_i[83]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(data_i[84]),
    .X(net111));
 sky130_fd_sc_hd__buf_1 input112 (.A(data_i[85]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(data_i[86]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(data_i[87]),
    .X(net114));
 sky130_fd_sc_hd__buf_2 input115 (.A(data_i[88]),
    .X(net115));
 sky130_fd_sc_hd__buf_1 input116 (.A(data_i[89]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(data_i[8]),
    .X(net117));
 sky130_fd_sc_hd__buf_4 input118 (.A(data_i[90]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(data_i[91]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(data_i[10]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(data_i[92]),
    .X(net120));
 sky130_fd_sc_hd__buf_1 input121 (.A(data_i[93]),
    .X(net121));
 sky130_fd_sc_hd__buf_2 input122 (.A(data_i[94]),
    .X(net122));
 sky130_fd_sc_hd__buf_1 input123 (.A(data_i[95]),
    .X(net123));
 sky130_fd_sc_hd__buf_1 input124 (.A(data_i[96]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_4 input125 (.A(data_i[97]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input126 (.A(data_i[98]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 input127 (.A(data_i[99]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 input128 (.A(data_i[9]),
    .X(net128));
 sky130_fd_sc_hd__buf_4 input129 (.A(decrypt_i),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(data_i[110]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input130 (.A(key_i[0]),
    .X(net130));
 sky130_fd_sc_hd__buf_4 input131 (.A(key_i[100]),
    .X(net131));
 sky130_fd_sc_hd__buf_1 input132 (.A(key_i[101]),
    .X(net132));
 sky130_fd_sc_hd__dlymetal6s2s_1 input133 (.A(key_i[102]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 input134 (.A(key_i[103]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 input135 (.A(key_i[104]),
    .X(net135));
 sky130_fd_sc_hd__buf_2 input136 (.A(key_i[105]),
    .X(net136));
 sky130_fd_sc_hd__dlymetal6s2s_1 input137 (.A(key_i[106]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 input138 (.A(key_i[107]),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(key_i[108]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input14 (.A(data_i[111]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input140 (.A(key_i[109]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_2 input141 (.A(key_i[10]),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input142 (.A(key_i[110]),
    .X(net142));
 sky130_fd_sc_hd__buf_2 input143 (.A(key_i[111]),
    .X(net143));
 sky130_fd_sc_hd__buf_2 input144 (.A(key_i[112]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(key_i[113]),
    .X(net145));
 sky130_fd_sc_hd__buf_2 input146 (.A(key_i[114]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(key_i[115]),
    .X(net147));
 sky130_fd_sc_hd__buf_2 input148 (.A(key_i[116]),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input149 (.A(key_i[117]),
    .X(net149));
 sky130_fd_sc_hd__buf_1 input15 (.A(data_i[112]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input150 (.A(key_i[118]),
    .X(net150));
 sky130_fd_sc_hd__dlymetal6s2s_1 input151 (.A(key_i[119]),
    .X(net151));
 sky130_fd_sc_hd__dlymetal6s2s_1 input152 (.A(key_i[11]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(key_i[120]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(key_i[121]),
    .X(net154));
 sky130_fd_sc_hd__buf_1 input155 (.A(key_i[122]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 input156 (.A(key_i[123]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(key_i[124]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 input158 (.A(key_i[125]),
    .X(net158));
 sky130_fd_sc_hd__buf_4 input159 (.A(key_i[126]),
    .X(net159));
 sky130_fd_sc_hd__buf_1 input16 (.A(data_i[113]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input160 (.A(key_i[127]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 input161 (.A(key_i[12]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 input162 (.A(key_i[13]),
    .X(net162));
 sky130_fd_sc_hd__buf_1 input163 (.A(key_i[14]),
    .X(net163));
 sky130_fd_sc_hd__buf_1 input164 (.A(key_i[15]),
    .X(net164));
 sky130_fd_sc_hd__buf_2 input165 (.A(key_i[16]),
    .X(net165));
 sky130_fd_sc_hd__buf_1 input166 (.A(key_i[17]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 input167 (.A(key_i[18]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 input168 (.A(key_i[19]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 input169 (.A(key_i[1]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(data_i[114]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input170 (.A(key_i[20]),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(key_i[21]),
    .X(net171));
 sky130_fd_sc_hd__buf_4 input172 (.A(key_i[22]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 input173 (.A(key_i[23]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 input174 (.A(key_i[24]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 input175 (.A(key_i[25]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_4 input176 (.A(key_i[26]),
    .X(net176));
 sky130_fd_sc_hd__buf_2 input177 (.A(key_i[27]),
    .X(net177));
 sky130_fd_sc_hd__buf_2 input178 (.A(key_i[28]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(key_i[29]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(data_i[115]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input180 (.A(key_i[2]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 input181 (.A(key_i[30]),
    .X(net181));
 sky130_fd_sc_hd__buf_1 input182 (.A(key_i[31]),
    .X(net182));
 sky130_fd_sc_hd__buf_1 input183 (.A(key_i[32]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 input184 (.A(key_i[33]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 input185 (.A(key_i[34]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 input186 (.A(key_i[35]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 input187 (.A(key_i[36]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 input188 (.A(key_i[37]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 input189 (.A(key_i[38]),
    .X(net189));
 sky130_fd_sc_hd__buf_4 input19 (.A(data_i[116]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input190 (.A(key_i[39]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 input191 (.A(key_i[3]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 input192 (.A(key_i[40]),
    .X(net192));
 sky130_fd_sc_hd__buf_2 input193 (.A(key_i[41]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 input194 (.A(key_i[42]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 input195 (.A(key_i[43]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 input196 (.A(key_i[44]),
    .X(net196));
 sky130_fd_sc_hd__buf_1 input197 (.A(key_i[45]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(key_i[46]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 input199 (.A(key_i[47]),
    .X(net199));
 sky130_fd_sc_hd__buf_1 input2 (.A(data_i[100]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(data_i[117]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input200 (.A(key_i[48]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 input201 (.A(key_i[49]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_4 input202 (.A(key_i[4]),
    .X(net202));
 sky130_fd_sc_hd__buf_1 input203 (.A(key_i[50]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_2 input204 (.A(key_i[51]),
    .X(net204));
 sky130_fd_sc_hd__buf_2 input205 (.A(key_i[52]),
    .X(net205));
 sky130_fd_sc_hd__buf_4 input206 (.A(key_i[53]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 input207 (.A(key_i[54]),
    .X(net207));
 sky130_fd_sc_hd__buf_2 input208 (.A(key_i[55]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 input209 (.A(key_i[56]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(data_i[118]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_4 input210 (.A(key_i[57]),
    .X(net210));
 sky130_fd_sc_hd__buf_2 input211 (.A(key_i[58]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 input212 (.A(key_i[59]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(key_i[5]),
    .X(net213));
 sky130_fd_sc_hd__buf_1 input214 (.A(key_i[60]),
    .X(net214));
 sky130_fd_sc_hd__buf_2 input215 (.A(key_i[61]),
    .X(net215));
 sky130_fd_sc_hd__dlymetal6s2s_1 input216 (.A(key_i[62]),
    .X(net216));
 sky130_fd_sc_hd__buf_2 input217 (.A(key_i[63]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 input218 (.A(key_i[64]),
    .X(net218));
 sky130_fd_sc_hd__buf_1 input219 (.A(key_i[65]),
    .X(net219));
 sky130_fd_sc_hd__buf_1 input22 (.A(data_i[119]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input220 (.A(key_i[66]),
    .X(net220));
 sky130_fd_sc_hd__dlymetal6s2s_1 input221 (.A(key_i[67]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 input222 (.A(key_i[68]),
    .X(net222));
 sky130_fd_sc_hd__buf_2 input223 (.A(key_i[69]),
    .X(net223));
 sky130_fd_sc_hd__buf_1 input224 (.A(key_i[6]),
    .X(net224));
 sky130_fd_sc_hd__buf_4 input225 (.A(key_i[70]),
    .X(net225));
 sky130_fd_sc_hd__dlymetal6s2s_1 input226 (.A(key_i[71]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 input227 (.A(key_i[72]),
    .X(net227));
 sky130_fd_sc_hd__dlymetal6s2s_1 input228 (.A(key_i[73]),
    .X(net228));
 sky130_fd_sc_hd__dlymetal6s2s_1 input229 (.A(key_i[74]),
    .X(net229));
 sky130_fd_sc_hd__buf_2 input23 (.A(data_i[11]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input230 (.A(key_i[75]),
    .X(net230));
 sky130_fd_sc_hd__buf_2 input231 (.A(key_i[76]),
    .X(net231));
 sky130_fd_sc_hd__dlymetal6s2s_1 input232 (.A(key_i[77]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_4 input233 (.A(key_i[78]),
    .X(net233));
 sky130_fd_sc_hd__buf_1 input234 (.A(key_i[79]),
    .X(net234));
 sky130_fd_sc_hd__buf_2 input235 (.A(key_i[7]),
    .X(net235));
 sky130_fd_sc_hd__buf_2 input236 (.A(key_i[80]),
    .X(net236));
 sky130_fd_sc_hd__buf_2 input237 (.A(key_i[81]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 input238 (.A(key_i[82]),
    .X(net238));
 sky130_fd_sc_hd__buf_4 input239 (.A(key_i[83]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(data_i[120]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input240 (.A(key_i[84]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 input241 (.A(key_i[85]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 input242 (.A(key_i[86]),
    .X(net242));
 sky130_fd_sc_hd__buf_2 input243 (.A(key_i[87]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 input244 (.A(key_i[88]),
    .X(net244));
 sky130_fd_sc_hd__buf_1 input245 (.A(key_i[89]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 input246 (.A(key_i[8]),
    .X(net246));
 sky130_fd_sc_hd__buf_2 input247 (.A(key_i[90]),
    .X(net247));
 sky130_fd_sc_hd__buf_2 input248 (.A(key_i[91]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 input249 (.A(key_i[92]),
    .X(net249));
 sky130_fd_sc_hd__buf_2 input25 (.A(data_i[121]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input250 (.A(key_i[93]),
    .X(net250));
 sky130_fd_sc_hd__buf_2 input251 (.A(key_i[94]),
    .X(net251));
 sky130_fd_sc_hd__buf_1 input252 (.A(key_i[95]),
    .X(net252));
 sky130_fd_sc_hd__buf_1 input253 (.A(key_i[96]),
    .X(net253));
 sky130_fd_sc_hd__buf_1 input254 (.A(key_i[97]),
    .X(net254));
 sky130_fd_sc_hd__buf_2 input255 (.A(key_i[98]),
    .X(net255));
 sky130_fd_sc_hd__buf_2 input256 (.A(key_i[99]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 input257 (.A(key_i[9]),
    .X(net257));
 sky130_fd_sc_hd__buf_2 input258 (.A(load_i),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 input259 (.A(reset),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(data_i[122]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(data_i[123]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 input28 (.A(data_i[124]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(data_i[125]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(data_i[101]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input30 (.A(data_i[126]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(data_i[127]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(data_i[12]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(data_i[13]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(data_i[14]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(data_i[15]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(data_i[16]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input37 (.A(data_i[17]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(data_i[18]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(data_i[19]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input4 (.A(data_i[102]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(data_i[1]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(data_i[20]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 input42 (.A(data_i[21]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(data_i[22]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(data_i[23]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(data_i[24]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(data_i[25]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input47 (.A(data_i[26]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(data_i[27]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(data_i[28]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 input5 (.A(data_i[103]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input50 (.A(data_i[29]),
    .X(net50));
 sky130_fd_sc_hd__buf_4 input51 (.A(data_i[2]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(data_i[30]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(data_i[31]),
    .X(net53));
 sky130_fd_sc_hd__buf_2 input54 (.A(data_i[32]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(data_i[33]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(data_i[34]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(data_i[35]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(data_i[36]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_4 input59 (.A(data_i[37]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(data_i[104]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input60 (.A(data_i[38]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 input61 (.A(data_i[39]),
    .X(net61));
 sky130_fd_sc_hd__buf_2 input62 (.A(data_i[3]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(data_i[40]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(data_i[41]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(data_i[42]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(data_i[43]),
    .X(net66));
 sky130_fd_sc_hd__buf_2 input67 (.A(data_i[44]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(data_i[45]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(data_i[46]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(data_i[105]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(data_i[47]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(data_i[48]),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 input72 (.A(data_i[49]),
    .X(net72));
 sky130_fd_sc_hd__buf_2 input73 (.A(data_i[4]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(data_i[50]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(data_i[51]),
    .X(net75));
 sky130_fd_sc_hd__dlymetal6s2s_1 input76 (.A(data_i[52]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(data_i[53]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(data_i[54]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(data_i[55]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input8 (.A(data_i[106]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(data_i[56]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 input81 (.A(data_i[57]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(data_i[58]),
    .X(net82));
 sky130_fd_sc_hd__buf_2 input83 (.A(data_i[59]),
    .X(net83));
 sky130_fd_sc_hd__dlymetal6s2s_1 input84 (.A(data_i[5]),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input85 (.A(data_i[60]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(data_i[61]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 input87 (.A(data_i[62]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(data_i[63]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(data_i[64]),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input9 (.A(data_i[107]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(data_i[65]),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(data_i[66]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(data_i[67]),
    .X(net92));
 sky130_fd_sc_hd__buf_2 input93 (.A(data_i[68]),
    .X(net93));
 sky130_fd_sc_hd__dlymetal6s2s_1 input94 (.A(data_i[69]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(data_i[6]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(data_i[70]),
    .X(net96));
 sky130_fd_sc_hd__buf_2 input97 (.A(data_i[71]),
    .X(net97));
 sky130_fd_sc_hd__buf_2 input98 (.A(data_i[72]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input99 (.A(data_i[73]),
    .X(net99));
 sky130_fd_sc_hd__buf_4 max_cap389 (.A(_0750_),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net260),
    .X(data_o[0]));
 sky130_fd_sc_hd__clkbuf_4 output261 (.A(net261),
    .X(data_o[100]));
 sky130_fd_sc_hd__clkbuf_4 output262 (.A(net262),
    .X(data_o[101]));
 sky130_fd_sc_hd__clkbuf_4 output263 (.A(net263),
    .X(data_o[102]));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net264),
    .X(data_o[103]));
 sky130_fd_sc_hd__clkbuf_4 output265 (.A(net265),
    .X(data_o[104]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(data_o[105]));
 sky130_fd_sc_hd__clkbuf_4 output267 (.A(net267),
    .X(data_o[106]));
 sky130_fd_sc_hd__clkbuf_4 output268 (.A(net268),
    .X(data_o[107]));
 sky130_fd_sc_hd__clkbuf_4 output269 (.A(net269),
    .X(data_o[108]));
 sky130_fd_sc_hd__clkbuf_4 output270 (.A(net270),
    .X(data_o[109]));
 sky130_fd_sc_hd__clkbuf_4 output271 (.A(net271),
    .X(data_o[10]));
 sky130_fd_sc_hd__clkbuf_4 output272 (.A(net272),
    .X(data_o[110]));
 sky130_fd_sc_hd__clkbuf_4 output273 (.A(net273),
    .X(data_o[111]));
 sky130_fd_sc_hd__clkbuf_4 output274 (.A(net274),
    .X(data_o[112]));
 sky130_fd_sc_hd__clkbuf_4 output275 (.A(net275),
    .X(data_o[113]));
 sky130_fd_sc_hd__clkbuf_4 output276 (.A(net276),
    .X(data_o[114]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(data_o[115]));
 sky130_fd_sc_hd__clkbuf_4 output278 (.A(net278),
    .X(data_o[116]));
 sky130_fd_sc_hd__clkbuf_4 output279 (.A(net279),
    .X(data_o[117]));
 sky130_fd_sc_hd__clkbuf_4 output280 (.A(net280),
    .X(data_o[118]));
 sky130_fd_sc_hd__clkbuf_4 output281 (.A(net281),
    .X(data_o[119]));
 sky130_fd_sc_hd__clkbuf_4 output282 (.A(net282),
    .X(data_o[11]));
 sky130_fd_sc_hd__clkbuf_4 output283 (.A(net283),
    .X(data_o[120]));
 sky130_fd_sc_hd__clkbuf_4 output284 (.A(net284),
    .X(data_o[121]));
 sky130_fd_sc_hd__clkbuf_4 output285 (.A(net285),
    .X(data_o[122]));
 sky130_fd_sc_hd__clkbuf_4 output286 (.A(net286),
    .X(data_o[123]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(data_o[124]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(data_o[125]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(data_o[126]));
 sky130_fd_sc_hd__clkbuf_4 output290 (.A(net290),
    .X(data_o[127]));
 sky130_fd_sc_hd__clkbuf_4 output291 (.A(net291),
    .X(data_o[12]));
 sky130_fd_sc_hd__clkbuf_4 output292 (.A(net292),
    .X(data_o[13]));
 sky130_fd_sc_hd__clkbuf_4 output293 (.A(net293),
    .X(data_o[14]));
 sky130_fd_sc_hd__clkbuf_4 output294 (.A(net294),
    .X(data_o[15]));
 sky130_fd_sc_hd__clkbuf_4 output295 (.A(net295),
    .X(data_o[16]));
 sky130_fd_sc_hd__clkbuf_4 output296 (.A(net296),
    .X(data_o[17]));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(data_o[18]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(data_o[19]));
 sky130_fd_sc_hd__clkbuf_4 output299 (.A(net299),
    .X(data_o[1]));
 sky130_fd_sc_hd__clkbuf_4 output300 (.A(net300),
    .X(data_o[20]));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(data_o[21]));
 sky130_fd_sc_hd__clkbuf_4 output302 (.A(net302),
    .X(data_o[22]));
 sky130_fd_sc_hd__clkbuf_4 output303 (.A(net303),
    .X(data_o[23]));
 sky130_fd_sc_hd__clkbuf_4 output304 (.A(net304),
    .X(data_o[24]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(data_o[25]));
 sky130_fd_sc_hd__clkbuf_4 output306 (.A(net306),
    .X(data_o[26]));
 sky130_fd_sc_hd__clkbuf_4 output307 (.A(net307),
    .X(data_o[27]));
 sky130_fd_sc_hd__clkbuf_4 output308 (.A(net308),
    .X(data_o[28]));
 sky130_fd_sc_hd__clkbuf_4 output309 (.A(net309),
    .X(data_o[29]));
 sky130_fd_sc_hd__clkbuf_4 output310 (.A(net310),
    .X(data_o[2]));
 sky130_fd_sc_hd__clkbuf_4 output311 (.A(net311),
    .X(data_o[30]));
 sky130_fd_sc_hd__clkbuf_4 output312 (.A(net312),
    .X(data_o[31]));
 sky130_fd_sc_hd__clkbuf_4 output313 (.A(net313),
    .X(data_o[32]));
 sky130_fd_sc_hd__clkbuf_4 output314 (.A(net314),
    .X(data_o[33]));
 sky130_fd_sc_hd__clkbuf_4 output315 (.A(net315),
    .X(data_o[34]));
 sky130_fd_sc_hd__clkbuf_4 output316 (.A(net316),
    .X(data_o[35]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .X(data_o[36]));
 sky130_fd_sc_hd__clkbuf_4 output318 (.A(net318),
    .X(data_o[37]));
 sky130_fd_sc_hd__clkbuf_4 output319 (.A(net319),
    .X(data_o[38]));
 sky130_fd_sc_hd__clkbuf_4 output320 (.A(net320),
    .X(data_o[39]));
 sky130_fd_sc_hd__clkbuf_4 output321 (.A(net321),
    .X(data_o[3]));
 sky130_fd_sc_hd__clkbuf_4 output322 (.A(net322),
    .X(data_o[40]));
 sky130_fd_sc_hd__clkbuf_4 output323 (.A(net323),
    .X(data_o[41]));
 sky130_fd_sc_hd__clkbuf_4 output324 (.A(net324),
    .X(data_o[42]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(data_o[43]));
 sky130_fd_sc_hd__clkbuf_4 output326 (.A(net326),
    .X(data_o[44]));
 sky130_fd_sc_hd__clkbuf_4 output327 (.A(net327),
    .X(data_o[45]));
 sky130_fd_sc_hd__clkbuf_4 output328 (.A(net328),
    .X(data_o[46]));
 sky130_fd_sc_hd__clkbuf_4 output329 (.A(net329),
    .X(data_o[47]));
 sky130_fd_sc_hd__clkbuf_4 output330 (.A(net330),
    .X(data_o[48]));
 sky130_fd_sc_hd__clkbuf_4 output331 (.A(net331),
    .X(data_o[49]));
 sky130_fd_sc_hd__clkbuf_4 output332 (.A(net332),
    .X(data_o[4]));
 sky130_fd_sc_hd__clkbuf_4 output333 (.A(net333),
    .X(data_o[50]));
 sky130_fd_sc_hd__clkbuf_4 output334 (.A(net334),
    .X(data_o[51]));
 sky130_fd_sc_hd__clkbuf_4 output335 (.A(net335),
    .X(data_o[52]));
 sky130_fd_sc_hd__clkbuf_4 output336 (.A(net336),
    .X(data_o[53]));
 sky130_fd_sc_hd__clkbuf_4 output337 (.A(net337),
    .X(data_o[54]));
 sky130_fd_sc_hd__clkbuf_4 output338 (.A(net338),
    .X(data_o[55]));
 sky130_fd_sc_hd__clkbuf_4 output339 (.A(net339),
    .X(data_o[56]));
 sky130_fd_sc_hd__clkbuf_4 output340 (.A(net340),
    .X(data_o[57]));
 sky130_fd_sc_hd__clkbuf_4 output341 (.A(net341),
    .X(data_o[58]));
 sky130_fd_sc_hd__clkbuf_4 output342 (.A(net342),
    .X(data_o[59]));
 sky130_fd_sc_hd__clkbuf_4 output343 (.A(net343),
    .X(data_o[5]));
 sky130_fd_sc_hd__clkbuf_4 output344 (.A(net344),
    .X(data_o[60]));
 sky130_fd_sc_hd__clkbuf_4 output345 (.A(net345),
    .X(data_o[61]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(data_o[62]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .X(data_o[63]));
 sky130_fd_sc_hd__clkbuf_4 output348 (.A(net348),
    .X(data_o[64]));
 sky130_fd_sc_hd__clkbuf_4 output349 (.A(net349),
    .X(data_o[65]));
 sky130_fd_sc_hd__clkbuf_4 output350 (.A(net350),
    .X(data_o[66]));
 sky130_fd_sc_hd__clkbuf_4 output351 (.A(net351),
    .X(data_o[67]));
 sky130_fd_sc_hd__clkbuf_4 output352 (.A(net352),
    .X(data_o[68]));
 sky130_fd_sc_hd__clkbuf_4 output353 (.A(net353),
    .X(data_o[69]));
 sky130_fd_sc_hd__clkbuf_4 output354 (.A(net354),
    .X(data_o[6]));
 sky130_fd_sc_hd__clkbuf_4 output355 (.A(net355),
    .X(data_o[70]));
 sky130_fd_sc_hd__clkbuf_4 output356 (.A(net356),
    .X(data_o[71]));
 sky130_fd_sc_hd__clkbuf_4 output357 (.A(net357),
    .X(data_o[72]));
 sky130_fd_sc_hd__clkbuf_4 output358 (.A(net358),
    .X(data_o[73]));
 sky130_fd_sc_hd__clkbuf_4 output359 (.A(net359),
    .X(data_o[74]));
 sky130_fd_sc_hd__clkbuf_4 output360 (.A(net360),
    .X(data_o[75]));
 sky130_fd_sc_hd__clkbuf_4 output361 (.A(net361),
    .X(data_o[76]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(data_o[77]));
 sky130_fd_sc_hd__clkbuf_4 output363 (.A(net363),
    .X(data_o[78]));
 sky130_fd_sc_hd__clkbuf_4 output364 (.A(net364),
    .X(data_o[79]));
 sky130_fd_sc_hd__clkbuf_4 output365 (.A(net365),
    .X(data_o[7]));
 sky130_fd_sc_hd__clkbuf_4 output366 (.A(net366),
    .X(data_o[80]));
 sky130_fd_sc_hd__buf_2 output367 (.A(net367),
    .X(data_o[81]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .X(data_o[82]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(data_o[83]));
 sky130_fd_sc_hd__clkbuf_4 output370 (.A(net370),
    .X(data_o[84]));
 sky130_fd_sc_hd__clkbuf_4 output371 (.A(net371),
    .X(data_o[85]));
 sky130_fd_sc_hd__clkbuf_4 output372 (.A(net372),
    .X(data_o[86]));
 sky130_fd_sc_hd__clkbuf_4 output373 (.A(net373),
    .X(data_o[87]));
 sky130_fd_sc_hd__clkbuf_4 output374 (.A(net374),
    .X(data_o[88]));
 sky130_fd_sc_hd__clkbuf_4 output375 (.A(net375),
    .X(data_o[89]));
 sky130_fd_sc_hd__clkbuf_4 output376 (.A(net376),
    .X(data_o[8]));
 sky130_fd_sc_hd__clkbuf_4 output377 (.A(net377),
    .X(data_o[90]));
 sky130_fd_sc_hd__clkbuf_4 output378 (.A(net378),
    .X(data_o[91]));
 sky130_fd_sc_hd__clkbuf_4 output379 (.A(net379),
    .X(data_o[92]));
 sky130_fd_sc_hd__clkbuf_4 output380 (.A(net380),
    .X(data_o[93]));
 sky130_fd_sc_hd__clkbuf_4 output381 (.A(net381),
    .X(data_o[94]));
 sky130_fd_sc_hd__clkbuf_4 output382 (.A(net382),
    .X(data_o[95]));
 sky130_fd_sc_hd__clkbuf_4 output383 (.A(net383),
    .X(data_o[96]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .X(data_o[97]));
 sky130_fd_sc_hd__clkbuf_4 output385 (.A(net385),
    .X(data_o[98]));
 sky130_fd_sc_hd__clkbuf_4 output386 (.A(net386),
    .X(data_o[99]));
 sky130_fd_sc_hd__clkbuf_4 output387 (.A(net387),
    .X(data_o[9]));
 sky130_fd_sc_hd__clkbuf_4 output388 (.A(net388),
    .X(ready_o));
endmodule

