VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO aes_Trojan
  CLASS BLOCK ;
  FOREIGN aes_Trojan ;
  ORIGIN 0.000 0.000 ;
  SIZE 650.000 BY 650.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END clk
  PIN data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 646.000 61.550 650.000 ;
    END
  END data_i[0]
  PIN data_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 325.310 646.000 325.590 650.000 ;
    END
  END data_i[100]
  PIN data_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END data_i[101]
  PIN data_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END data_i[102]
  PIN data_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END data_i[103]
  PIN data_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 197.240 650.000 197.840 ;
    END
  END data_i[104]
  PIN data_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END data_i[105]
  PIN data_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END data_i[106]
  PIN data_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END data_i[107]
  PIN data_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END data_i[108]
  PIN data_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 336.640 650.000 337.240 ;
    END
  END data_i[109]
  PIN data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 513.440 650.000 514.040 ;
    END
  END data_i[10]
  PIN data_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 74.840 650.000 75.440 ;
    END
  END data_i[110]
  PIN data_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END data_i[111]
  PIN data_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 646.000 22.910 650.000 ;
    END
  END data_i[112]
  PIN data_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END data_i[113]
  PIN data_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END data_i[114]
  PIN data_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 560.370 646.000 560.650 650.000 ;
    END
  END data_i[115]
  PIN data_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END data_i[116]
  PIN data_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 343.440 650.000 344.040 ;
    END
  END data_i[117]
  PIN data_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 646.000 13.250 650.000 ;
    END
  END data_i[118]
  PIN data_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 293.110 646.000 293.390 650.000 ;
    END
  END data_i[119]
  PIN data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 622.240 650.000 622.840 ;
    END
  END data_i[11]
  PIN data_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END data_i[120]
  PIN data_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 412.250 646.000 412.530 650.000 ;
    END
  END data_i[121]
  PIN data_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END data_i[122]
  PIN data_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 142.840 650.000 143.440 ;
    END
  END data_i[123]
  PIN data_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 386.490 646.000 386.770 650.000 ;
    END
  END data_i[124]
  PIN data_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END data_i[125]
  PIN data_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END data_i[126]
  PIN data_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END data_i[127]
  PIN data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 646.000 6.810 650.000 ;
    END
  END data_i[12]
  PIN data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 495.970 646.000 496.250 650.000 ;
    END
  END data_i[13]
  PIN data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 360.730 646.000 361.010 650.000 ;
    END
  END data_i[14]
  PIN data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END data_i[15]
  PIN data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END data_i[16]
  PIN data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END data_i[17]
  PIN data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 254.470 646.000 254.750 650.000 ;
    END
  END data_i[18]
  PIN data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END data_i[19]
  PIN data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 646.000 286.950 650.000 ;
    END
  END data_i[1]
  PIN data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END data_i[20]
  PIN data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 646.000 35.790 650.000 ;
    END
  END data_i[21]
  PIN data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 499.840 650.000 500.440 ;
    END
  END data_i[22]
  PIN data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END data_i[23]
  PIN data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 235.150 646.000 235.430 650.000 ;
    END
  END data_i[24]
  PIN data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 579.690 646.000 579.970 650.000 ;
    END
  END data_i[25]
  PIN data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END data_i[26]
  PIN data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 515.290 646.000 515.570 650.000 ;
    END
  END data_i[27]
  PIN data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 404.640 650.000 405.240 ;
    END
  END data_i[28]
  PIN data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 431.840 650.000 432.440 ;
    END
  END data_i[29]
  PIN data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 581.440 650.000 582.040 ;
    END
  END data_i[2]
  PIN data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END data_i[30]
  PIN data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END data_i[31]
  PIN data_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END data_i[32]
  PIN data_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END data_i[33]
  PIN data_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 646.000 100.190 650.000 ;
    END
  END data_i[34]
  PIN data_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 646.000 164.590 650.000 ;
    END
  END data_i[35]
  PIN data_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 312.430 646.000 312.710 650.000 ;
    END
  END data_i[36]
  PIN data_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END data_i[37]
  PIN data_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 534.610 646.000 534.890 650.000 ;
    END
  END data_i[38]
  PIN data_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END data_i[39]
  PIN data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 156.440 650.000 157.040 ;
    END
  END data_i[3]
  PIN data_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 483.090 646.000 483.370 650.000 ;
    END
  END data_i[40]
  PIN data_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END data_i[41]
  PIN data_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 102.040 650.000 102.640 ;
    END
  END data_i[42]
  PIN data_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END data_i[43]
  PIN data_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END data_i[44]
  PIN data_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 644.090 646.000 644.370 650.000 ;
    END
  END data_i[45]
  PIN data_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END data_i[46]
  PIN data_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END data_i[47]
  PIN data_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 646.000 228.990 650.000 ;
    END
  END data_i[48]
  PIN data_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 646.000 393.210 650.000 ;
    END
  END data_i[49]
  PIN data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 61.240 650.000 61.840 ;
    END
  END data_i[4]
  PIN data_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END data_i[50]
  PIN data_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END data_i[51]
  PIN data_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END data_i[52]
  PIN data_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 566.810 646.000 567.090 650.000 ;
    END
  END data_i[53]
  PIN data_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END data_i[54]
  PIN data_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 642.640 650.000 643.240 ;
    END
  END data_i[55]
  PIN data_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END data_i[56]
  PIN data_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 248.030 646.000 248.310 650.000 ;
    END
  END data_i[57]
  PIN data_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 224.440 650.000 225.040 ;
    END
  END data_i[58]
  PIN data_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 533.840 650.000 534.440 ;
    END
  END data_i[59]
  PIN data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 646.000 145.270 650.000 ;
    END
  END data_i[5]
  PIN data_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 574.640 650.000 575.240 ;
    END
  END data_i[60]
  PIN data_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END data_i[61]
  PIN data_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END data_i[62]
  PIN data_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 329.840 650.000 330.440 ;
    END
  END data_i[63]
  PIN data_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END data_i[64]
  PIN data_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 115.640 650.000 116.240 ;
    END
  END data_i[65]
  PIN data_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 646.000 48.670 650.000 ;
    END
  END data_i[66]
  PIN data_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 646.000 299.830 650.000 ;
    END
  END data_i[67]
  PIN data_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END data_i[68]
  PIN data_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 238.040 650.000 238.640 ;
    END
  END data_i[69]
  PIN data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 646.000 380.330 650.000 ;
    END
  END data_i[6]
  PIN data_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 399.370 646.000 399.650 650.000 ;
    END
  END data_i[70]
  PIN data_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 40.840 650.000 41.440 ;
    END
  END data_i[71]
  PIN data_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 334.970 646.000 335.250 650.000 ;
    END
  END data_i[72]
  PIN data_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END data_i[73]
  PIN data_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 384.240 650.000 384.840 ;
    END
  END data_i[74]
  PIN data_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 646.000 138.830 650.000 ;
    END
  END data_i[75]
  PIN data_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END data_i[76]
  PIN data_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END data_i[77]
  PIN data_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END data_i[78]
  PIN data_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 222.270 646.000 222.550 650.000 ;
    END
  END data_i[79]
  PIN data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 68.040 650.000 68.640 ;
    END
  END data_i[7]
  PIN data_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 452.240 650.000 452.840 ;
    END
  END data_i[80]
  PIN data_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 646.000 171.030 650.000 ;
    END
  END data_i[81]
  PIN data_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END data_i[82]
  PIN data_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 527.040 650.000 527.640 ;
    END
  END data_i[83]
  PIN data_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END data_i[84]
  PIN data_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END data_i[85]
  PIN data_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 299.240 650.000 299.840 ;
    END
  END data_i[86]
  PIN data_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END data_i[87]
  PIN data_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END data_i[88]
  PIN data_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END data_i[89]
  PIN data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 540.640 650.000 541.240 ;
    END
  END data_i[8]
  PIN data_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 444.450 646.000 444.730 650.000 ;
    END
  END data_i[90]
  PIN data_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 615.440 650.000 616.040 ;
    END
  END data_i[91]
  PIN data_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 95.240 650.000 95.840 ;
    END
  END data_i[92]
  PIN data_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END data_i[93]
  PIN data_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 646.000 80.870 650.000 ;
    END
  END data_i[94]
  PIN data_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END data_i[95]
  PIN data_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 646.000 55.110 650.000 ;
    END
  END data_i[96]
  PIN data_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END data_i[97]
  PIN data_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 67.710 646.000 67.990 650.000 ;
    END
  END data_i[98]
  PIN data_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END data_i[99]
  PIN data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 646.000 132.390 650.000 ;
    END
  END data_i[9]
  PIN data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END data_o[0]
  PIN data_o[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END data_o[100]
  PIN data_o[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END data_o[101]
  PIN data_o[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END data_o[102]
  PIN data_o[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END data_o[103]
  PIN data_o[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 459.040 650.000 459.640 ;
    END
  END data_o[104]
  PIN data_o[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 418.240 650.000 418.840 ;
    END
  END data_o[105]
  PIN data_o[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END data_o[106]
  PIN data_o[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END data_o[107]
  PIN data_o[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END data_o[108]
  PIN data_o[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 646.000 113.070 650.000 ;
    END
  END data_o[109]
  PIN data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END data_o[10]
  PIN data_o[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 608.640 650.000 609.240 ;
    END
  END data_o[110]
  PIN data_o[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END data_o[111]
  PIN data_o[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 204.040 650.000 204.640 ;
    END
  END data_o[112]
  PIN data_o[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END data_o[113]
  PIN data_o[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END data_o[114]
  PIN data_o[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 486.240 650.000 486.840 ;
    END
  END data_o[115]
  PIN data_o[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 151.430 646.000 151.710 650.000 ;
    END
  END data_o[116]
  PIN data_o[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 136.040 650.000 136.640 ;
    END
  END data_o[117]
  PIN data_o[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END data_o[118]
  PIN data_o[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END data_o[119]
  PIN data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 231.240 650.000 231.840 ;
    END
  END data_o[11]
  PIN data_o[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END data_o[120]
  PIN data_o[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END data_o[121]
  PIN data_o[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END data_o[122]
  PIN data_o[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END data_o[123]
  PIN data_o[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 554.240 650.000 554.840 ;
    END
  END data_o[124]
  PIN data_o[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 520.240 650.000 520.840 ;
    END
  END data_o[125]
  PIN data_o[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 258.440 650.000 259.040 ;
    END
  END data_o[126]
  PIN data_o[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END data_o[127]
  PIN data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END data_o[12]
  PIN data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 605.450 646.000 605.730 650.000 ;
    END
  END data_o[13]
  PIN data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 210.840 650.000 211.440 ;
    END
  END data_o[14]
  PIN data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 637.650 646.000 637.930 650.000 ;
    END
  END data_o[15]
  PIN data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 646.000 0.370 650.000 ;
    END
  END data_o[16]
  PIN data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END data_o[17]
  PIN data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 418.690 646.000 418.970 650.000 ;
    END
  END data_o[18]
  PIN data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 108.840 650.000 109.440 ;
    END
  END data_o[19]
  PIN data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 347.850 646.000 348.130 650.000 ;
    END
  END data_o[1]
  PIN data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END data_o[20]
  PIN data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END data_o[21]
  PIN data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 425.040 650.000 425.640 ;
    END
  END data_o[22]
  PIN data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END data_o[23]
  PIN data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END data_o[24]
  PIN data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 217.640 650.000 218.240 ;
    END
  END data_o[25]
  PIN data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END data_o[26]
  PIN data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 318.870 646.000 319.150 650.000 ;
    END
  END data_o[27]
  PIN data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 646.000 47.640 650.000 48.240 ;
    END
  END data_o[28]
  PIN data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END data_o[29]
  PIN data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END data_o[2]
  PIN data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 438.640 650.000 439.240 ;
    END
  END data_o[30]
  PIN data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 176.840 650.000 177.440 ;
    END
  END data_o[31]
  PIN data_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END data_o[32]
  PIN data_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 20.440 650.000 21.040 ;
    END
  END data_o[33]
  PIN data_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END data_o[34]
  PIN data_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.870 646.000 158.150 650.000 ;
    END
  END data_o[35]
  PIN data_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 646.000 129.240 650.000 129.840 ;
    END
  END data_o[36]
  PIN data_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.950 646.000 42.230 650.000 ;
    END
  END data_o[37]
  PIN data_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END data_o[38]
  PIN data_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END data_o[39]
  PIN data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END data_o[3]
  PIN data_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END data_o[40]
  PIN data_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END data_o[41]
  PIN data_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END data_o[42]
  PIN data_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 405.810 646.000 406.090 650.000 ;
    END
  END data_o[43]
  PIN data_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END data_o[44]
  PIN data_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END data_o[45]
  PIN data_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END data_o[46]
  PIN data_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END data_o[47]
  PIN data_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END data_o[48]
  PIN data_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 202.950 646.000 203.230 650.000 ;
    END
  END data_o[49]
  PIN data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END data_o[4]
  PIN data_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 646.000 88.440 650.000 89.040 ;
    END
  END data_o[50]
  PIN data_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 573.250 646.000 573.530 650.000 ;
    END
  END data_o[51]
  PIN data_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END data_o[52]
  PIN data_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 367.170 646.000 367.450 650.000 ;
    END
  END data_o[53]
  PIN data_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END data_o[54]
  PIN data_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 599.010 646.000 599.290 650.000 ;
    END
  END data_o[55]
  PIN data_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 119.230 646.000 119.510 650.000 ;
    END
  END data_o[56]
  PIN data_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END data_o[57]
  PIN data_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END data_o[58]
  PIN data_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END data_o[59]
  PIN data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 373.610 646.000 373.890 650.000 ;
    END
  END data_o[5]
  PIN data_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END data_o[60]
  PIN data_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 251.640 650.000 252.240 ;
    END
  END data_o[61]
  PIN data_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 183.640 650.000 184.240 ;
    END
  END data_o[62]
  PIN data_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 397.840 650.000 398.440 ;
    END
  END data_o[63]
  PIN data_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END data_o[64]
  PIN data_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 106.350 646.000 106.630 650.000 ;
    END
  END data_o[65]
  PIN data_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 646.000 323.040 650.000 323.640 ;
    END
  END data_o[66]
  PIN data_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END data_o[67]
  PIN data_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END data_o[68]
  PIN data_o[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END data_o[69]
  PIN data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END data_o[6]
  PIN data_o[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END data_o[70]
  PIN data_o[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 646.000 6.840 650.000 7.440 ;
    END
  END data_o[71]
  PIN data_o[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 278.840 650.000 279.440 ;
    END
  END data_o[72]
  PIN data_o[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 635.840 650.000 636.440 ;
    END
  END data_o[73]
  PIN data_o[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END data_o[74]
  PIN data_o[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 547.490 646.000 547.770 650.000 ;
    END
  END data_o[75]
  PIN data_o[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END data_o[76]
  PIN data_o[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 646.000 350.240 650.000 350.840 ;
    END
  END data_o[77]
  PIN data_o[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END data_o[78]
  PIN data_o[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 508.850 646.000 509.130 650.000 ;
    END
  END data_o[79]
  PIN data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END data_o[7]
  PIN data_o[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 190.070 646.000 190.350 650.000 ;
    END
  END data_o[80]
  PIN data_o[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 561.040 650.000 561.640 ;
    END
  END data_o[81]
  PIN data_o[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 601.840 650.000 602.440 ;
    END
  END data_o[82]
  PIN data_o[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 506.640 650.000 507.240 ;
    END
  END data_o[83]
  PIN data_o[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END data_o[84]
  PIN data_o[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 479.440 650.000 480.040 ;
    END
  END data_o[85]
  PIN data_o[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END data_o[86]
  PIN data_o[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END data_o[87]
  PIN data_o[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 280.230 646.000 280.510 650.000 ;
    END
  END data_o[88]
  PIN data_o[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END data_o[89]
  PIN data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END data_o[8]
  PIN data_o[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END data_o[90]
  PIN data_o[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END data_o[91]
  PIN data_o[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 629.040 650.000 629.640 ;
    END
  END data_o[92]
  PIN data_o[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 646.000 34.040 650.000 34.640 ;
    END
  END data_o[93]
  PIN data_o[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 305.990 646.000 306.270 650.000 ;
    END
  END data_o[94]
  PIN data_o[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END data_o[95]
  PIN data_o[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END data_o[96]
  PIN data_o[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END data_o[97]
  PIN data_o[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 586.130 646.000 586.410 650.000 ;
    END
  END data_o[98]
  PIN data_o[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END data_o[99]
  PIN data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END data_o[9]
  PIN decrypt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END decrypt_i
  PIN key_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 272.040 650.000 272.640 ;
    END
  END key_i[0]
  PIN key_i[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END key_i[100]
  PIN key_i[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END key_i[101]
  PIN key_i[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 273.790 646.000 274.070 650.000 ;
    END
  END key_i[102]
  PIN key_i[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END key_i[103]
  PIN key_i[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END key_i[104]
  PIN key_i[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 489.530 646.000 489.810 650.000 ;
    END
  END key_i[105]
  PIN key_i[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 292.440 650.000 293.040 ;
    END
  END key_i[106]
  PIN key_i[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END key_i[107]
  PIN key_i[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 611.890 646.000 612.170 650.000 ;
    END
  END key_i[108]
  PIN key_i[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 27.240 650.000 27.840 ;
    END
  END key_i[109]
  PIN key_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 431.570 646.000 431.850 650.000 ;
    END
  END key_i[10]
  PIN key_i[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END key_i[110]
  PIN key_i[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END key_i[111]
  PIN key_i[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END key_i[112]
  PIN key_i[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 285.640 650.000 286.240 ;
    END
  END key_i[113]
  PIN key_i[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 646.000 29.350 650.000 ;
    END
  END key_i[114]
  PIN key_i[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 391.040 650.000 391.640 ;
    END
  END key_i[115]
  PIN key_i[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END key_i[116]
  PIN key_i[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END key_i[117]
  PIN key_i[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END key_i[118]
  PIN key_i[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 592.570 646.000 592.850 650.000 ;
    END
  END key_i[119]
  PIN key_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 465.840 650.000 466.440 ;
    END
  END key_i[11]
  PIN key_i[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 646.000 216.110 650.000 ;
    END
  END key_i[120]
  PIN key_i[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 267.350 646.000 267.630 650.000 ;
    END
  END key_i[121]
  PIN key_i[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 81.640 650.000 82.240 ;
    END
  END key_i[122]
  PIN key_i[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 646.000 177.470 650.000 ;
    END
  END key_i[123]
  PIN key_i[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END key_i[124]
  PIN key_i[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 470.210 646.000 470.490 650.000 ;
    END
  END key_i[125]
  PIN key_i[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 341.410 646.000 341.690 650.000 ;
    END
  END key_i[126]
  PIN key_i[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 646.000 93.750 650.000 ;
    END
  END key_i[127]
  PIN key_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END key_i[12]
  PIN key_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END key_i[13]
  PIN key_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 445.440 650.000 446.040 ;
    END
  END key_i[14]
  PIN key_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 411.440 650.000 412.040 ;
    END
  END key_i[15]
  PIN key_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END key_i[16]
  PIN key_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 363.840 650.000 364.440 ;
    END
  END key_i[17]
  PIN key_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END key_i[18]
  PIN key_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END key_i[19]
  PIN key_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 450.890 646.000 451.170 650.000 ;
    END
  END key_i[1]
  PIN key_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 624.770 646.000 625.050 650.000 ;
    END
  END key_i[20]
  PIN key_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END key_i[21]
  PIN key_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END key_i[22]
  PIN key_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 122.440 650.000 123.040 ;
    END
  END key_i[23]
  PIN key_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 646.000 125.950 650.000 ;
    END
  END key_i[24]
  PIN key_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END key_i[25]
  PIN key_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END key_i[26]
  PIN key_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 260.910 646.000 261.190 650.000 ;
    END
  END key_i[27]
  PIN key_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END key_i[28]
  PIN key_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 595.040 650.000 595.640 ;
    END
  END key_i[29]
  PIN key_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END key_i[2]
  PIN key_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 541.050 646.000 541.330 650.000 ;
    END
  END key_i[30]
  PIN key_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 244.840 650.000 245.440 ;
    END
  END key_i[31]
  PIN key_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END key_i[32]
  PIN key_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 521.730 646.000 522.010 650.000 ;
    END
  END key_i[33]
  PIN key_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END key_i[34]
  PIN key_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END key_i[35]
  PIN key_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END key_i[36]
  PIN key_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END key_i[37]
  PIN key_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 149.640 650.000 150.240 ;
    END
  END key_i[38]
  PIN key_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 241.590 646.000 241.870 650.000 ;
    END
  END key_i[39]
  PIN key_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 547.440 650.000 548.040 ;
    END
  END key_i[3]
  PIN key_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END key_i[40]
  PIN key_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END key_i[41]
  PIN key_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END key_i[42]
  PIN key_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END key_i[43]
  PIN key_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END key_i[44]
  PIN key_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 316.240 650.000 316.840 ;
    END
  END key_i[45]
  PIN key_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END key_i[46]
  PIN key_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 463.770 646.000 464.050 650.000 ;
    END
  END key_i[47]
  PIN key_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 618.330 646.000 618.610 650.000 ;
    END
  END key_i[48]
  PIN key_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 74.150 646.000 74.430 650.000 ;
    END
  END key_i[49]
  PIN key_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END key_i[4]
  PIN key_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 370.640 650.000 371.240 ;
    END
  END key_i[50]
  PIN key_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 631.210 646.000 631.490 650.000 ;
    END
  END key_i[51]
  PIN key_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END key_i[52]
  PIN key_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END key_i[53]
  PIN key_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 190.440 650.000 191.040 ;
    END
  END key_i[54]
  PIN key_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END key_i[55]
  PIN key_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 553.930 646.000 554.210 650.000 ;
    END
  END key_i[56]
  PIN key_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 183.630 646.000 183.910 650.000 ;
    END
  END key_i[57]
  PIN key_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END key_i[58]
  PIN key_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 377.440 650.000 378.040 ;
    END
  END key_i[59]
  PIN key_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END key_i[5]
  PIN key_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 170.040 650.000 170.640 ;
    END
  END key_i[60]
  PIN key_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END key_i[61]
  PIN key_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 0.040 650.000 0.640 ;
    END
  END key_i[62]
  PIN key_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END key_i[63]
  PIN key_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END key_i[64]
  PIN key_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 265.240 650.000 265.840 ;
    END
  END key_i[65]
  PIN key_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 528.170 646.000 528.450 650.000 ;
    END
  END key_i[66]
  PIN key_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 567.840 650.000 568.440 ;
    END
  END key_i[67]
  PIN key_i[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 13.640 650.000 14.240 ;
    END
  END key_i[68]
  PIN key_i[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END key_i[69]
  PIN key_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 357.040 650.000 357.640 ;
    END
  END key_i[6]
  PIN key_i[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END key_i[70]
  PIN key_i[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 588.240 650.000 588.840 ;
    END
  END key_i[71]
  PIN key_i[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 502.410 646.000 502.690 650.000 ;
    END
  END key_i[72]
  PIN key_i[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 54.440 650.000 55.040 ;
    END
  END key_i[73]
  PIN key_i[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 476.650 646.000 476.930 650.000 ;
    END
  END key_i[74]
  PIN key_i[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END key_i[75]
  PIN key_i[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END key_i[76]
  PIN key_i[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END key_i[77]
  PIN key_i[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END key_i[78]
  PIN key_i[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END key_i[79]
  PIN key_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END key_i[7]
  PIN key_i[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END key_i[80]
  PIN key_i[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 646.000 196.790 650.000 ;
    END
  END key_i[81]
  PIN key_i[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END key_i[82]
  PIN key_i[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END key_i[83]
  PIN key_i[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END key_i[84]
  PIN key_i[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 354.290 646.000 354.570 650.000 ;
    END
  END key_i[85]
  PIN key_i[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 209.390 646.000 209.670 650.000 ;
    END
  END key_i[86]
  PIN key_i[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END key_i[87]
  PIN key_i[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 457.330 646.000 457.610 650.000 ;
    END
  END key_i[88]
  PIN key_i[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 163.240 650.000 163.840 ;
    END
  END key_i[89]
  PIN key_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END key_i[8]
  PIN key_i[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 493.040 650.000 493.640 ;
    END
  END key_i[90]
  PIN key_i[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END key_i[91]
  PIN key_i[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END key_i[92]
  PIN key_i[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END key_i[93]
  PIN key_i[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 646.000 472.640 650.000 473.240 ;
    END
  END key_i[94]
  PIN key_i[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END key_i[95]
  PIN key_i[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 438.010 646.000 438.290 650.000 ;
    END
  END key_i[96]
  PIN key_i[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 425.130 646.000 425.410 650.000 ;
    END
  END key_i[97]
  PIN key_i[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END key_i[98]
  PIN key_i[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 646.000 87.310 650.000 ;
    END
  END key_i[99]
  PIN key_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END key_i[9]
  PIN load_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END load_i
  PIN ready_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END ready_o
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 646.000 306.040 650.000 306.640 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.720 10.640 191.320 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.720 10.640 371.320 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 549.720 10.640 551.320 636.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 99.720 10.640 101.320 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.720 10.640 281.320 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.720 10.640 461.320 636.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 639.720 10.640 641.320 636.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 644.460 636.565 ;
      LAYER met1 ;
        RECT 0.070 9.220 648.990 638.480 ;
      LAYER met2 ;
        RECT 0.650 645.720 6.250 646.410 ;
        RECT 7.090 645.720 12.690 646.410 ;
        RECT 13.530 645.720 22.350 646.410 ;
        RECT 23.190 645.720 28.790 646.410 ;
        RECT 29.630 645.720 35.230 646.410 ;
        RECT 36.070 645.720 41.670 646.410 ;
        RECT 42.510 645.720 48.110 646.410 ;
        RECT 48.950 645.720 54.550 646.410 ;
        RECT 55.390 645.720 60.990 646.410 ;
        RECT 61.830 645.720 67.430 646.410 ;
        RECT 68.270 645.720 73.870 646.410 ;
        RECT 74.710 645.720 80.310 646.410 ;
        RECT 81.150 645.720 86.750 646.410 ;
        RECT 87.590 645.720 93.190 646.410 ;
        RECT 94.030 645.720 99.630 646.410 ;
        RECT 100.470 645.720 106.070 646.410 ;
        RECT 106.910 645.720 112.510 646.410 ;
        RECT 113.350 645.720 118.950 646.410 ;
        RECT 119.790 645.720 125.390 646.410 ;
        RECT 126.230 645.720 131.830 646.410 ;
        RECT 132.670 645.720 138.270 646.410 ;
        RECT 139.110 645.720 144.710 646.410 ;
        RECT 145.550 645.720 151.150 646.410 ;
        RECT 151.990 645.720 157.590 646.410 ;
        RECT 158.430 645.720 164.030 646.410 ;
        RECT 164.870 645.720 170.470 646.410 ;
        RECT 171.310 645.720 176.910 646.410 ;
        RECT 177.750 645.720 183.350 646.410 ;
        RECT 184.190 645.720 189.790 646.410 ;
        RECT 190.630 645.720 196.230 646.410 ;
        RECT 197.070 645.720 202.670 646.410 ;
        RECT 203.510 645.720 209.110 646.410 ;
        RECT 209.950 645.720 215.550 646.410 ;
        RECT 216.390 645.720 221.990 646.410 ;
        RECT 222.830 645.720 228.430 646.410 ;
        RECT 229.270 645.720 234.870 646.410 ;
        RECT 235.710 645.720 241.310 646.410 ;
        RECT 242.150 645.720 247.750 646.410 ;
        RECT 248.590 645.720 254.190 646.410 ;
        RECT 255.030 645.720 260.630 646.410 ;
        RECT 261.470 645.720 267.070 646.410 ;
        RECT 267.910 645.720 273.510 646.410 ;
        RECT 274.350 645.720 279.950 646.410 ;
        RECT 280.790 645.720 286.390 646.410 ;
        RECT 287.230 645.720 292.830 646.410 ;
        RECT 293.670 645.720 299.270 646.410 ;
        RECT 300.110 645.720 305.710 646.410 ;
        RECT 306.550 645.720 312.150 646.410 ;
        RECT 312.990 645.720 318.590 646.410 ;
        RECT 319.430 645.720 325.030 646.410 ;
        RECT 325.870 645.720 334.690 646.410 ;
        RECT 335.530 645.720 341.130 646.410 ;
        RECT 341.970 645.720 347.570 646.410 ;
        RECT 348.410 645.720 354.010 646.410 ;
        RECT 354.850 645.720 360.450 646.410 ;
        RECT 361.290 645.720 366.890 646.410 ;
        RECT 367.730 645.720 373.330 646.410 ;
        RECT 374.170 645.720 379.770 646.410 ;
        RECT 380.610 645.720 386.210 646.410 ;
        RECT 387.050 645.720 392.650 646.410 ;
        RECT 393.490 645.720 399.090 646.410 ;
        RECT 399.930 645.720 405.530 646.410 ;
        RECT 406.370 645.720 411.970 646.410 ;
        RECT 412.810 645.720 418.410 646.410 ;
        RECT 419.250 645.720 424.850 646.410 ;
        RECT 425.690 645.720 431.290 646.410 ;
        RECT 432.130 645.720 437.730 646.410 ;
        RECT 438.570 645.720 444.170 646.410 ;
        RECT 445.010 645.720 450.610 646.410 ;
        RECT 451.450 645.720 457.050 646.410 ;
        RECT 457.890 645.720 463.490 646.410 ;
        RECT 464.330 645.720 469.930 646.410 ;
        RECT 470.770 645.720 476.370 646.410 ;
        RECT 477.210 645.720 482.810 646.410 ;
        RECT 483.650 645.720 489.250 646.410 ;
        RECT 490.090 645.720 495.690 646.410 ;
        RECT 496.530 645.720 502.130 646.410 ;
        RECT 502.970 645.720 508.570 646.410 ;
        RECT 509.410 645.720 515.010 646.410 ;
        RECT 515.850 645.720 521.450 646.410 ;
        RECT 522.290 645.720 527.890 646.410 ;
        RECT 528.730 645.720 534.330 646.410 ;
        RECT 535.170 645.720 540.770 646.410 ;
        RECT 541.610 645.720 547.210 646.410 ;
        RECT 548.050 645.720 553.650 646.410 ;
        RECT 554.490 645.720 560.090 646.410 ;
        RECT 560.930 645.720 566.530 646.410 ;
        RECT 567.370 645.720 572.970 646.410 ;
        RECT 573.810 645.720 579.410 646.410 ;
        RECT 580.250 645.720 585.850 646.410 ;
        RECT 586.690 645.720 592.290 646.410 ;
        RECT 593.130 645.720 598.730 646.410 ;
        RECT 599.570 645.720 605.170 646.410 ;
        RECT 606.010 645.720 611.610 646.410 ;
        RECT 612.450 645.720 618.050 646.410 ;
        RECT 618.890 645.720 624.490 646.410 ;
        RECT 625.330 645.720 630.930 646.410 ;
        RECT 631.770 645.720 637.370 646.410 ;
        RECT 638.210 645.720 643.810 646.410 ;
        RECT 644.650 645.720 648.970 646.410 ;
        RECT 0.100 4.280 648.970 645.720 ;
        RECT 0.650 0.155 6.250 4.280 ;
        RECT 7.090 0.155 12.690 4.280 ;
        RECT 13.530 0.155 19.130 4.280 ;
        RECT 19.970 0.155 25.570 4.280 ;
        RECT 26.410 0.155 32.010 4.280 ;
        RECT 32.850 0.155 38.450 4.280 ;
        RECT 39.290 0.155 44.890 4.280 ;
        RECT 45.730 0.155 51.330 4.280 ;
        RECT 52.170 0.155 57.770 4.280 ;
        RECT 58.610 0.155 64.210 4.280 ;
        RECT 65.050 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 83.530 4.280 ;
        RECT 84.370 0.155 89.970 4.280 ;
        RECT 90.810 0.155 96.410 4.280 ;
        RECT 97.250 0.155 102.850 4.280 ;
        RECT 103.690 0.155 109.290 4.280 ;
        RECT 110.130 0.155 115.730 4.280 ;
        RECT 116.570 0.155 122.170 4.280 ;
        RECT 123.010 0.155 128.610 4.280 ;
        RECT 129.450 0.155 135.050 4.280 ;
        RECT 135.890 0.155 141.490 4.280 ;
        RECT 142.330 0.155 147.930 4.280 ;
        RECT 148.770 0.155 154.370 4.280 ;
        RECT 155.210 0.155 160.810 4.280 ;
        RECT 161.650 0.155 167.250 4.280 ;
        RECT 168.090 0.155 173.690 4.280 ;
        RECT 174.530 0.155 180.130 4.280 ;
        RECT 180.970 0.155 186.570 4.280 ;
        RECT 187.410 0.155 193.010 4.280 ;
        RECT 193.850 0.155 199.450 4.280 ;
        RECT 200.290 0.155 205.890 4.280 ;
        RECT 206.730 0.155 212.330 4.280 ;
        RECT 213.170 0.155 218.770 4.280 ;
        RECT 219.610 0.155 225.210 4.280 ;
        RECT 226.050 0.155 231.650 4.280 ;
        RECT 232.490 0.155 238.090 4.280 ;
        RECT 238.930 0.155 244.530 4.280 ;
        RECT 245.370 0.155 250.970 4.280 ;
        RECT 251.810 0.155 257.410 4.280 ;
        RECT 258.250 0.155 263.850 4.280 ;
        RECT 264.690 0.155 270.290 4.280 ;
        RECT 271.130 0.155 276.730 4.280 ;
        RECT 277.570 0.155 283.170 4.280 ;
        RECT 284.010 0.155 289.610 4.280 ;
        RECT 290.450 0.155 296.050 4.280 ;
        RECT 296.890 0.155 302.490 4.280 ;
        RECT 303.330 0.155 308.930 4.280 ;
        RECT 309.770 0.155 318.590 4.280 ;
        RECT 319.430 0.155 325.030 4.280 ;
        RECT 325.870 0.155 331.470 4.280 ;
        RECT 332.310 0.155 337.910 4.280 ;
        RECT 338.750 0.155 344.350 4.280 ;
        RECT 345.190 0.155 350.790 4.280 ;
        RECT 351.630 0.155 357.230 4.280 ;
        RECT 358.070 0.155 363.670 4.280 ;
        RECT 364.510 0.155 370.110 4.280 ;
        RECT 370.950 0.155 376.550 4.280 ;
        RECT 377.390 0.155 382.990 4.280 ;
        RECT 383.830 0.155 389.430 4.280 ;
        RECT 390.270 0.155 395.870 4.280 ;
        RECT 396.710 0.155 402.310 4.280 ;
        RECT 403.150 0.155 408.750 4.280 ;
        RECT 409.590 0.155 415.190 4.280 ;
        RECT 416.030 0.155 421.630 4.280 ;
        RECT 422.470 0.155 428.070 4.280 ;
        RECT 428.910 0.155 434.510 4.280 ;
        RECT 435.350 0.155 440.950 4.280 ;
        RECT 441.790 0.155 447.390 4.280 ;
        RECT 448.230 0.155 453.830 4.280 ;
        RECT 454.670 0.155 460.270 4.280 ;
        RECT 461.110 0.155 466.710 4.280 ;
        RECT 467.550 0.155 473.150 4.280 ;
        RECT 473.990 0.155 479.590 4.280 ;
        RECT 480.430 0.155 486.030 4.280 ;
        RECT 486.870 0.155 492.470 4.280 ;
        RECT 493.310 0.155 498.910 4.280 ;
        RECT 499.750 0.155 505.350 4.280 ;
        RECT 506.190 0.155 511.790 4.280 ;
        RECT 512.630 0.155 518.230 4.280 ;
        RECT 519.070 0.155 524.670 4.280 ;
        RECT 525.510 0.155 531.110 4.280 ;
        RECT 531.950 0.155 537.550 4.280 ;
        RECT 538.390 0.155 543.990 4.280 ;
        RECT 544.830 0.155 550.430 4.280 ;
        RECT 551.270 0.155 556.870 4.280 ;
        RECT 557.710 0.155 563.310 4.280 ;
        RECT 564.150 0.155 569.750 4.280 ;
        RECT 570.590 0.155 576.190 4.280 ;
        RECT 577.030 0.155 582.630 4.280 ;
        RECT 583.470 0.155 589.070 4.280 ;
        RECT 589.910 0.155 595.510 4.280 ;
        RECT 596.350 0.155 601.950 4.280 ;
        RECT 602.790 0.155 608.390 4.280 ;
        RECT 609.230 0.155 614.830 4.280 ;
        RECT 615.670 0.155 621.270 4.280 ;
        RECT 622.110 0.155 627.710 4.280 ;
        RECT 628.550 0.155 637.370 4.280 ;
        RECT 638.210 0.155 643.810 4.280 ;
        RECT 644.650 0.155 648.970 4.280 ;
      LAYER met3 ;
        RECT 4.400 642.240 645.600 643.105 ;
        RECT 3.990 636.840 648.995 642.240 ;
        RECT 4.400 635.440 645.600 636.840 ;
        RECT 3.990 630.040 648.995 635.440 ;
        RECT 4.400 628.640 645.600 630.040 ;
        RECT 3.990 623.240 648.995 628.640 ;
        RECT 4.400 621.840 645.600 623.240 ;
        RECT 3.990 616.440 648.995 621.840 ;
        RECT 4.400 615.040 645.600 616.440 ;
        RECT 3.990 609.640 648.995 615.040 ;
        RECT 4.400 608.240 645.600 609.640 ;
        RECT 3.990 602.840 648.995 608.240 ;
        RECT 4.400 601.440 645.600 602.840 ;
        RECT 3.990 596.040 648.995 601.440 ;
        RECT 4.400 594.640 645.600 596.040 ;
        RECT 3.990 589.240 648.995 594.640 ;
        RECT 4.400 587.840 645.600 589.240 ;
        RECT 3.990 582.440 648.995 587.840 ;
        RECT 4.400 581.040 645.600 582.440 ;
        RECT 3.990 575.640 648.995 581.040 ;
        RECT 4.400 574.240 645.600 575.640 ;
        RECT 3.990 568.840 648.995 574.240 ;
        RECT 4.400 567.440 645.600 568.840 ;
        RECT 3.990 562.040 648.995 567.440 ;
        RECT 4.400 560.640 645.600 562.040 ;
        RECT 3.990 555.240 648.995 560.640 ;
        RECT 4.400 553.840 645.600 555.240 ;
        RECT 3.990 548.440 648.995 553.840 ;
        RECT 4.400 547.040 645.600 548.440 ;
        RECT 3.990 541.640 648.995 547.040 ;
        RECT 4.400 540.240 645.600 541.640 ;
        RECT 3.990 534.840 648.995 540.240 ;
        RECT 4.400 533.440 645.600 534.840 ;
        RECT 3.990 528.040 648.995 533.440 ;
        RECT 4.400 526.640 645.600 528.040 ;
        RECT 3.990 521.240 648.995 526.640 ;
        RECT 4.400 519.840 645.600 521.240 ;
        RECT 3.990 514.440 648.995 519.840 ;
        RECT 4.400 513.040 645.600 514.440 ;
        RECT 3.990 507.640 648.995 513.040 ;
        RECT 4.400 506.240 645.600 507.640 ;
        RECT 3.990 500.840 648.995 506.240 ;
        RECT 4.400 499.440 645.600 500.840 ;
        RECT 3.990 494.040 648.995 499.440 ;
        RECT 4.400 492.640 645.600 494.040 ;
        RECT 3.990 487.240 648.995 492.640 ;
        RECT 4.400 485.840 645.600 487.240 ;
        RECT 3.990 480.440 648.995 485.840 ;
        RECT 4.400 479.040 645.600 480.440 ;
        RECT 3.990 473.640 648.995 479.040 ;
        RECT 4.400 472.240 645.600 473.640 ;
        RECT 3.990 466.840 648.995 472.240 ;
        RECT 4.400 465.440 645.600 466.840 ;
        RECT 3.990 460.040 648.995 465.440 ;
        RECT 4.400 458.640 645.600 460.040 ;
        RECT 3.990 453.240 648.995 458.640 ;
        RECT 4.400 451.840 645.600 453.240 ;
        RECT 3.990 446.440 648.995 451.840 ;
        RECT 4.400 445.040 645.600 446.440 ;
        RECT 3.990 439.640 648.995 445.040 ;
        RECT 4.400 438.240 645.600 439.640 ;
        RECT 3.990 432.840 648.995 438.240 ;
        RECT 4.400 431.440 645.600 432.840 ;
        RECT 3.990 426.040 648.995 431.440 ;
        RECT 4.400 424.640 645.600 426.040 ;
        RECT 3.990 419.240 648.995 424.640 ;
        RECT 4.400 417.840 645.600 419.240 ;
        RECT 3.990 412.440 648.995 417.840 ;
        RECT 4.400 411.040 645.600 412.440 ;
        RECT 3.990 405.640 648.995 411.040 ;
        RECT 4.400 404.240 645.600 405.640 ;
        RECT 3.990 398.840 648.995 404.240 ;
        RECT 4.400 397.440 645.600 398.840 ;
        RECT 3.990 392.040 648.995 397.440 ;
        RECT 4.400 390.640 645.600 392.040 ;
        RECT 3.990 385.240 648.995 390.640 ;
        RECT 4.400 383.840 645.600 385.240 ;
        RECT 3.990 378.440 648.995 383.840 ;
        RECT 4.400 377.040 645.600 378.440 ;
        RECT 3.990 371.640 648.995 377.040 ;
        RECT 4.400 370.240 645.600 371.640 ;
        RECT 3.990 364.840 648.995 370.240 ;
        RECT 4.400 363.440 645.600 364.840 ;
        RECT 3.990 358.040 648.995 363.440 ;
        RECT 4.400 356.640 645.600 358.040 ;
        RECT 3.990 351.240 648.995 356.640 ;
        RECT 4.400 349.840 645.600 351.240 ;
        RECT 3.990 344.440 648.995 349.840 ;
        RECT 4.400 343.040 645.600 344.440 ;
        RECT 3.990 337.640 648.995 343.040 ;
        RECT 4.400 336.240 645.600 337.640 ;
        RECT 3.990 330.840 648.995 336.240 ;
        RECT 3.990 329.440 645.600 330.840 ;
        RECT 3.990 327.440 648.995 329.440 ;
        RECT 4.400 326.040 648.995 327.440 ;
        RECT 3.990 324.040 648.995 326.040 ;
        RECT 3.990 322.640 645.600 324.040 ;
        RECT 3.990 320.640 648.995 322.640 ;
        RECT 4.400 319.240 648.995 320.640 ;
        RECT 3.990 317.240 648.995 319.240 ;
        RECT 3.990 315.840 645.600 317.240 ;
        RECT 3.990 313.840 648.995 315.840 ;
        RECT 4.400 312.440 648.995 313.840 ;
        RECT 3.990 307.040 648.995 312.440 ;
        RECT 4.400 305.640 645.600 307.040 ;
        RECT 3.990 300.240 648.995 305.640 ;
        RECT 4.400 298.840 645.600 300.240 ;
        RECT 3.990 293.440 648.995 298.840 ;
        RECT 4.400 292.040 645.600 293.440 ;
        RECT 3.990 286.640 648.995 292.040 ;
        RECT 4.400 285.240 645.600 286.640 ;
        RECT 3.990 279.840 648.995 285.240 ;
        RECT 4.400 278.440 645.600 279.840 ;
        RECT 3.990 273.040 648.995 278.440 ;
        RECT 4.400 271.640 645.600 273.040 ;
        RECT 3.990 266.240 648.995 271.640 ;
        RECT 4.400 264.840 645.600 266.240 ;
        RECT 3.990 259.440 648.995 264.840 ;
        RECT 4.400 258.040 645.600 259.440 ;
        RECT 3.990 252.640 648.995 258.040 ;
        RECT 4.400 251.240 645.600 252.640 ;
        RECT 3.990 245.840 648.995 251.240 ;
        RECT 4.400 244.440 645.600 245.840 ;
        RECT 3.990 239.040 648.995 244.440 ;
        RECT 4.400 237.640 645.600 239.040 ;
        RECT 3.990 232.240 648.995 237.640 ;
        RECT 4.400 230.840 645.600 232.240 ;
        RECT 3.990 225.440 648.995 230.840 ;
        RECT 4.400 224.040 645.600 225.440 ;
        RECT 3.990 218.640 648.995 224.040 ;
        RECT 4.400 217.240 645.600 218.640 ;
        RECT 3.990 211.840 648.995 217.240 ;
        RECT 4.400 210.440 645.600 211.840 ;
        RECT 3.990 205.040 648.995 210.440 ;
        RECT 4.400 203.640 645.600 205.040 ;
        RECT 3.990 198.240 648.995 203.640 ;
        RECT 4.400 196.840 645.600 198.240 ;
        RECT 3.990 191.440 648.995 196.840 ;
        RECT 4.400 190.040 645.600 191.440 ;
        RECT 3.990 184.640 648.995 190.040 ;
        RECT 4.400 183.240 645.600 184.640 ;
        RECT 3.990 177.840 648.995 183.240 ;
        RECT 4.400 176.440 645.600 177.840 ;
        RECT 3.990 171.040 648.995 176.440 ;
        RECT 4.400 169.640 645.600 171.040 ;
        RECT 3.990 164.240 648.995 169.640 ;
        RECT 4.400 162.840 645.600 164.240 ;
        RECT 3.990 157.440 648.995 162.840 ;
        RECT 4.400 156.040 645.600 157.440 ;
        RECT 3.990 150.640 648.995 156.040 ;
        RECT 4.400 149.240 645.600 150.640 ;
        RECT 3.990 143.840 648.995 149.240 ;
        RECT 4.400 142.440 645.600 143.840 ;
        RECT 3.990 137.040 648.995 142.440 ;
        RECT 4.400 135.640 645.600 137.040 ;
        RECT 3.990 130.240 648.995 135.640 ;
        RECT 4.400 128.840 645.600 130.240 ;
        RECT 3.990 123.440 648.995 128.840 ;
        RECT 4.400 122.040 645.600 123.440 ;
        RECT 3.990 116.640 648.995 122.040 ;
        RECT 4.400 115.240 645.600 116.640 ;
        RECT 3.990 109.840 648.995 115.240 ;
        RECT 4.400 108.440 645.600 109.840 ;
        RECT 3.990 103.040 648.995 108.440 ;
        RECT 4.400 101.640 645.600 103.040 ;
        RECT 3.990 96.240 648.995 101.640 ;
        RECT 4.400 94.840 645.600 96.240 ;
        RECT 3.990 89.440 648.995 94.840 ;
        RECT 4.400 88.040 645.600 89.440 ;
        RECT 3.990 82.640 648.995 88.040 ;
        RECT 4.400 81.240 645.600 82.640 ;
        RECT 3.990 75.840 648.995 81.240 ;
        RECT 4.400 74.440 645.600 75.840 ;
        RECT 3.990 69.040 648.995 74.440 ;
        RECT 4.400 67.640 645.600 69.040 ;
        RECT 3.990 62.240 648.995 67.640 ;
        RECT 4.400 60.840 645.600 62.240 ;
        RECT 3.990 55.440 648.995 60.840 ;
        RECT 4.400 54.040 645.600 55.440 ;
        RECT 3.990 48.640 648.995 54.040 ;
        RECT 4.400 47.240 645.600 48.640 ;
        RECT 3.990 41.840 648.995 47.240 ;
        RECT 4.400 40.440 645.600 41.840 ;
        RECT 3.990 35.040 648.995 40.440 ;
        RECT 4.400 33.640 645.600 35.040 ;
        RECT 3.990 28.240 648.995 33.640 ;
        RECT 4.400 26.840 645.600 28.240 ;
        RECT 3.990 21.440 648.995 26.840 ;
        RECT 4.400 20.040 645.600 21.440 ;
        RECT 3.990 14.640 648.995 20.040 ;
        RECT 4.400 13.240 645.600 14.640 ;
        RECT 3.990 7.840 648.995 13.240 ;
        RECT 4.400 6.440 645.600 7.840 ;
        RECT 3.990 1.040 648.995 6.440 ;
        RECT 3.990 0.175 645.600 1.040 ;
      LAYER met4 ;
        RECT 119.895 637.120 589.425 639.025 ;
        RECT 119.895 10.240 189.320 637.120 ;
        RECT 191.720 10.240 279.320 637.120 ;
        RECT 281.720 10.240 369.320 637.120 ;
        RECT 371.720 10.240 459.320 637.120 ;
        RECT 461.720 10.240 549.320 637.120 ;
        RECT 551.720 10.240 589.425 637.120 ;
        RECT 119.895 7.655 589.425 10.240 ;
  END
END aes_Trojan
END LIBRARY

