// This is the unpowered netlist.
module des (clk,
    decrypt,
    desIn,
    desOut,
    key,
    roundSel);
 input clk;
 input decrypt;
 input [63:0] desIn;
 output [63:0] desOut;
 input [55:0] key;
 input [3:0] roundSel;

 wire \L[10] ;
 wire \L[11] ;
 wire \L[12] ;
 wire \L[13] ;
 wire \L[14] ;
 wire \L[15] ;
 wire \L[16] ;
 wire \L[17] ;
 wire \L[18] ;
 wire \L[19] ;
 wire \L[1] ;
 wire \L[20] ;
 wire \L[21] ;
 wire \L[22] ;
 wire \L[23] ;
 wire \L[24] ;
 wire \L[25] ;
 wire \L[26] ;
 wire \L[27] ;
 wire \L[28] ;
 wire \L[29] ;
 wire \L[2] ;
 wire \L[30] ;
 wire \L[31] ;
 wire \L[32] ;
 wire \L[3] ;
 wire \L[4] ;
 wire \L[5] ;
 wire \L[6] ;
 wire \L[7] ;
 wire \L[8] ;
 wire \L[9] ;
 wire \R[10] ;
 wire \R[11] ;
 wire \R[12] ;
 wire \R[13] ;
 wire \R[14] ;
 wire \R[15] ;
 wire \R[16] ;
 wire \R[17] ;
 wire \R[18] ;
 wire \R[19] ;
 wire \R[1] ;
 wire \R[20] ;
 wire \R[21] ;
 wire \R[22] ;
 wire \R[23] ;
 wire \R[24] ;
 wire \R[25] ;
 wire \R[26] ;
 wire \R[27] ;
 wire \R[28] ;
 wire \R[29] ;
 wire \R[2] ;
 wire \R[30] ;
 wire \R[31] ;
 wire \R[32] ;
 wire \R[3] ;
 wire \R[4] ;
 wire \R[5] ;
 wire \R[6] ;
 wire \R[7] ;
 wire \R[8] ;
 wire \R[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net142));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__buf_6 _1309_ (.A(net125),
    .X(_0599_));
 sky130_fd_sc_hd__nor4_4 _1310_ (.A(_0599_),
    .B(net124),
    .C(net122),
    .D(net123),
    .Y(_0600_));
 sky130_fd_sc_hd__mux2_1 _1311_ (.A0(\R[32] ),
    .A1(net54),
    .S(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__clkbuf_4 _1312_ (.A(_0601_),
    .X(net178));
 sky130_fd_sc_hd__mux2_1 _1313_ (.A0(\R[31] ),
    .A1(net45),
    .S(net190),
    .X(_0602_));
 sky130_fd_sc_hd__buf_2 _1314_ (.A(_0602_),
    .X(net169));
 sky130_fd_sc_hd__mux2_1 _1315_ (.A0(\R[30] ),
    .A1(net37),
    .S(net190),
    .X(_0603_));
 sky130_fd_sc_hd__clkbuf_2 _1316_ (.A(_0603_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 _1317_ (.A(net190),
    .X(_0604_));
 sky130_fd_sc_hd__buf_6 _1318_ (.A(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _1319_ (.A0(\R[29] ),
    .A1(net28),
    .S(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__clkbuf_4 _1320_ (.A(_0606_),
    .X(net152));
 sky130_fd_sc_hd__mux2_1 _1321_ (.A0(\R[28] ),
    .A1(net19),
    .S(_0600_),
    .X(_0607_));
 sky130_fd_sc_hd__buf_4 _1322_ (.A(_0607_),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_8 _1323_ (.A(net190),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _1324_ (.A0(\R[27] ),
    .A1(net10),
    .S(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__buf_2 _1325_ (.A(_0609_),
    .X(net134));
 sky130_fd_sc_hd__mux2_1 _1326_ (.A0(\R[26] ),
    .A1(net65),
    .S(net190),
    .X(_0610_));
 sky130_fd_sc_hd__buf_2 _1327_ (.A(_0610_),
    .X(net189));
 sky130_fd_sc_hd__mux2_1 _1328_ (.A0(\R[25] ),
    .A1(net13),
    .S(_0604_),
    .X(_0611_));
 sky130_fd_sc_hd__clkbuf_8 _1329_ (.A(_0611_),
    .X(net137));
 sky130_fd_sc_hd__mux2_1 _1330_ (.A0(\R[24] ),
    .A1(net56),
    .S(_0604_),
    .X(_0612_));
 sky130_fd_sc_hd__buf_4 _1331_ (.A(_0612_),
    .X(net180));
 sky130_fd_sc_hd__mux2_1 _1332_ (.A0(\R[23] ),
    .A1(net48),
    .S(_0608_),
    .X(_0613_));
 sky130_fd_sc_hd__clkbuf_4 _1333_ (.A(_0613_),
    .X(net172));
 sky130_fd_sc_hd__mux2_1 _1334_ (.A0(\R[22] ),
    .A1(net39),
    .S(_0604_),
    .X(_0614_));
 sky130_fd_sc_hd__buf_4 _1335_ (.A(_0614_),
    .X(net163));
 sky130_fd_sc_hd__mux2_1 _1336_ (.A0(\R[21] ),
    .A1(net30),
    .S(_0604_),
    .X(_0615_));
 sky130_fd_sc_hd__clkbuf_8 _1337_ (.A(_0615_),
    .X(net154));
 sky130_fd_sc_hd__mux2_1 _1338_ (.A0(\R[20] ),
    .A1(net21),
    .S(_0608_),
    .X(_0616_));
 sky130_fd_sc_hd__buf_4 _1339_ (.A(_0616_),
    .X(net145));
 sky130_fd_sc_hd__mux2_1 _1340_ (.A0(\R[19] ),
    .A1(net12),
    .S(_0608_),
    .X(_0617_));
 sky130_fd_sc_hd__buf_2 _1341_ (.A(_0617_),
    .X(net136));
 sky130_fd_sc_hd__mux2_1 _1342_ (.A0(\R[18] ),
    .A1(net4),
    .S(_0604_),
    .X(_0618_));
 sky130_fd_sc_hd__buf_4 _1343_ (.A(_0618_),
    .X(net128));
 sky130_fd_sc_hd__mux2_1 _1344_ (.A0(\R[17] ),
    .A1(net35),
    .S(_0605_),
    .X(_0619_));
 sky130_fd_sc_hd__buf_4 _1345_ (.A(_0619_),
    .X(net159));
 sky130_fd_sc_hd__mux2_1 _1346_ (.A0(\R[16] ),
    .A1(net59),
    .S(net190),
    .X(_0620_));
 sky130_fd_sc_hd__buf_4 _1347_ (.A(_0620_),
    .X(net183));
 sky130_fd_sc_hd__or4_4 _1348_ (.A(_0599_),
    .B(net124),
    .C(net122),
    .D(net123),
    .X(_0621_));
 sky130_fd_sc_hd__or2_1 _1349_ (.A(net193),
    .B(_0608_),
    .X(_0622_));
 sky130_fd_sc_hd__o21ai_4 _1350_ (.A1(net50),
    .A2(_0621_),
    .B1(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _1351_ (.A(_0623_),
    .Y(net174));
 sky130_fd_sc_hd__mux2_1 _1352_ (.A0(\R[14] ),
    .A1(net41),
    .S(_0604_),
    .X(_0624_));
 sky130_fd_sc_hd__buf_4 _1353_ (.A(_0624_),
    .X(net165));
 sky130_fd_sc_hd__mux2_1 _1354_ (.A0(\R[13] ),
    .A1(net32),
    .S(_0605_),
    .X(_0625_));
 sky130_fd_sc_hd__buf_6 _1355_ (.A(_0625_),
    .X(net156));
 sky130_fd_sc_hd__or2_1 _1356_ (.A(\R[12] ),
    .B(_0604_),
    .X(_0626_));
 sky130_fd_sc_hd__o21ai_4 _1357_ (.A1(net23),
    .A2(_0621_),
    .B1(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__inv_2 _1358_ (.A(_0627_),
    .Y(net147));
 sky130_fd_sc_hd__mux2_1 _1359_ (.A0(\R[11] ),
    .A1(net15),
    .S(_0608_),
    .X(_0628_));
 sky130_fd_sc_hd__buf_2 _1360_ (.A(_0628_),
    .X(net139));
 sky130_fd_sc_hd__mux2_1 _1361_ (.A0(\R[10] ),
    .A1(net6),
    .S(_0604_),
    .X(_0629_));
 sky130_fd_sc_hd__clkbuf_4 _1362_ (.A(_0629_),
    .X(net130));
 sky130_fd_sc_hd__mux2_1 _1363_ (.A0(\R[9] ),
    .A1(net57),
    .S(_0605_),
    .X(_0630_));
 sky130_fd_sc_hd__clkbuf_8 _1364_ (.A(_0630_),
    .X(net181));
 sky130_fd_sc_hd__mux2_1 _1365_ (.A0(\R[8] ),
    .A1(net61),
    .S(_0608_),
    .X(_0631_));
 sky130_fd_sc_hd__buf_4 _1366_ (.A(_0631_),
    .X(net185));
 sky130_fd_sc_hd__mux2_1 _1367_ (.A0(\R[7] ),
    .A1(net52),
    .S(_0600_),
    .X(_0632_));
 sky130_fd_sc_hd__clkbuf_2 _1368_ (.A(_0632_),
    .X(net176));
 sky130_fd_sc_hd__mux2_1 _1369_ (.A0(\R[6] ),
    .A1(net43),
    .S(_0608_),
    .X(_0633_));
 sky130_fd_sc_hd__clkbuf_4 _1370_ (.A(_0633_),
    .X(net167));
 sky130_fd_sc_hd__mux2_1 _1371_ (.A0(\R[5] ),
    .A1(net34),
    .S(_0604_),
    .X(_0634_));
 sky130_fd_sc_hd__buf_4 _1372_ (.A(_0634_),
    .X(net158));
 sky130_fd_sc_hd__mux2_1 _1373_ (.A0(\R[4] ),
    .A1(net26),
    .S(_0608_),
    .X(_0635_));
 sky130_fd_sc_hd__buf_4 _1374_ (.A(_0635_),
    .X(net150));
 sky130_fd_sc_hd__mux2_1 _1375_ (.A0(\R[3] ),
    .A1(net17),
    .S(net190),
    .X(_0636_));
 sky130_fd_sc_hd__buf_2 _1376_ (.A(_0636_),
    .X(net141));
 sky130_fd_sc_hd__mux2_1 _1377_ (.A0(\R[2] ),
    .A1(net8),
    .S(_0608_),
    .X(_0637_));
 sky130_fd_sc_hd__buf_2 _1378_ (.A(_0637_),
    .X(net132));
 sky130_fd_sc_hd__mux2_1 _1379_ (.A0(\R[1] ),
    .A1(net63),
    .S(_0605_),
    .X(_0638_));
 sky130_fd_sc_hd__clkbuf_8 _1380_ (.A(_0638_),
    .X(net187));
 sky130_fd_sc_hd__xnor2_1 _1381_ (.A(_0599_),
    .B(net122),
    .Y(_0639_));
 sky130_fd_sc_hd__xor2_2 _1382_ (.A(_0599_),
    .B(net123),
    .X(_0640_));
 sky130_fd_sc_hd__xnor2_2 _1383_ (.A(_0599_),
    .B(net124),
    .Y(_0641_));
 sky130_fd_sc_hd__and3_1 _1384_ (.A(_0639_),
    .B(_0640_),
    .C(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__clkbuf_4 _1385_ (.A(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__buf_4 _1386_ (.A(_0643_),
    .X(_0644_));
 sky130_fd_sc_hd__xnor2_2 _1387_ (.A(_0599_),
    .B(net1),
    .Y(_0645_));
 sky130_fd_sc_hd__buf_2 _1388_ (.A(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__clkbuf_4 _1389_ (.A(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__or2_4 _1390_ (.A(net121),
    .B(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__xor2_4 _1391_ (.A(_0599_),
    .B(net1),
    .X(_0649_));
 sky130_fd_sc_hd__buf_2 _1392_ (.A(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__clkbuf_4 _1393_ (.A(_0650_),
    .X(_0651_));
 sky130_fd_sc_hd__or2_2 _1394_ (.A(net90),
    .B(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__xor2_2 _1395_ (.A(_0599_),
    .B(net122),
    .X(_0653_));
 sky130_fd_sc_hd__xnor2_1 _1396_ (.A(_0599_),
    .B(net123),
    .Y(_0654_));
 sky130_fd_sc_hd__and3_1 _1397_ (.A(_0653_),
    .B(_0654_),
    .C(_0641_),
    .X(_0655_));
 sky130_fd_sc_hd__clkbuf_4 _1398_ (.A(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__clkbuf_4 _1399_ (.A(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__clkbuf_4 _1400_ (.A(_0645_),
    .X(_0658_));
 sky130_fd_sc_hd__clkbuf_4 _1401_ (.A(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__or2_2 _1402_ (.A(net81),
    .B(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__clkbuf_4 _1403_ (.A(_0649_),
    .X(_0661_));
 sky130_fd_sc_hd__or2_2 _1404_ (.A(net104),
    .B(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__and3_1 _1405_ (.A(_0657_),
    .B(_0660_),
    .C(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__a31o_1 _1406_ (.A1(_0644_),
    .A2(_0648_),
    .A3(_0652_),
    .B1(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__xor2_1 _1407_ (.A(_0599_),
    .B(net124),
    .X(_0665_));
 sky130_fd_sc_hd__and3_1 _1408_ (.A(_0639_),
    .B(_0640_),
    .C(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__clkbuf_4 _1409_ (.A(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__clkbuf_4 _1410_ (.A(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__or2_2 _1411_ (.A(net86),
    .B(_0661_),
    .X(_0669_));
 sky130_fd_sc_hd__clkbuf_4 _1412_ (.A(_0645_),
    .X(_0670_));
 sky130_fd_sc_hd__or2_1 _1413_ (.A(net120),
    .B(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__and3_1 _1414_ (.A(_0653_),
    .B(_0640_),
    .C(_0665_),
    .X(_0672_));
 sky130_fd_sc_hd__clkbuf_4 _1415_ (.A(_0672_),
    .X(_0673_));
 sky130_fd_sc_hd__clkbuf_4 _1416_ (.A(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_4 _1417_ (.A(_0649_),
    .X(_0675_));
 sky130_fd_sc_hd__or2_2 _1418_ (.A(net102),
    .B(_0675_),
    .X(_0676_));
 sky130_fd_sc_hd__or2_2 _1419_ (.A(net109),
    .B(_0658_),
    .X(_0677_));
 sky130_fd_sc_hd__and3_1 _1420_ (.A(_0674_),
    .B(_0676_),
    .C(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__a31o_1 _1421_ (.A1(_0668_),
    .A2(_0669_),
    .A3(_0671_),
    .B1(_0678_),
    .X(_0679_));
 sky130_fd_sc_hd__and3_1 _1422_ (.A(_0653_),
    .B(_0640_),
    .C(_0641_),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_4 _1423_ (.A(_0680_),
    .X(_0681_));
 sky130_fd_sc_hd__buf_4 _1424_ (.A(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__or2_4 _1425_ (.A(net111),
    .B(_0647_),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_4 _1426_ (.A(_0650_),
    .X(_0684_));
 sky130_fd_sc_hd__or2_1 _1427_ (.A(net105),
    .B(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__and3_1 _1428_ (.A(_0653_),
    .B(_0654_),
    .C(_0665_),
    .X(_0686_));
 sky130_fd_sc_hd__clkbuf_4 _1429_ (.A(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__clkbuf_4 _1430_ (.A(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_4 _1431_ (.A(_0646_),
    .X(_0689_));
 sky130_fd_sc_hd__or2_2 _1432_ (.A(net80),
    .B(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__buf_2 _1433_ (.A(_0649_),
    .X(_0691_));
 sky130_fd_sc_hd__or2_4 _1434_ (.A(net71),
    .B(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__and3_2 _1435_ (.A(_0639_),
    .B(_0654_),
    .C(_0641_),
    .X(_0693_));
 sky130_fd_sc_hd__a31o_1 _1436_ (.A1(_0688_),
    .A2(_0690_),
    .A3(_0692_),
    .B1(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__and3_1 _1437_ (.A(_0639_),
    .B(_0654_),
    .C(_0665_),
    .X(_0695_));
 sky130_fd_sc_hd__buf_4 _1438_ (.A(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__clkbuf_4 _1439_ (.A(_0646_),
    .X(_0697_));
 sky130_fd_sc_hd__or2_2 _1440_ (.A(net95),
    .B(_0697_),
    .X(_0698_));
 sky130_fd_sc_hd__or2_2 _1441_ (.A(net66),
    .B(_0684_),
    .X(_0699_));
 sky130_fd_sc_hd__and3_1 _1442_ (.A(_0696_),
    .B(_0698_),
    .C(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__a311o_1 _1443_ (.A1(_0682_),
    .A2(_0683_),
    .A3(_0685_),
    .B1(_0694_),
    .C1(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__clkbuf_4 _1444_ (.A(_0675_),
    .X(_0702_));
 sky130_fd_sc_hd__or2_2 _1445_ (.A(net96),
    .B(_0702_),
    .X(_0703_));
 sky130_fd_sc_hd__or2_2 _1446_ (.A(net89),
    .B(_0646_),
    .X(_0704_));
 sky130_fd_sc_hd__nor2_1 _1447_ (.A(_0653_),
    .B(_0640_),
    .Y(_0705_));
 sky130_fd_sc_hd__clkbuf_4 _1448_ (.A(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__clkbuf_4 _1449_ (.A(_0641_),
    .X(_0707_));
 sky130_fd_sc_hd__nand2_2 _1450_ (.A(_0706_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__buf_4 _1451_ (.A(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__a21o_1 _1452_ (.A1(_0703_),
    .A2(_0704_),
    .B1(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__o31a_4 _1453_ (.A1(_0664_),
    .A2(_0679_),
    .A3(_0701_),
    .B1(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__xor2_4 _1454_ (.A(net137),
    .B(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__or2_2 _1455_ (.A(net90),
    .B(_0697_),
    .X(_0713_));
 sky130_fd_sc_hd__or2_2 _1456_ (.A(net79),
    .B(_0650_),
    .X(_0714_));
 sky130_fd_sc_hd__mux2_1 _1457_ (.A0(net94),
    .A1(net104),
    .S(_0651_),
    .X(_0715_));
 sky130_fd_sc_hd__clkbuf_4 _1458_ (.A(_0680_),
    .X(_0716_));
 sky130_fd_sc_hd__a32o_1 _1459_ (.A1(_0643_),
    .A2(_0713_),
    .A3(_0714_),
    .B1(_0715_),
    .B2(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__or2_2 _1460_ (.A(net120),
    .B(_0675_),
    .X(_0718_));
 sky130_fd_sc_hd__or2_2 _1461_ (.A(net73),
    .B(_0646_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _1462_ (.A0(net80),
    .A1(net88),
    .S(_0651_),
    .X(_0720_));
 sky130_fd_sc_hd__clkbuf_4 _1463_ (.A(_0667_),
    .X(_0721_));
 sky130_fd_sc_hd__a32o_1 _1464_ (.A1(_0688_),
    .A2(_0718_),
    .A3(_0719_),
    .B1(_0720_),
    .B2(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__or2_2 _1465_ (.A(net105),
    .B(_0647_),
    .X(_0723_));
 sky130_fd_sc_hd__or2_1 _1466_ (.A(net119),
    .B(_0684_),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _1467_ (.A0(net95),
    .A1(net103),
    .S(_0651_),
    .X(_0725_));
 sky130_fd_sc_hd__a32o_1 _1468_ (.A1(_0657_),
    .A2(_0723_),
    .A3(_0724_),
    .B1(_0725_),
    .B2(_0674_),
    .X(_0726_));
 sky130_fd_sc_hd__clkbuf_4 _1469_ (.A(_0641_),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _1470_ (.A0(net89),
    .A1(net109),
    .S(_0659_),
    .X(_0728_));
 sky130_fd_sc_hd__clkbuf_4 _1471_ (.A(_0705_),
    .X(_0729_));
 sky130_fd_sc_hd__o21a_1 _1472_ (.A1(_0727_),
    .A2(_0728_),
    .B1(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__or4_2 _1473_ (.A(_0717_),
    .B(_0722_),
    .C(_0726_),
    .D(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__or2_2 _1474_ (.A(net113),
    .B(_0658_),
    .X(_0732_));
 sky130_fd_sc_hd__a21o_1 _1475_ (.A1(_0699_),
    .A2(_0732_),
    .B1(_0709_),
    .X(_0733_));
 sky130_fd_sc_hd__nand3b_2 _1476_ (.A_N(net134),
    .B(_0731_),
    .C(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__a21bo_1 _1477_ (.A1(_0731_),
    .A2(_0733_),
    .B1_N(net134),
    .X(_0735_));
 sky130_fd_sc_hd__nand2_1 _1478_ (.A(_0734_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__clkbuf_4 _1479_ (.A(_0642_),
    .X(_0737_));
 sky130_fd_sc_hd__or2_2 _1480_ (.A(net103),
    .B(_0661_),
    .X(_0738_));
 sky130_fd_sc_hd__and3_1 _1481_ (.A(_0737_),
    .B(_0677_),
    .C(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__or2_2 _1482_ (.A(net79),
    .B(_0658_),
    .X(_0740_));
 sky130_fd_sc_hd__or2_2 _1483_ (.A(net73),
    .B(_0661_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(net89),
    .A1(net119),
    .S(_0661_),
    .X(_0742_));
 sky130_fd_sc_hd__a32o_1 _1485_ (.A1(_0696_),
    .A2(_0740_),
    .A3(_0741_),
    .B1(_0742_),
    .B2(_0687_),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(net90),
    .A1(net97),
    .S(_0661_),
    .X(_0744_));
 sky130_fd_sc_hd__a32o_1 _1487_ (.A1(_0662_),
    .A2(_0667_),
    .A3(_0732_),
    .B1(_0744_),
    .B2(_0673_),
    .X(_0745_));
 sky130_fd_sc_hd__or2_2 _1488_ (.A(net87),
    .B(_0675_),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _1489_ (.A0(net94),
    .A1(net88),
    .S(_0658_),
    .X(_0747_));
 sky130_fd_sc_hd__clkbuf_4 _1490_ (.A(_0680_),
    .X(_0748_));
 sky130_fd_sc_hd__a32o_1 _1491_ (.A1(_0656_),
    .A2(_0671_),
    .A3(_0746_),
    .B1(_0747_),
    .B2(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__or4_2 _1492_ (.A(_0739_),
    .B(_0743_),
    .C(_0745_),
    .D(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__clkbuf_4 _1493_ (.A(_0693_),
    .X(_0751_));
 sky130_fd_sc_hd__or2_2 _1494_ (.A(net80),
    .B(_0675_),
    .X(_0752_));
 sky130_fd_sc_hd__clkbuf_4 _1495_ (.A(_0670_),
    .X(_0753_));
 sky130_fd_sc_hd__or2_2 _1496_ (.A(net72),
    .B(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__and3_1 _1497_ (.A(_0751_),
    .B(_0752_),
    .C(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__o21ai_2 _1498_ (.A1(_0750_),
    .A2(_0755_),
    .B1(net189),
    .Y(_0756_));
 sky130_fd_sc_hd__or3_2 _1499_ (.A(net189),
    .B(_0750_),
    .C(_0755_),
    .X(_0757_));
 sky130_fd_sc_hd__and2_1 _1500_ (.A(_0756_),
    .B(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__buf_2 _1501_ (.A(_0758_),
    .X(_0759_));
 sky130_fd_sc_hd__nor2_1 _1502_ (.A(_0736_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__buf_2 _1503_ (.A(_0645_),
    .X(_0761_));
 sky130_fd_sc_hd__or2_2 _1504_ (.A(net71),
    .B(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__clkbuf_4 _1505_ (.A(_0649_),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_1 _1506_ (.A0(net80),
    .A1(net66),
    .S(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__a32o_1 _1507_ (.A1(_0643_),
    .A2(_0762_),
    .A3(_0718_),
    .B1(_0681_),
    .B2(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__or2_2 _1508_ (.A(net121),
    .B(_0763_),
    .X(_0766_));
 sky130_fd_sc_hd__or2_2 _1509_ (.A(net104),
    .B(_0761_),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _1510_ (.A0(net111),
    .A1(net90),
    .S(_0763_),
    .X(_0768_));
 sky130_fd_sc_hd__a32o_1 _1511_ (.A1(_0667_),
    .A2(_0766_),
    .A3(_0767_),
    .B1(_0768_),
    .B2(_0687_),
    .X(_0769_));
 sky130_fd_sc_hd__clkbuf_4 _1512_ (.A(_0650_),
    .X(_0770_));
 sky130_fd_sc_hd__or2_2 _1513_ (.A(net81),
    .B(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_1 _1514_ (.A0(net86),
    .A1(net109),
    .S(_0647_),
    .X(_0772_));
 sky130_fd_sc_hd__clkbuf_4 _1515_ (.A(_0655_),
    .X(_0773_));
 sky130_fd_sc_hd__a32o_1 _1516_ (.A1(_0673_),
    .A2(_0704_),
    .A3(_0771_),
    .B1(_0772_),
    .B2(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _1517_ (.A0(net105),
    .A1(net95),
    .S(_0761_),
    .X(_0775_));
 sky130_fd_sc_hd__o21a_1 _1518_ (.A1(_0707_),
    .A2(_0775_),
    .B1(_0706_),
    .X(_0776_));
 sky130_fd_sc_hd__or4_2 _1519_ (.A(_0765_),
    .B(_0769_),
    .C(_0774_),
    .D(_0776_),
    .X(_0777_));
 sky130_fd_sc_hd__or2_2 _1520_ (.A(net94),
    .B(_0670_),
    .X(_0778_));
 sky130_fd_sc_hd__clkbuf_4 _1521_ (.A(_0708_),
    .X(_0779_));
 sky130_fd_sc_hd__a21o_1 _1522_ (.A1(_0676_),
    .A2(_0778_),
    .B1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__nand3_2 _1523_ (.A(net143),
    .B(_0777_),
    .C(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__a21o_1 _1524_ (.A1(_0777_),
    .A2(_0780_),
    .B1(net143),
    .X(_0782_));
 sky130_fd_sc_hd__a22o_2 _1525_ (.A1(_0781_),
    .A2(_0782_),
    .B1(_0734_),
    .B2(_0735_),
    .X(_0783_));
 sky130_fd_sc_hd__nand4_4 _1526_ (.A(_0781_),
    .B(_0782_),
    .C(_0734_),
    .D(_0735_),
    .Y(_0784_));
 sky130_fd_sc_hd__nand2_4 _1527_ (.A(_0756_),
    .B(_0757_),
    .Y(_0785_));
 sky130_fd_sc_hd__a21o_1 _1528_ (.A1(_0783_),
    .A2(_0784_),
    .B1(_0785_),
    .X(_0786_));
 sky130_fd_sc_hd__and2b_1 _1529_ (.A_N(_0760_),
    .B(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__clkbuf_4 _1530_ (.A(_0751_),
    .X(_0788_));
 sky130_fd_sc_hd__or2_2 _1531_ (.A(net97),
    .B(_0650_),
    .X(_0789_));
 sky130_fd_sc_hd__clkbuf_4 _1532_ (.A(_0686_),
    .X(_0790_));
 sky130_fd_sc_hd__and3_1 _1533_ (.A(_0683_),
    .B(_0676_),
    .C(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__or2_2 _1534_ (.A(net112),
    .B(_0670_),
    .X(_0792_));
 sky130_fd_sc_hd__and3_1 _1535_ (.A(_0773_),
    .B(_0685_),
    .C(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__a311o_1 _1536_ (.A1(_0660_),
    .A2(_0682_),
    .A3(_0692_),
    .B1(_0791_),
    .C1(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__clkbuf_4 _1537_ (.A(_0702_),
    .X(_0795_));
 sky130_fd_sc_hd__buf_4 _1538_ (.A(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__clkbuf_4 _1539_ (.A(_0673_),
    .X(_0797_));
 sky130_fd_sc_hd__o211a_1 _1540_ (.A1(net72),
    .A2(_0796_),
    .B1(_0797_),
    .C1(_0690_),
    .X(_0798_));
 sky130_fd_sc_hd__buf_4 _1541_ (.A(_0696_),
    .X(_0799_));
 sky130_fd_sc_hd__and3_1 _1542_ (.A(_0648_),
    .B(_0799_),
    .C(_0669_),
    .X(_0800_));
 sky130_fd_sc_hd__or2_2 _1543_ (.A(net96),
    .B(_0689_),
    .X(_0801_));
 sky130_fd_sc_hd__or2_2 _1544_ (.A(net77),
    .B(_0691_),
    .X(_0802_));
 sky130_fd_sc_hd__and3_1 _1545_ (.A(_0698_),
    .B(_0721_),
    .C(_0802_),
    .X(_0803_));
 sky130_fd_sc_hd__a31o_1 _1546_ (.A1(_0644_),
    .A2(_0699_),
    .A3(_0801_),
    .B1(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__or4_2 _1547_ (.A(_0794_),
    .B(_0798_),
    .C(_0800_),
    .D(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__a31oi_2 _1548_ (.A1(_0788_),
    .A2(_0713_),
    .A3(_0789_),
    .B1(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__xnor2_2 _1549_ (.A(net152),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__inv_2 _1550_ (.A(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__nand2_1 _1551_ (.A(_0781_),
    .B(_0782_),
    .Y(_0809_));
 sky130_fd_sc_hd__buf_2 _1552_ (.A(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__nor2_1 _1553_ (.A(_0810_),
    .B(_0759_),
    .Y(_0811_));
 sky130_fd_sc_hd__xnor2_4 _1554_ (.A(net137),
    .B(_0711_),
    .Y(_0812_));
 sky130_fd_sc_hd__a31oi_1 _1555_ (.A1(_0810_),
    .A2(_0736_),
    .A3(_0759_),
    .B1(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__or3b_1 _1556_ (.A(_0760_),
    .B(_0811_),
    .C_N(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__o211a_1 _1557_ (.A1(_0712_),
    .A2(_0787_),
    .B1(_0808_),
    .C1(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__nand2_2 _1558_ (.A(_0783_),
    .B(_0784_),
    .Y(_0816_));
 sky130_fd_sc_hd__nand2_1 _1559_ (.A(_0712_),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__or3b_1 _1560_ (.A(_0712_),
    .B(_0811_),
    .C_N(_0783_),
    .X(_0818_));
 sky130_fd_sc_hd__buf_6 _1561_ (.A(_0788_),
    .X(_0819_));
 sky130_fd_sc_hd__or2_1 _1562_ (.A(net88),
    .B(_0770_),
    .X(_0820_));
 sky130_fd_sc_hd__buf_4 _1563_ (.A(_0668_),
    .X(_0821_));
 sky130_fd_sc_hd__buf_2 _1564_ (.A(_0646_),
    .X(_0822_));
 sky130_fd_sc_hd__or2_2 _1565_ (.A(net86),
    .B(_0822_),
    .X(_0823_));
 sky130_fd_sc_hd__or2_2 _1566_ (.A(net113),
    .B(_0702_),
    .X(_0824_));
 sky130_fd_sc_hd__clkbuf_4 _1567_ (.A(_0797_),
    .X(_0825_));
 sky130_fd_sc_hd__clkbuf_4 _1568_ (.A(_0716_),
    .X(_0826_));
 sky130_fd_sc_hd__and3_1 _1569_ (.A(_0826_),
    .B(_0703_),
    .C(_0754_),
    .X(_0827_));
 sky130_fd_sc_hd__a31o_1 _1570_ (.A1(_0825_),
    .A2(_0762_),
    .A3(_0724_),
    .B1(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__clkbuf_4 _1571_ (.A(_0696_),
    .X(_0829_));
 sky130_fd_sc_hd__or2_4 _1572_ (.A(net77),
    .B(_0646_),
    .X(_0830_));
 sky130_fd_sc_hd__or2_2 _1573_ (.A(net112),
    .B(_0650_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_4 _1574_ (.A(_0644_),
    .X(_0832_));
 sky130_fd_sc_hd__or2_2 _1575_ (.A(net87),
    .B(_0646_),
    .X(_0833_));
 sky130_fd_sc_hd__clkbuf_4 _1576_ (.A(_0687_),
    .X(_0834_));
 sky130_fd_sc_hd__or2_2 _1577_ (.A(net102),
    .B(_0647_),
    .X(_0835_));
 sky130_fd_sc_hd__and3_1 _1578_ (.A(_0834_),
    .B(_0789_),
    .C(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__a31o_1 _1579_ (.A1(_0832_),
    .A2(_0771_),
    .A3(_0833_),
    .B1(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__buf_4 _1580_ (.A(_0753_),
    .X(_0838_));
 sky130_fd_sc_hd__buf_4 _1581_ (.A(_0656_),
    .X(_0839_));
 sky130_fd_sc_hd__clkbuf_4 _1582_ (.A(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__o211a_1 _1583_ (.A1(net103),
    .A2(_0838_),
    .B1(_0840_),
    .C1(_0766_),
    .X(_0841_));
 sky130_fd_sc_hd__a311o_1 _1584_ (.A1(_0829_),
    .A2(_0830_),
    .A3(_0831_),
    .B1(_0837_),
    .C1(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__a311o_1 _1585_ (.A1(_0821_),
    .A2(_0823_),
    .A3(_0824_),
    .B1(_0828_),
    .C1(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__a31o_2 _1586_ (.A1(_0683_),
    .A2(_0819_),
    .A3(_0820_),
    .B1(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__xnor2_4 _1587_ (.A(net180),
    .B(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__a31o_1 _1588_ (.A1(_0807_),
    .A2(_0817_),
    .A3(_0818_),
    .B1(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__xnor2_1 _1589_ (.A(_0785_),
    .B(_0816_),
    .Y(_0847_));
 sky130_fd_sc_hd__xnor2_1 _1590_ (.A(_0810_),
    .B(_0759_),
    .Y(_0848_));
 sky130_fd_sc_hd__and2_1 _1591_ (.A(_0734_),
    .B(_0735_),
    .X(_0849_));
 sky130_fd_sc_hd__nor2_1 _1592_ (.A(_0849_),
    .B(_0785_),
    .Y(_0850_));
 sky130_fd_sc_hd__or2b_1 _1593_ (.A(_0850_),
    .B_N(_0816_),
    .X(_0851_));
 sky130_fd_sc_hd__nor2_1 _1594_ (.A(_0850_),
    .B(_0848_),
    .Y(_0852_));
 sky130_fd_sc_hd__mux4_1 _1595_ (.A0(_0847_),
    .A1(_0848_),
    .A2(_0851_),
    .A3(_0852_),
    .S0(_0812_),
    .S1(_0808_),
    .X(_0853_));
 sky130_fd_sc_hd__a2bb2o_1 _1596_ (.A1_N(_0815_),
    .A2_N(_0846_),
    .B1(_0853_),
    .B2(_0845_),
    .X(_0854_));
 sky130_fd_sc_hd__buf_6 _1597_ (.A(_0605_),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _1598_ (.A0(net194),
    .A1(net53),
    .S(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__xnor2_1 _1599_ (.A(_0854_),
    .B(_0856_),
    .Y(net177));
 sky130_fd_sc_hd__or2_2 _1600_ (.A(net70),
    .B(_0691_),
    .X(_0857_));
 sky130_fd_sc_hd__or2_2 _1601_ (.A(net118),
    .B(_0822_),
    .X(_0858_));
 sky130_fd_sc_hd__a21o_1 _1602_ (.A1(_0857_),
    .A2(_0858_),
    .B1(_0709_),
    .X(_0859_));
 sky130_fd_sc_hd__clkbuf_4 _1603_ (.A(_0650_),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _1604_ (.A0(net117),
    .A1(net98),
    .S(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__o21a_1 _1605_ (.A1(_0727_),
    .A2(_0861_),
    .B1(_0729_),
    .X(_0862_));
 sky130_fd_sc_hd__clkbuf_4 _1606_ (.A(_0737_),
    .X(_0863_));
 sky130_fd_sc_hd__or2_2 _1607_ (.A(net67),
    .B(_0689_),
    .X(_0864_));
 sky130_fd_sc_hd__or2_2 _1608_ (.A(net93),
    .B(_0691_),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _1609_ (.A0(net114),
    .A1(net108),
    .S(_0659_),
    .X(_0866_));
 sky130_fd_sc_hd__a32o_1 _1610_ (.A1(_0863_),
    .A2(_0864_),
    .A3(_0865_),
    .B1(_0866_),
    .B2(_0716_),
    .X(_0867_));
 sky130_fd_sc_hd__or2_2 _1611_ (.A(net92),
    .B(_0770_),
    .X(_0868_));
 sky130_fd_sc_hd__or2_2 _1612_ (.A(net68),
    .B(_0761_),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _1613_ (.A0(net76),
    .A1(net83),
    .S(_0860_),
    .X(_0870_));
 sky130_fd_sc_hd__a32o_1 _1614_ (.A1(_0721_),
    .A2(_0868_),
    .A3(_0869_),
    .B1(_0870_),
    .B2(_0688_),
    .X(_0871_));
 sky130_fd_sc_hd__or2_2 _1615_ (.A(net82),
    .B(_0697_),
    .X(_0872_));
 sky130_fd_sc_hd__or2_2 _1616_ (.A(net78),
    .B(_0684_),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _1617_ (.A0(net107),
    .A1(net115),
    .S(_0860_),
    .X(_0874_));
 sky130_fd_sc_hd__a32o_1 _1618_ (.A1(_0657_),
    .A2(_0872_),
    .A3(_0873_),
    .B1(_0874_),
    .B2(_0674_),
    .X(_0875_));
 sky130_fd_sc_hd__or4_2 _1619_ (.A(_0862_),
    .B(_0867_),
    .C(_0871_),
    .D(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__nand3b_4 _1620_ (.A_N(net150),
    .B(_0859_),
    .C(_0876_),
    .Y(_0877_));
 sky130_fd_sc_hd__a21bo_2 _1621_ (.A1(_0859_),
    .A2(_0876_),
    .B1_N(net150),
    .X(_0878_));
 sky130_fd_sc_hd__or2_4 _1622_ (.A(net110),
    .B(_0650_),
    .X(_0879_));
 sky130_fd_sc_hd__or2_2 _1623_ (.A(net101),
    .B(_0689_),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _1624_ (.A0(net116),
    .A1(net107),
    .S(_0689_),
    .X(_0881_));
 sky130_fd_sc_hd__a32o_1 _1625_ (.A1(_0681_),
    .A2(_0879_),
    .A3(_0880_),
    .B1(_0881_),
    .B2(_0643_),
    .X(_0882_));
 sky130_fd_sc_hd__or2_2 _1626_ (.A(net70),
    .B(_0646_),
    .X(_0883_));
 sky130_fd_sc_hd__or2_2 _1627_ (.A(net91),
    .B(_0651_),
    .X(_0884_));
 sky130_fd_sc_hd__clkbuf_4 _1628_ (.A(net85),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _1629_ (.A0(_0885_),
    .A1(net75),
    .S(_0689_),
    .X(_0886_));
 sky130_fd_sc_hd__a32o_1 _1630_ (.A1(_0790_),
    .A2(_0883_),
    .A3(_0884_),
    .B1(_0886_),
    .B2(_0696_),
    .X(_0887_));
 sky130_fd_sc_hd__or2_4 _1631_ (.A(net69),
    .B(_0658_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _1632_ (.A0(net99),
    .A1(net67),
    .S(_0770_),
    .X(_0889_));
 sky130_fd_sc_hd__clkbuf_4 _1633_ (.A(_0672_),
    .X(_0890_));
 sky130_fd_sc_hd__a32o_1 _1634_ (.A1(_0773_),
    .A2(_0868_),
    .A3(_0888_),
    .B1(_0889_),
    .B2(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__clkbuf_4 _1635_ (.A(_0666_),
    .X(_0892_));
 sky130_fd_sc_hd__or2_2 _1636_ (.A(net106),
    .B(_0691_),
    .X(_0893_));
 sky130_fd_sc_hd__a31o_1 _1637_ (.A1(_0892_),
    .A2(_0872_),
    .A3(_0893_),
    .B1(_0693_),
    .X(_0894_));
 sky130_fd_sc_hd__or4_2 _1638_ (.A(_0882_),
    .B(_0887_),
    .C(_0891_),
    .D(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__or2_2 _1639_ (.A(net76),
    .B(_0822_),
    .X(_0896_));
 sky130_fd_sc_hd__or2_2 _1640_ (.A(net84),
    .B(_0770_),
    .X(_0897_));
 sky130_fd_sc_hd__a21o_1 _1641_ (.A1(_0896_),
    .A2(_0897_),
    .B1(_0779_),
    .X(_0898_));
 sky130_fd_sc_hd__nand3b_2 _1642_ (.A_N(net132),
    .B(_0895_),
    .C(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__a21bo_1 _1643_ (.A1(_0895_),
    .A2(_0898_),
    .B1_N(net132),
    .X(_0900_));
 sky130_fd_sc_hd__a22o_1 _1644_ (.A1(_0877_),
    .A2(_0878_),
    .B1(_0899_),
    .B2(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__nand4_4 _1645_ (.A(_0877_),
    .B(_0878_),
    .C(_0899_),
    .D(_0900_),
    .Y(_0902_));
 sky130_fd_sc_hd__inv_2 _1646_ (.A(net141),
    .Y(_0903_));
 sky130_fd_sc_hd__or2_2 _1647_ (.A(net114),
    .B(_0659_),
    .X(_0904_));
 sky130_fd_sc_hd__or2_4 _1648_ (.A(net99),
    .B(_0661_),
    .X(_0905_));
 sky130_fd_sc_hd__a21o_1 _1649_ (.A1(_0904_),
    .A2(_0905_),
    .B1(_0709_),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _1650_ (.A0(net110),
    .A1(_0885_),
    .S(_0659_),
    .X(_0907_));
 sky130_fd_sc_hd__o21a_1 _1651_ (.A1(_0727_),
    .A2(_0907_),
    .B1(_0729_),
    .X(_0908_));
 sky130_fd_sc_hd__or2_2 _1652_ (.A(net75),
    .B(_0670_),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _1653_ (.A0(net82),
    .A1(net91),
    .S(_0651_),
    .X(_0910_));
 sky130_fd_sc_hd__a32o_1 _1654_ (.A1(_0681_),
    .A2(_0857_),
    .A3(_0909_),
    .B1(_0910_),
    .B2(_0863_),
    .X(_0911_));
 sky130_fd_sc_hd__or2_2 _1655_ (.A(net92),
    .B(_0689_),
    .X(_0912_));
 sky130_fd_sc_hd__or2_2 _1656_ (.A(net116),
    .B(_0684_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _1657_ (.A0(net101),
    .A1(net107),
    .S(_0651_),
    .X(_0914_));
 sky130_fd_sc_hd__a32o_1 _1658_ (.A1(_0892_),
    .A2(_0912_),
    .A3(_0913_),
    .B1(_0914_),
    .B2(_0688_),
    .X(_0915_));
 sky130_fd_sc_hd__or2_2 _1659_ (.A(net69),
    .B(_0763_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _1660_ (.A0(net106),
    .A1(net67),
    .S(_0697_),
    .X(_0917_));
 sky130_fd_sc_hd__a32o_1 _1661_ (.A1(_0674_),
    .A2(_0896_),
    .A3(_0916_),
    .B1(_0917_),
    .B2(_0657_),
    .X(_0918_));
 sky130_fd_sc_hd__or4_4 _1662_ (.A(_0908_),
    .B(_0911_),
    .C(_0915_),
    .D(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__and3_2 _1663_ (.A(_0903_),
    .B(_0906_),
    .C(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__a21oi_4 _1664_ (.A1(_0906_),
    .A2(_0919_),
    .B1(_0903_),
    .Y(_0921_));
 sky130_fd_sc_hd__nor2_2 _1665_ (.A(_0920_),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__a21oi_1 _1666_ (.A1(_0901_),
    .A2(_0902_),
    .B1(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__or2_2 _1667_ (.A(net84),
    .B(_0658_),
    .X(_0924_));
 sky130_fd_sc_hd__or2_1 _1668_ (.A(net116),
    .B(_0753_),
    .X(_0925_));
 sky130_fd_sc_hd__o211a_1 _1669_ (.A1(net74),
    .A2(_0795_),
    .B1(_0834_),
    .C1(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__o211a_1 _1670_ (.A1(_0885_),
    .A2(_0838_),
    .B1(_0797_),
    .C1(_0873_),
    .X(_0927_));
 sky130_fd_sc_hd__a311o_1 _1671_ (.A1(_0682_),
    .A2(_0893_),
    .A3(_0924_),
    .B1(_0926_),
    .C1(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__or2_2 _1672_ (.A(net100),
    .B(_0761_),
    .X(_0929_));
 sky130_fd_sc_hd__or2_1 _1673_ (.A(net118),
    .B(_0770_),
    .X(_0930_));
 sky130_fd_sc_hd__and3_1 _1674_ (.A(_0721_),
    .B(_0880_),
    .C(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _1675_ (.A0(net75),
    .A1(net115),
    .S(_0702_),
    .X(_0932_));
 sky130_fd_sc_hd__a32o_1 _1676_ (.A1(_0799_),
    .A2(_0905_),
    .A3(_0888_),
    .B1(_0932_),
    .B2(_0839_),
    .X(_0933_));
 sky130_fd_sc_hd__a311o_1 _1677_ (.A1(_0832_),
    .A2(_0884_),
    .A3(_0929_),
    .B1(_0931_),
    .C1(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__or2_1 _1678_ (.A(net110),
    .B(_0822_),
    .X(_0935_));
 sky130_fd_sc_hd__or2_2 _1679_ (.A(net68),
    .B(_0770_),
    .X(_0936_));
 sky130_fd_sc_hd__and3_1 _1680_ (.A(_0751_),
    .B(_0935_),
    .C(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__or3_2 _1681_ (.A(_0928_),
    .B(_0934_),
    .C(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__xnor2_4 _1682_ (.A(net187),
    .B(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__buf_2 _1683_ (.A(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__and3b_1 _1684_ (.A_N(net132),
    .B(_0895_),
    .C(_0898_),
    .X(_0941_));
 sky130_fd_sc_hd__a21boi_1 _1685_ (.A1(_0895_),
    .A2(_0898_),
    .B1_N(net132),
    .Y(_0942_));
 sky130_fd_sc_hd__nor2_2 _1686_ (.A(_0941_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__buf_2 _1687_ (.A(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__nand2_1 _1688_ (.A(_0922_),
    .B(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__or3b_1 _1689_ (.A(_0923_),
    .B(_0940_),
    .C_N(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__inv_2 _1690_ (.A(_0939_),
    .Y(_0947_));
 sky130_fd_sc_hd__nor2_1 _1691_ (.A(_0922_),
    .B(_0944_),
    .Y(_0948_));
 sky130_fd_sc_hd__o211ai_4 _1692_ (.A1(_0920_),
    .A2(_0921_),
    .B1(_0877_),
    .C1(_0878_),
    .Y(_0949_));
 sky130_fd_sc_hd__a21boi_1 _1693_ (.A1(_0901_),
    .A2(_0902_),
    .B1_N(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__or3_1 _1694_ (.A(_0947_),
    .B(_0948_),
    .C(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__or2_2 _1695_ (.A(net93),
    .B(_0753_),
    .X(_0952_));
 sky130_fd_sc_hd__or2_2 _1696_ (.A(net101),
    .B(_0702_),
    .X(_0953_));
 sky130_fd_sc_hd__or2_2 _1697_ (.A(net98),
    .B(_0761_),
    .X(_0954_));
 sky130_fd_sc_hd__or2_2 _1698_ (.A(net76),
    .B(_0691_),
    .X(_0955_));
 sky130_fd_sc_hd__or2_2 _1699_ (.A(net108),
    .B(_0860_),
    .X(_0956_));
 sky130_fd_sc_hd__o211a_1 _1700_ (.A1(_0885_),
    .A2(_0838_),
    .B1(_0839_),
    .C1(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__a31o_1 _1701_ (.A1(_0826_),
    .A2(_0955_),
    .A3(_0872_),
    .B1(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__or2_2 _1702_ (.A(net117),
    .B(_0795_),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _1703_ (.A0(net75),
    .A1(net83),
    .S(_0702_),
    .X(_0960_));
 sky130_fd_sc_hd__a32o_1 _1704_ (.A1(_0799_),
    .A2(_0868_),
    .A3(_0864_),
    .B1(_0797_),
    .B2(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__or2_2 _1705_ (.A(net107),
    .B(_0650_),
    .X(_0962_));
 sky130_fd_sc_hd__and3_1 _1706_ (.A(_0834_),
    .B(_0962_),
    .C(_0904_),
    .X(_0963_));
 sky130_fd_sc_hd__a311o_1 _1707_ (.A1(_0832_),
    .A2(_0883_),
    .A3(_0959_),
    .B1(_0961_),
    .C1(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__a311o_1 _1708_ (.A1(_0821_),
    .A2(_0954_),
    .A3(_0879_),
    .B1(_0958_),
    .C1(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__a31oi_4 _1709_ (.A1(_0819_),
    .A2(_0952_),
    .A3(_0953_),
    .B1(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__xnor2_4 _1710_ (.A(net158),
    .B(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__inv_2 _1711_ (.A(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__a21oi_1 _1712_ (.A1(_0946_),
    .A2(_0951_),
    .B1(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__or2_2 _1713_ (.A(net115),
    .B(_0860_),
    .X(_0970_));
 sky130_fd_sc_hd__or2_2 _1714_ (.A(net83),
    .B(_0770_),
    .X(_0971_));
 sky130_fd_sc_hd__o211a_1 _1715_ (.A1(net117),
    .A2(_0838_),
    .B1(_0826_),
    .C1(_0971_),
    .X(_0972_));
 sky130_fd_sc_hd__or2_2 _1716_ (.A(net78),
    .B(_0753_),
    .X(_0973_));
 sky130_fd_sc_hd__o211a_1 _1717_ (.A1(net67),
    .A2(_0796_),
    .B1(_0821_),
    .C1(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__a311o_1 _1718_ (.A1(_0840_),
    .A2(_0912_),
    .A3(_0970_),
    .B1(_0972_),
    .C1(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__or2_1 _1719_ (.A(net82),
    .B(_0795_),
    .X(_0976_));
 sky130_fd_sc_hd__and3_1 _1720_ (.A(_0825_),
    .B(_0976_),
    .C(_0858_),
    .X(_0977_));
 sky130_fd_sc_hd__or2_2 _1721_ (.A(net108),
    .B(_0822_),
    .X(_0978_));
 sky130_fd_sc_hd__or2_2 _1722_ (.A(net98),
    .B(_0763_),
    .X(_0979_));
 sky130_fd_sc_hd__and3_1 _1723_ (.A(_0829_),
    .B(_0978_),
    .C(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__clkbuf_4 _1724_ (.A(_0688_),
    .X(_0981_));
 sky130_fd_sc_hd__or2_2 _1725_ (.A(net114),
    .B(_0763_),
    .X(_0982_));
 sky130_fd_sc_hd__and3_1 _1726_ (.A(_0981_),
    .B(_0952_),
    .C(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__and3_1 _1727_ (.A(_0832_),
    .B(_0896_),
    .C(_0936_),
    .X(_0984_));
 sky130_fd_sc_hd__or4_1 _1728_ (.A(_0977_),
    .B(_0980_),
    .C(_0983_),
    .D(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__and3_1 _1729_ (.A(_0819_),
    .B(_0962_),
    .C(_0929_),
    .X(_0986_));
 sky130_fd_sc_hd__nor3_2 _1730_ (.A(_0975_),
    .B(_0985_),
    .C(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__xnor2_2 _1731_ (.A(net178),
    .B(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__inv_2 _1732_ (.A(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__a211o_2 _1733_ (.A1(_0877_),
    .A2(_0878_),
    .B1(_0920_),
    .C1(_0921_),
    .X(_0990_));
 sky130_fd_sc_hd__nor2b_2 _1734_ (.A(_0939_),
    .B_N(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__a21o_2 _1735_ (.A1(_0949_),
    .A2(_0990_),
    .B1(_0944_),
    .X(_0992_));
 sky130_fd_sc_hd__nand2_1 _1736_ (.A(_0944_),
    .B(_0990_),
    .Y(_0993_));
 sky130_fd_sc_hd__and3_1 _1737_ (.A(_0940_),
    .B(_0992_),
    .C(_0993_),
    .X(_0994_));
 sky130_fd_sc_hd__a211oi_1 _1738_ (.A1(_0901_),
    .A2(_0991_),
    .B1(_0994_),
    .C1(_0967_),
    .Y(_0995_));
 sky130_fd_sc_hd__or3_2 _1739_ (.A(_0922_),
    .B(_0941_),
    .C(_0942_),
    .X(_0996_));
 sky130_fd_sc_hd__a21oi_1 _1740_ (.A1(_0992_),
    .A2(_0996_),
    .B1(_0991_),
    .Y(_0997_));
 sky130_fd_sc_hd__a31o_1 _1741_ (.A1(_0992_),
    .A2(_0991_),
    .A3(_0996_),
    .B1(_0967_),
    .X(_0998_));
 sky130_fd_sc_hd__nor2_1 _1742_ (.A(_0997_),
    .B(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__and2b_1 _1743_ (.A_N(_0943_),
    .B(_0922_),
    .X(_1000_));
 sky130_fd_sc_hd__a311o_1 _1744_ (.A1(_0944_),
    .A2(_0949_),
    .A3(_0990_),
    .B1(_1000_),
    .C1(_0947_),
    .X(_1001_));
 sky130_fd_sc_hd__a31o_1 _1745_ (.A1(_0967_),
    .A2(_0946_),
    .A3(_1001_),
    .B1(_0988_),
    .X(_1002_));
 sky130_fd_sc_hd__o32a_2 _1746_ (.A1(_0969_),
    .A2(_0989_),
    .A3(_0995_),
    .B1(_0999_),
    .B2(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _1747_ (.A0(\L[31] ),
    .A1(net44),
    .S(_0855_),
    .X(_1004_));
 sky130_fd_sc_hd__xnor2_2 _1748_ (.A(_1003_),
    .B(_1004_),
    .Y(net168));
 sky130_fd_sc_hd__or2_2 _1749_ (.A(net106),
    .B(_0689_),
    .X(_1005_));
 sky130_fd_sc_hd__and3_1 _1750_ (.A(_0839_),
    .B(_0954_),
    .C(_0905_),
    .X(_1006_));
 sky130_fd_sc_hd__and3_1 _1751_ (.A(_0834_),
    .B(_0865_),
    .C(_0929_),
    .X(_1007_));
 sky130_fd_sc_hd__a311o_1 _1752_ (.A1(_0825_),
    .A2(_0959_),
    .A3(_0888_),
    .B1(_1006_),
    .C1(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__or2_2 _1753_ (.A(net83),
    .B(_0822_),
    .X(_1009_));
 sky130_fd_sc_hd__o211a_1 _1754_ (.A1(net74),
    .A2(_0796_),
    .B1(_1009_),
    .C1(_0644_),
    .X(_1010_));
 sky130_fd_sc_hd__a31o_1 _1755_ (.A1(_0826_),
    .A2(_0869_),
    .A3(_0930_),
    .B1(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__or2_2 _1756_ (.A(net115),
    .B(_0761_),
    .X(_1012_));
 sky130_fd_sc_hd__and3_1 _1757_ (.A(_0829_),
    .B(_0873_),
    .C(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__and3_1 _1758_ (.A(_0821_),
    .B(_0956_),
    .C(_0924_),
    .X(_1014_));
 sky130_fd_sc_hd__or4_1 _1759_ (.A(_1008_),
    .B(_1011_),
    .C(_1013_),
    .D(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__a31o_1 _1760_ (.A1(_0819_),
    .A2(_1005_),
    .A3(_0982_),
    .B1(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__xor2_4 _1761_ (.A(net185),
    .B(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__inv_2 _1762_ (.A(_1017_),
    .Y(_1018_));
 sky130_fd_sc_hd__or2_2 _1763_ (.A(net100),
    .B(_0860_),
    .X(_1019_));
 sky130_fd_sc_hd__and3_1 _1764_ (.A(_0773_),
    .B(_0916_),
    .C(_0978_),
    .X(_1020_));
 sky130_fd_sc_hd__or2_2 _1765_ (.A(net74),
    .B(_0761_),
    .X(_1021_));
 sky130_fd_sc_hd__and3_1 _1766_ (.A(_0790_),
    .B(_0936_),
    .C(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__a311o_1 _1767_ (.A1(_0716_),
    .A2(_0973_),
    .A3(_1019_),
    .B1(_1020_),
    .C1(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__and3_1 _1768_ (.A(_0797_),
    .B(_1005_),
    .C(_0979_),
    .X(_1024_));
 sky130_fd_sc_hd__and3_1 _1769_ (.A(_0799_),
    .B(_0858_),
    .C(_0970_),
    .X(_1025_));
 sky130_fd_sc_hd__or2_1 _1770_ (.A(net99),
    .B(_0697_),
    .X(_1026_));
 sky130_fd_sc_hd__and3_1 _1771_ (.A(_0892_),
    .B(_0971_),
    .C(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__a31o_1 _1772_ (.A1(_0644_),
    .A2(_0952_),
    .A3(_0897_),
    .B1(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__or4_1 _1773_ (.A(_1023_),
    .B(_1024_),
    .C(_1025_),
    .D(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__a31o_1 _1774_ (.A1(_0788_),
    .A2(_0959_),
    .A3(_0925_),
    .B1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__xor2_2 _1775_ (.A(net156),
    .B(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__inv_2 _1776_ (.A(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__o21a_1 _1777_ (.A1(net74),
    .A2(_0795_),
    .B1(_0864_),
    .X(_1033_));
 sky130_fd_sc_hd__or2_2 _1778_ (.A(_0779_),
    .B(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__mux2_1 _1779_ (.A0(net101),
    .A1(net75),
    .S(_0651_),
    .X(_1035_));
 sky130_fd_sc_hd__o21a_1 _1780_ (.A1(_0727_),
    .A2(_1035_),
    .B1(_0729_),
    .X(_1036_));
 sky130_fd_sc_hd__mux2_1 _1781_ (.A0(net99),
    .A1(net82),
    .S(_0689_),
    .X(_1037_));
 sky130_fd_sc_hd__a32o_1 _1782_ (.A1(_0890_),
    .A2(_0912_),
    .A3(_0897_),
    .B1(_1037_),
    .B2(_0773_),
    .X(_1038_));
 sky130_fd_sc_hd__or2_2 _1783_ (.A(net107),
    .B(_0697_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _1784_ (.A0(net116),
    .A1(net110),
    .S(_0770_),
    .X(_1040_));
 sky130_fd_sc_hd__a32o_1 _1785_ (.A1(_0892_),
    .A2(_1039_),
    .A3(_0916_),
    .B1(_1040_),
    .B2(_0790_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _1786_ (.A0(_0885_),
    .A1(net91),
    .S(_0770_),
    .X(_1042_));
 sky130_fd_sc_hd__a32o_1 _1787_ (.A1(_0643_),
    .A2(_1005_),
    .A3(_0857_),
    .B1(_1042_),
    .B2(_0681_),
    .X(_1043_));
 sky130_fd_sc_hd__or4_2 _1788_ (.A(_1036_),
    .B(_1038_),
    .C(_1041_),
    .D(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__nand3_2 _1789_ (.A(_0627_),
    .B(_1034_),
    .C(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a21o_1 _1790_ (.A1(_1034_),
    .A2(_1044_),
    .B1(_0627_),
    .X(_1046_));
 sky130_fd_sc_hd__o21a_1 _1791_ (.A1(_0885_),
    .A2(_0838_),
    .B1(_0865_),
    .X(_1047_));
 sky130_fd_sc_hd__or2_1 _1792_ (.A(_0779_),
    .B(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_1 _1793_ (.A0(net99),
    .A1(net84),
    .S(_0659_),
    .X(_1049_));
 sky130_fd_sc_hd__o21a_1 _1794_ (.A1(_0727_),
    .A2(_1049_),
    .B1(_0729_),
    .X(_1050_));
 sky130_fd_sc_hd__mux2_1 _1795_ (.A0(net101),
    .A1(net78),
    .S(_0651_),
    .X(_1051_));
 sky130_fd_sc_hd__a32o_1 _1796_ (.A1(_0890_),
    .A2(_0909_),
    .A3(_0936_),
    .B1(_1051_),
    .B2(_0657_),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _1797_ (.A0(net91),
    .A1(net115),
    .S(_0697_),
    .X(_1053_));
 sky130_fd_sc_hd__a32o_1 _1798_ (.A1(_0790_),
    .A2(_1005_),
    .A3(_1019_),
    .B1(_1053_),
    .B2(_0721_),
    .X(_1054_));
 sky130_fd_sc_hd__mux2_1 _1799_ (.A0(net116),
    .A1(net118),
    .S(_0684_),
    .X(_1055_));
 sky130_fd_sc_hd__a32o_1 _1800_ (.A1(_0681_),
    .A2(_0916_),
    .A3(_1021_),
    .B1(_1055_),
    .B2(_0863_),
    .X(_1056_));
 sky130_fd_sc_hd__or4_1 _1801_ (.A(_1050_),
    .B(_1052_),
    .C(_1054_),
    .D(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__and3b_2 _1802_ (.A_N(net139),
    .B(_1048_),
    .C(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__a21boi_2 _1803_ (.A1(_1048_),
    .A2(_1057_),
    .B1_N(net139),
    .Y(_1059_));
 sky130_fd_sc_hd__a211o_2 _1804_ (.A1(_1045_),
    .A2(_1046_),
    .B1(_1058_),
    .C1(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__o211ai_4 _1805_ (.A1(_1058_),
    .A2(_1059_),
    .B1(_1045_),
    .C1(_1046_),
    .Y(_1061_));
 sky130_fd_sc_hd__nand2_1 _1806_ (.A(_1060_),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__and3_1 _1807_ (.A(_0892_),
    .B(_0858_),
    .C(_0982_),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _1808_ (.A0(net67),
    .A1(net74),
    .S(_0684_),
    .X(_1064_));
 sky130_fd_sc_hd__a32o_1 _1809_ (.A1(_0657_),
    .A2(_0896_),
    .A3(_1019_),
    .B1(_1064_),
    .B2(_0674_),
    .X(_1065_));
 sky130_fd_sc_hd__a311o_1 _1810_ (.A1(_0834_),
    .A2(_0973_),
    .A3(_0979_),
    .B1(_1063_),
    .C1(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__a21o_1 _1811_ (.A1(_0952_),
    .A2(_0971_),
    .B1(_0727_),
    .X(_1067_));
 sky130_fd_sc_hd__o211a_1 _1812_ (.A1(net117),
    .A2(_0753_),
    .B1(_0970_),
    .C1(_0863_),
    .X(_1068_));
 sky130_fd_sc_hd__and3_1 _1813_ (.A(_0716_),
    .B(_0936_),
    .C(_0978_),
    .X(_1069_));
 sky130_fd_sc_hd__a211o_1 _1814_ (.A1(_0729_),
    .A2(_1067_),
    .B1(_1068_),
    .C1(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__a21o_1 _1815_ (.A1(_0868_),
    .A2(_0924_),
    .B1(_0709_),
    .X(_1071_));
 sky130_fd_sc_hd__o21ai_4 _1816_ (.A1(_1066_),
    .A2(_1070_),
    .B1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__xnor2_4 _1817_ (.A(net130),
    .B(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__nor2_2 _1818_ (.A(_1058_),
    .B(_1059_),
    .Y(_1074_));
 sky130_fd_sc_hd__or2_1 _1819_ (.A(_1073_),
    .B(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__and3_1 _1820_ (.A(_0674_),
    .B(_0865_),
    .C(_0880_),
    .X(_1076_));
 sky130_fd_sc_hd__and3_1 _1821_ (.A(_0688_),
    .B(_0888_),
    .C(_0930_),
    .X(_1077_));
 sky130_fd_sc_hd__a311o_1 _1822_ (.A1(_0682_),
    .A2(_0905_),
    .A3(_0929_),
    .B1(_1076_),
    .C1(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__o211a_1 _1823_ (.A1(net74),
    .A2(_0795_),
    .B1(_0696_),
    .C1(_0924_),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _1824_ (.A0(net116),
    .A1(net78),
    .S(_0659_),
    .X(_1080_));
 sky130_fd_sc_hd__a32o_1 _1825_ (.A1(_0863_),
    .A2(_1012_),
    .A3(_0893_),
    .B1(_1080_),
    .B2(_0721_),
    .X(_1081_));
 sky130_fd_sc_hd__a311o_1 _1826_ (.A1(_0839_),
    .A2(_0869_),
    .A3(_0884_),
    .B1(_1079_),
    .C1(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__and3_1 _1827_ (.A(_0751_),
    .B(_0909_),
    .C(_0971_),
    .X(_1083_));
 sky130_fd_sc_hd__or3_2 _1828_ (.A(_1078_),
    .B(_1082_),
    .C(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__xnor2_4 _1829_ (.A(net181),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__inv_2 _1830_ (.A(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__a21o_1 _1831_ (.A1(_1062_),
    .A2(_1075_),
    .B1(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__xor2_2 _1832_ (.A(net130),
    .B(_1072_),
    .X(_1088_));
 sky130_fd_sc_hd__and3_1 _1833_ (.A(_0627_),
    .B(_1034_),
    .C(_1044_),
    .X(_1089_));
 sky130_fd_sc_hd__a21oi_1 _1834_ (.A1(_1034_),
    .A2(_1044_),
    .B1(_0627_),
    .Y(_1090_));
 sky130_fd_sc_hd__nor2_2 _1835_ (.A(_1089_),
    .B(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__xnor2_2 _1836_ (.A(_1088_),
    .B(_1091_),
    .Y(_1092_));
 sky130_fd_sc_hd__or3b_1 _1837_ (.A(_1092_),
    .B(_1085_),
    .C_N(_1061_),
    .X(_1093_));
 sky130_fd_sc_hd__and3_1 _1838_ (.A(_1032_),
    .B(_1087_),
    .C(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__buf_2 _1839_ (.A(_1088_),
    .X(_1095_));
 sky130_fd_sc_hd__nor2_1 _1840_ (.A(_1095_),
    .B(_1062_),
    .Y(_1096_));
 sky130_fd_sc_hd__o211a_1 _1841_ (.A1(_1089_),
    .A2(_1090_),
    .B1(_1095_),
    .C1(_1074_),
    .X(_1097_));
 sky130_fd_sc_hd__buf_2 _1842_ (.A(_1085_),
    .X(_1098_));
 sky130_fd_sc_hd__nor2_1 _1843_ (.A(_1074_),
    .B(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__or4_1 _1844_ (.A(_1095_),
    .B(_1074_),
    .C(_1091_),
    .D(_1085_),
    .X(_1100_));
 sky130_fd_sc_hd__buf_2 _1845_ (.A(_1031_),
    .X(_1101_));
 sky130_fd_sc_hd__o311a_1 _1846_ (.A1(_1096_),
    .A2(_1097_),
    .A3(_1099_),
    .B1(_1100_),
    .C1(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__nand2_1 _1847_ (.A(_1074_),
    .B(_1098_),
    .Y(_1103_));
 sky130_fd_sc_hd__a211o_1 _1848_ (.A1(_1092_),
    .A2(_1103_),
    .B1(_1097_),
    .C1(_1101_),
    .X(_1104_));
 sky130_fd_sc_hd__nand2_1 _1849_ (.A(_1018_),
    .B(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__or2_1 _1850_ (.A(_1095_),
    .B(_1060_),
    .X(_1106_));
 sky130_fd_sc_hd__nand2_1 _1851_ (.A(_1095_),
    .B(_1060_),
    .Y(_1107_));
 sky130_fd_sc_hd__and3_1 _1852_ (.A(_1106_),
    .B(_1098_),
    .C(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__nand3_2 _1853_ (.A(_1073_),
    .B(_1060_),
    .C(_1061_),
    .Y(_1109_));
 sky130_fd_sc_hd__a21o_1 _1854_ (.A1(_1060_),
    .A2(_1061_),
    .B1(_1073_),
    .X(_1110_));
 sky130_fd_sc_hd__and3_1 _1855_ (.A(_1086_),
    .B(_1109_),
    .C(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__o21a_1 _1856_ (.A1(_1108_),
    .A2(_1111_),
    .B1(_1101_),
    .X(_1112_));
 sky130_fd_sc_hd__o32a_4 _1857_ (.A1(_1018_),
    .A2(_1094_),
    .A3(_1102_),
    .B1(_1105_),
    .B2(_1112_),
    .X(_1113_));
 sky130_fd_sc_hd__clkbuf_8 _1858_ (.A(_0605_),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_2 _1859_ (.A0(\L[30] ),
    .A1(net36),
    .S(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__xor2_4 _1860_ (.A(_1113_),
    .B(_1115_),
    .X(net160));
 sky130_fd_sc_hd__or2_2 _1861_ (.A(net119),
    .B(_0670_),
    .X(_1116_));
 sky130_fd_sc_hd__o211a_1 _1862_ (.A1(net95),
    .A2(_0796_),
    .B1(_0821_),
    .C1(_0719_),
    .X(_1117_));
 sky130_fd_sc_hd__or2_1 _1863_ (.A(net109),
    .B(_0650_),
    .X(_1118_));
 sky130_fd_sc_hd__and3_1 _1864_ (.A(_0826_),
    .B(_0713_),
    .C(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__nor2_1 _1865_ (.A(net66),
    .B(_0753_),
    .Y(_1120_));
 sky130_fd_sc_hd__and3b_1 _1866_ (.A_N(_1120_),
    .B(_0714_),
    .C(_0840_),
    .X(_1121_));
 sky130_fd_sc_hd__or2_2 _1867_ (.A(net111),
    .B(_0860_),
    .X(_1122_));
 sky130_fd_sc_hd__or2_2 _1868_ (.A(net88),
    .B(_0753_),
    .X(_1123_));
 sky130_fd_sc_hd__and3_1 _1869_ (.A(_0799_),
    .B(_0718_),
    .C(_0767_),
    .X(_1124_));
 sky130_fd_sc_hd__a31o_1 _1870_ (.A1(_0797_),
    .A2(_1122_),
    .A3(_1123_),
    .B1(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__o211a_1 _1871_ (.A1(net94),
    .A2(_0796_),
    .B1(_0723_),
    .C1(_0832_),
    .X(_1126_));
 sky130_fd_sc_hd__a311o_1 _1872_ (.A1(_0981_),
    .A2(_0704_),
    .A3(_0752_),
    .B1(_1125_),
    .C1(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__or4_2 _1873_ (.A(_1117_),
    .B(_1119_),
    .C(_1121_),
    .D(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__a31oi_4 _1874_ (.A1(_0819_),
    .A2(_0692_),
    .A3(_1116_),
    .B1(_1128_),
    .Y(_1129_));
 sky130_fd_sc_hd__xor2_4 _1875_ (.A(net145),
    .B(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__and3_1 _1876_ (.A(_0863_),
    .B(_0660_),
    .C(_0685_),
    .X(_1131_));
 sky130_fd_sc_hd__a31o_1 _1877_ (.A1(_0648_),
    .A2(_0699_),
    .A3(_0682_),
    .B1(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__a21o_1 _1878_ (.A1(_0683_),
    .A2(_0692_),
    .B1(_0727_),
    .X(_1133_));
 sky130_fd_sc_hd__mux2_1 _1879_ (.A0(net120),
    .A1(net77),
    .S(_0689_),
    .X(_1134_));
 sky130_fd_sc_hd__a32o_1 _1880_ (.A1(_0652_),
    .A2(_0773_),
    .A3(_0801_),
    .B1(_1134_),
    .B2(_0890_),
    .X(_1135_));
 sky130_fd_sc_hd__and3_1 _1881_ (.A(_0892_),
    .B(_0676_),
    .C(_0690_),
    .X(_1136_));
 sky130_fd_sc_hd__and3_1 _1882_ (.A(_0698_),
    .B(_0669_),
    .C(_0790_),
    .X(_1137_));
 sky130_fd_sc_hd__a2111o_1 _1883_ (.A1(_0729_),
    .A2(_1133_),
    .B1(_1135_),
    .C1(_1136_),
    .D1(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__a21o_1 _1884_ (.A1(_0767_),
    .A2(_0831_),
    .B1(_0779_),
    .X(_1139_));
 sky130_fd_sc_hd__o21ai_2 _1885_ (.A1(_1132_),
    .A2(_1138_),
    .B1(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__xnor2_2 _1886_ (.A(net163),
    .B(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__o21a_1 _1887_ (.A1(net94),
    .A2(_0795_),
    .B1(_0823_),
    .X(_1142_));
 sky130_fd_sc_hd__or2_2 _1888_ (.A(_0709_),
    .B(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _1889_ (.A0(net81),
    .A1(net73),
    .S(_0659_),
    .X(_1144_));
 sky130_fd_sc_hd__a32o_1 _1890_ (.A1(_0657_),
    .A2(_0676_),
    .A3(_0740_),
    .B1(_1144_),
    .B2(_0674_),
    .X(_1145_));
 sky130_fd_sc_hd__mux2_1 _1891_ (.A0(net88),
    .A1(net96),
    .S(_0684_),
    .X(_1146_));
 sky130_fd_sc_hd__a32o_1 _1892_ (.A1(_0688_),
    .A2(_0738_),
    .A3(_0792_),
    .B1(_1146_),
    .B2(_0721_),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_1 _1893_ (.A0(net72),
    .A1(net113),
    .S(_0684_),
    .X(_1148_));
 sky130_fd_sc_hd__a32o_1 _1894_ (.A1(_0643_),
    .A2(_1116_),
    .A3(_0802_),
    .B1(_1148_),
    .B2(_0716_),
    .X(_1149_));
 sky130_fd_sc_hd__mux2_1 _1895_ (.A0(net97),
    .A1(net87),
    .S(_0659_),
    .X(_1150_));
 sky130_fd_sc_hd__o21a_1 _1896_ (.A1(_0727_),
    .A2(_1150_),
    .B1(_0729_),
    .X(_1151_));
 sky130_fd_sc_hd__or4_2 _1897_ (.A(_1145_),
    .B(_1147_),
    .C(_1149_),
    .D(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__nand3_4 _1898_ (.A(net180),
    .B(_1143_),
    .C(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__a21o_2 _1899_ (.A1(_1143_),
    .A2(_1152_),
    .B1(net180),
    .X(_1154_));
 sky130_fd_sc_hd__a21o_1 _1900_ (.A1(_0766_),
    .A2(_1123_),
    .B1(_0709_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _1901_ (.A0(net111),
    .A1(net73),
    .S(_0659_),
    .X(_1156_));
 sky130_fd_sc_hd__a32o_1 _1902_ (.A1(_0674_),
    .A2(_0692_),
    .A3(_0740_),
    .B1(_1156_),
    .B2(_0657_),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _1903_ (.A0(net105),
    .A1(net109),
    .S(_0860_),
    .X(_1158_));
 sky130_fd_sc_hd__a32o_1 _1904_ (.A1(_0699_),
    .A2(_0721_),
    .A3(_0778_),
    .B1(_1158_),
    .B2(_0688_),
    .X(_1159_));
 sky130_fd_sc_hd__mux2_1 _1905_ (.A0(net89),
    .A1(net95),
    .S(_0684_),
    .X(_1160_));
 sky130_fd_sc_hd__a32o_1 _1906_ (.A1(_0662_),
    .A2(_0716_),
    .A3(_0690_),
    .B1(_1160_),
    .B2(_0863_),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_1 _1907_ (.A0(net90),
    .A1(net120),
    .S(_0860_),
    .X(_1162_));
 sky130_fd_sc_hd__o21a_1 _1908_ (.A1(_0727_),
    .A2(_1162_),
    .B1(_0729_),
    .X(_1163_));
 sky130_fd_sc_hd__or4_2 _1909_ (.A(_1157_),
    .B(_1159_),
    .C(_1161_),
    .D(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__nand3b_4 _1910_ (.A_N(net172),
    .B(_1155_),
    .C(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__a21bo_2 _1911_ (.A1(_1155_),
    .A2(_1164_),
    .B1_N(net172),
    .X(_1166_));
 sky130_fd_sc_hd__a22o_2 _1912_ (.A1(_1153_),
    .A2(_1154_),
    .B1(_1165_),
    .B2(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__nand4_4 _1913_ (.A(_1153_),
    .B(_1154_),
    .C(_1165_),
    .D(_1166_),
    .Y(_1168_));
 sky130_fd_sc_hd__a21o_1 _1914_ (.A1(_1167_),
    .A2(_1168_),
    .B1(_1141_),
    .X(_1169_));
 sky130_fd_sc_hd__a21bo_1 _1915_ (.A1(_1141_),
    .A2(_1167_),
    .B1_N(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__and3_1 _1916_ (.A(_0834_),
    .B(_0724_),
    .C(_0754_),
    .X(_1171_));
 sky130_fd_sc_hd__and3_1 _1917_ (.A(_0839_),
    .B(_0703_),
    .C(_0719_),
    .X(_1172_));
 sky130_fd_sc_hd__a311o_1 _1918_ (.A1(_0832_),
    .A2(_1123_),
    .A3(_0831_),
    .B1(_1171_),
    .C1(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__mux2_1 _1919_ (.A0(net94),
    .A1(net102),
    .S(_0702_),
    .X(_1174_));
 sky130_fd_sc_hd__a32o_1 _1920_ (.A1(_0799_),
    .A2(_0824_),
    .A3(_0833_),
    .B1(_1174_),
    .B2(_0797_),
    .X(_1175_));
 sky130_fd_sc_hd__o211a_1 _1921_ (.A1(net103),
    .A2(_0838_),
    .B1(_0682_),
    .C1(_0789_),
    .X(_1176_));
 sky130_fd_sc_hd__a311o_1 _1922_ (.A1(_0821_),
    .A2(_0714_),
    .A3(_0830_),
    .B1(_1175_),
    .C1(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__or2_1 _1923_ (.A(net89),
    .B(_0691_),
    .X(_1178_));
 sky130_fd_sc_hd__and3_1 _1924_ (.A(_0660_),
    .B(_0788_),
    .C(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__or3_1 _1925_ (.A(_1173_),
    .B(_1177_),
    .C(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__xor2_1 _1926_ (.A(net137),
    .B(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__buf_2 _1927_ (.A(_1181_),
    .X(_1182_));
 sky130_fd_sc_hd__and3_1 _1928_ (.A(_0863_),
    .B(_1122_),
    .C(_0830_),
    .X(_1183_));
 sky130_fd_sc_hd__and3_1 _1929_ (.A(_0688_),
    .B(_0703_),
    .C(_0762_),
    .X(_1184_));
 sky130_fd_sc_hd__a311o_1 _1930_ (.A1(_0829_),
    .A2(_0823_),
    .A3(_0771_),
    .B1(_1183_),
    .C1(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__o211a_1 _1931_ (.A1(net95),
    .A2(_0795_),
    .B1(_0657_),
    .C1(_0754_),
    .X(_1186_));
 sky130_fd_sc_hd__and3b_1 _1932_ (.A_N(_1120_),
    .B(_0831_),
    .C(_0892_),
    .X(_1187_));
 sky130_fd_sc_hd__and3_1 _1933_ (.A(_0681_),
    .B(_0766_),
    .C(_0835_),
    .X(_1188_));
 sky130_fd_sc_hd__and3_1 _1934_ (.A(_0890_),
    .B(_0723_),
    .C(_0789_),
    .X(_1189_));
 sky130_fd_sc_hd__or4_2 _1935_ (.A(_1186_),
    .B(_1187_),
    .C(_1188_),
    .D(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__and3_1 _1936_ (.A(_0751_),
    .B(_0690_),
    .C(_0746_),
    .X(_1191_));
 sky130_fd_sc_hd__nor3_4 _1937_ (.A(_1185_),
    .B(_1190_),
    .C(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__xnor2_1 _1938_ (.A(net154),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__buf_2 _1939_ (.A(_1193_),
    .X(_1194_));
 sky130_fd_sc_hd__nand2_4 _1940_ (.A(_1165_),
    .B(_1166_),
    .Y(_1195_));
 sky130_fd_sc_hd__xor2_4 _1941_ (.A(net154),
    .B(_1192_),
    .X(_1196_));
 sky130_fd_sc_hd__o21ba_1 _1942_ (.A1(_1195_),
    .A2(_1196_),
    .B1_N(_1181_),
    .X(_1197_));
 sky130_fd_sc_hd__a31o_1 _1943_ (.A1(_1167_),
    .A2(_1182_),
    .A3(_1194_),
    .B1(_1197_),
    .X(_1198_));
 sky130_fd_sc_hd__xnor2_1 _1944_ (.A(_1170_),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__nand3_1 _1945_ (.A(_1141_),
    .B(_1167_),
    .C(_1168_),
    .Y(_1200_));
 sky130_fd_sc_hd__and3_1 _1946_ (.A(_1169_),
    .B(_1196_),
    .C(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__xor2_1 _1947_ (.A(net163),
    .B(_1140_),
    .X(_1202_));
 sky130_fd_sc_hd__clkbuf_4 _1948_ (.A(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__and2_1 _1949_ (.A(_1167_),
    .B(_1168_),
    .X(_1204_));
 sky130_fd_sc_hd__nand2_4 _1950_ (.A(_1153_),
    .B(_1154_),
    .Y(_1205_));
 sky130_fd_sc_hd__nand2_1 _1951_ (.A(_1203_),
    .B(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__o211a_1 _1952_ (.A1(_1203_),
    .A2(_1204_),
    .B1(_1194_),
    .C1(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__o21ai_1 _1953_ (.A1(_1201_),
    .A2(_1207_),
    .B1(_1182_),
    .Y(_1208_));
 sky130_fd_sc_hd__xnor2_1 _1954_ (.A(_1203_),
    .B(_1205_),
    .Y(_1209_));
 sky130_fd_sc_hd__nand2_1 _1955_ (.A(_1167_),
    .B(_1196_),
    .Y(_1210_));
 sky130_fd_sc_hd__nor2_1 _1956_ (.A(_1141_),
    .B(_1205_),
    .Y(_1211_));
 sky130_fd_sc_hd__inv_2 _1957_ (.A(_1181_),
    .Y(_1212_));
 sky130_fd_sc_hd__o221a_1 _1958_ (.A1(_1196_),
    .A2(_1209_),
    .B1(_1210_),
    .B2(_1211_),
    .C1(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__nor2_1 _1959_ (.A(_1130_),
    .B(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__a22o_1 _1960_ (.A1(_1130_),
    .A2(_1199_),
    .B1(_1208_),
    .B2(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__mux2_1 _1961_ (.A0(net195),
    .A1(net27),
    .S(_0855_),
    .X(_1216_));
 sky130_fd_sc_hd__xnor2_2 _1962_ (.A(_1215_),
    .B(_1216_),
    .Y(net151));
 sky130_fd_sc_hd__mux2_1 _1963_ (.A0(net116),
    .A1(net108),
    .S(_0822_),
    .X(_1217_));
 sky130_fd_sc_hd__a32o_1 _1964_ (.A1(_0773_),
    .A2(_1009_),
    .A3(_0893_),
    .B1(_1217_),
    .B2(_0890_),
    .X(_1218_));
 sky130_fd_sc_hd__mux2_1 _1965_ (.A0(net84),
    .A1(net78),
    .S(_0822_),
    .X(_1219_));
 sky130_fd_sc_hd__a32o_1 _1966_ (.A1(_0892_),
    .A2(_0865_),
    .A3(_0888_),
    .B1(_1219_),
    .B2(_0790_),
    .X(_1220_));
 sky130_fd_sc_hd__mux2_1 _1967_ (.A0(net115),
    .A1(net74),
    .S(_0822_),
    .X(_1221_));
 sky130_fd_sc_hd__a32o_1 _1968_ (.A1(_0737_),
    .A2(_0905_),
    .A3(_0869_),
    .B1(_1221_),
    .B2(_0681_),
    .X(_1222_));
 sky130_fd_sc_hd__mux2_1 _1969_ (.A0(net118),
    .A1(net100),
    .S(_0691_),
    .X(_1223_));
 sky130_fd_sc_hd__o21a_1 _1970_ (.A1(_0707_),
    .A2(_1223_),
    .B1(_0706_),
    .X(_1224_));
 sky130_fd_sc_hd__or4_4 _1971_ (.A(_1218_),
    .B(_1220_),
    .C(_1222_),
    .D(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__or2_2 _1972_ (.A(net91),
    .B(_0761_),
    .X(_1226_));
 sky130_fd_sc_hd__a21o_1 _1973_ (.A1(_1226_),
    .A2(_0979_),
    .B1(_0779_),
    .X(_1227_));
 sky130_fd_sc_hd__nand3_1 _1974_ (.A(net185),
    .B(_1225_),
    .C(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__a21o_1 _1975_ (.A1(_1225_),
    .A2(_1227_),
    .B1(net185),
    .X(_1229_));
 sky130_fd_sc_hd__inv_2 _1976_ (.A(net176),
    .Y(_1230_));
 sky130_fd_sc_hd__mux2_1 _1977_ (.A0(net116),
    .A1(net93),
    .S(_0691_),
    .X(_1231_));
 sky130_fd_sc_hd__a32o_1 _1978_ (.A1(_0890_),
    .A2(_1226_),
    .A3(_0971_),
    .B1(_1231_),
    .B2(_0773_),
    .X(_1232_));
 sky130_fd_sc_hd__mux2_1 _1979_ (.A0(net99),
    .A1(net115),
    .S(_0822_),
    .X(_1233_));
 sky130_fd_sc_hd__a32o_1 _1980_ (.A1(_0892_),
    .A2(_1005_),
    .A3(_0936_),
    .B1(_1233_),
    .B2(_0790_),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_1 _1981_ (.A0(net69),
    .A1(net78),
    .S(_0763_),
    .X(_1235_));
 sky130_fd_sc_hd__a32o_1 _1982_ (.A1(_0748_),
    .A2(_0858_),
    .A3(_0897_),
    .B1(_1235_),
    .B2(_0643_),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _1983_ (.A0(net74),
    .A1(net100),
    .S(_0761_),
    .X(_1237_));
 sky130_fd_sc_hd__o21a_1 _1984_ (.A1(_0707_),
    .A2(_1237_),
    .B1(_0706_),
    .X(_1238_));
 sky130_fd_sc_hd__or4_2 _1985_ (.A(_1232_),
    .B(_1234_),
    .C(_1236_),
    .D(_1238_),
    .X(_1239_));
 sky130_fd_sc_hd__a21o_1 _1986_ (.A1(_0956_),
    .A2(_0880_),
    .B1(_0779_),
    .X(_1240_));
 sky130_fd_sc_hd__and3_1 _1987_ (.A(_1230_),
    .B(_1239_),
    .C(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__a21oi_2 _1988_ (.A1(_1239_),
    .A2(_1240_),
    .B1(_1230_),
    .Y(_1242_));
 sky130_fd_sc_hd__a211o_2 _1989_ (.A1(_1228_),
    .A2(_1229_),
    .B1(_1241_),
    .C1(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__nand3_1 _1990_ (.A(_1230_),
    .B(_1239_),
    .C(_1240_),
    .Y(_1244_));
 sky130_fd_sc_hd__a21o_1 _1991_ (.A1(_1239_),
    .A2(_1240_),
    .B1(_1230_),
    .X(_1245_));
 sky130_fd_sc_hd__and3_1 _1992_ (.A(net185),
    .B(_1225_),
    .C(_1227_),
    .X(_1246_));
 sky130_fd_sc_hd__a21oi_2 _1993_ (.A1(_1225_),
    .A2(_1227_),
    .B1(net185),
    .Y(_1247_));
 sky130_fd_sc_hd__a211o_2 _1994_ (.A1(_1244_),
    .A2(_1245_),
    .B1(_1246_),
    .C1(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__and2_1 _1995_ (.A(_1243_),
    .B(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__and3_1 _1996_ (.A(_0716_),
    .B(_0953_),
    .C(_1005_),
    .X(_1250_));
 sky130_fd_sc_hd__and3_1 _1997_ (.A(_0668_),
    .B(_0935_),
    .C(_0897_),
    .X(_1251_));
 sky130_fd_sc_hd__a311o_1 _1998_ (.A1(_0981_),
    .A2(_0916_),
    .A3(_0909_),
    .B1(_1250_),
    .C1(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__and3_1 _1999_ (.A(_0657_),
    .B(_0857_),
    .C(_1021_),
    .X(_1253_));
 sky130_fd_sc_hd__and3_1 _2000_ (.A(_0696_),
    .B(_1226_),
    .C(_0913_),
    .X(_1254_));
 sky130_fd_sc_hd__or2_2 _2001_ (.A(_0885_),
    .B(_0860_),
    .X(_1255_));
 sky130_fd_sc_hd__and3_1 _2002_ (.A(_0643_),
    .B(_1255_),
    .C(_1026_),
    .X(_1256_));
 sky130_fd_sc_hd__and3_1 _2003_ (.A(_0674_),
    .B(_1039_),
    .C(_1019_),
    .X(_1257_));
 sky130_fd_sc_hd__or4_2 _2004_ (.A(_1253_),
    .B(_1254_),
    .C(_1256_),
    .D(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__and3_1 _2005_ (.A(_0788_),
    .B(_0872_),
    .C(_0930_),
    .X(_1259_));
 sky130_fd_sc_hd__nor3_4 _2006_ (.A(_1252_),
    .B(_1258_),
    .C(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__xor2_1 _2007_ (.A(net158),
    .B(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__buf_2 _2008_ (.A(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__o211a_1 _2009_ (.A1(net117),
    .A2(_0838_),
    .B1(_0839_),
    .C1(_0897_),
    .X(_1263_));
 sky130_fd_sc_hd__a31o_1 _2010_ (.A1(_0826_),
    .A2(_0952_),
    .A3(_0970_),
    .B1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__and3_1 _2011_ (.A(_0674_),
    .B(_0982_),
    .C(_1026_),
    .X(_1265_));
 sky130_fd_sc_hd__and3_1 _2012_ (.A(_0696_),
    .B(_0936_),
    .C(_0973_),
    .X(_1266_));
 sky130_fd_sc_hd__and3_1 _2013_ (.A(_0688_),
    .B(_0858_),
    .C(_0971_),
    .X(_1267_));
 sky130_fd_sc_hd__and3_1 _2014_ (.A(_0863_),
    .B(_0978_),
    .C(_1019_),
    .X(_1268_));
 sky130_fd_sc_hd__or4_1 _2015_ (.A(_1265_),
    .B(_1266_),
    .C(_1267_),
    .D(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__a311o_1 _2016_ (.A1(_0821_),
    .A2(_0979_),
    .A3(_1021_),
    .B1(_1264_),
    .C1(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__a31oi_4 _2017_ (.A1(_0819_),
    .A2(_0955_),
    .A3(_0888_),
    .B1(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__xnor2_4 _2018_ (.A(net181),
    .B(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__a21o_1 _2019_ (.A1(_1249_),
    .A2(_1262_),
    .B1(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__a21o_1 _2020_ (.A1(_1039_),
    .A2(_0970_),
    .B1(_0709_),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_1 _2021_ (.A0(net116),
    .A1(net106),
    .S(_0697_),
    .X(_1275_));
 sky130_fd_sc_hd__o21a_1 _2022_ (.A1(_0727_),
    .A2(_1275_),
    .B1(_0729_),
    .X(_1276_));
 sky130_fd_sc_hd__mux2_1 _2023_ (.A0(_0885_),
    .A1(net74),
    .S(_0697_),
    .X(_1277_));
 sky130_fd_sc_hd__a32o_1 _2024_ (.A1(_0790_),
    .A2(_0905_),
    .A3(_0880_),
    .B1(_1277_),
    .B2(_0721_),
    .X(_1278_));
 sky130_fd_sc_hd__mux2_1 _2025_ (.A0(net70),
    .A1(net118),
    .S(_0697_),
    .X(_1279_));
 sky130_fd_sc_hd__a32o_1 _2026_ (.A1(_0773_),
    .A2(_0879_),
    .A3(_0929_),
    .B1(_1279_),
    .B2(_0890_),
    .X(_1280_));
 sky130_fd_sc_hd__mux2_1 _2027_ (.A0(net75),
    .A1(net84),
    .S(_0651_),
    .X(_1281_));
 sky130_fd_sc_hd__a32o_1 _2028_ (.A1(_0681_),
    .A2(_0884_),
    .A3(_0888_),
    .B1(_1281_),
    .B2(_0643_),
    .X(_1282_));
 sky130_fd_sc_hd__or4_2 _2029_ (.A(_1276_),
    .B(_1278_),
    .C(_1280_),
    .D(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__nand3_1 _2030_ (.A(net167),
    .B(_1274_),
    .C(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__a21o_1 _2031_ (.A1(_1274_),
    .A2(_1283_),
    .B1(net167),
    .X(_1285_));
 sky130_fd_sc_hd__a211o_1 _2032_ (.A1(_1284_),
    .A2(_1285_),
    .B1(_1246_),
    .C1(_1247_),
    .X(_1286_));
 sky130_fd_sc_hd__and3_1 _2033_ (.A(net167),
    .B(_1274_),
    .C(_1283_),
    .X(_1287_));
 sky130_fd_sc_hd__a21oi_2 _2034_ (.A1(_1274_),
    .A2(_1283_),
    .B1(net167),
    .Y(_1288_));
 sky130_fd_sc_hd__a211o_2 _2035_ (.A1(_1228_),
    .A2(_1229_),
    .B1(_1287_),
    .C1(_1288_),
    .X(_1289_));
 sky130_fd_sc_hd__nand2_1 _2036_ (.A(_1286_),
    .B(_1289_),
    .Y(_1290_));
 sky130_fd_sc_hd__nor2_1 _2037_ (.A(_1262_),
    .B(_1290_),
    .Y(_1291_));
 sky130_fd_sc_hd__nor2_2 _2038_ (.A(_1287_),
    .B(_1288_),
    .Y(_1292_));
 sky130_fd_sc_hd__o211a_1 _2039_ (.A1(_1287_),
    .A2(_1288_),
    .B1(_1244_),
    .C1(_1245_),
    .X(_1293_));
 sky130_fd_sc_hd__a31o_1 _2040_ (.A1(_1292_),
    .A2(_1243_),
    .A3(_1248_),
    .B1(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__nand2_2 _2041_ (.A(_1284_),
    .B(_1285_),
    .Y(_1295_));
 sky130_fd_sc_hd__xnor2_4 _2042_ (.A(net158),
    .B(_1260_),
    .Y(_1296_));
 sky130_fd_sc_hd__nand2_1 _2043_ (.A(_1295_),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__xor2_4 _2044_ (.A(net181),
    .B(_1271_),
    .X(_1298_));
 sky130_fd_sc_hd__and3_1 _2045_ (.A(_1295_),
    .B(_1243_),
    .C(_1296_),
    .X(_1299_));
 sky130_fd_sc_hd__a311o_1 _2046_ (.A1(_1294_),
    .A2(_1286_),
    .A3(_1297_),
    .B1(_1298_),
    .C1(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__o21a_1 _2047_ (.A1(_1273_),
    .A2(_1291_),
    .B1(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__or4_1 _2048_ (.A(_1241_),
    .B(_1242_),
    .C(_1246_),
    .D(_1247_),
    .X(_1302_));
 sky130_fd_sc_hd__and3_1 _2049_ (.A(_1296_),
    .B(_1289_),
    .C(_1302_),
    .X(_1303_));
 sky130_fd_sc_hd__o21ai_1 _2050_ (.A1(_1273_),
    .A2(_1303_),
    .B1(_1300_),
    .Y(_1304_));
 sky130_fd_sc_hd__and3_1 _2051_ (.A(_0668_),
    .B(_1009_),
    .C(_0962_),
    .X(_1305_));
 sky130_fd_sc_hd__and3_1 _2052_ (.A(_0840_),
    .B(_0883_),
    .C(_0865_),
    .X(_1306_));
 sky130_fd_sc_hd__a311o_1 _2053_ (.A1(_0826_),
    .A2(_0864_),
    .A3(_0959_),
    .B1(_1305_),
    .C1(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__and3_1 _2054_ (.A(_0825_),
    .B(_0879_),
    .C(_0869_),
    .X(_1308_));
 sky130_fd_sc_hd__and3_1 _2055_ (.A(_0829_),
    .B(_0955_),
    .C(_0904_),
    .X(_0000_));
 sky130_fd_sc_hd__and3_1 _2056_ (.A(_0981_),
    .B(_0954_),
    .C(_0868_),
    .X(_0001_));
 sky130_fd_sc_hd__a31o_1 _2057_ (.A1(_0832_),
    .A2(_0872_),
    .A3(_0956_),
    .B1(_0001_),
    .X(_0002_));
 sky130_fd_sc_hd__or4_2 _2058_ (.A(_1307_),
    .B(_1308_),
    .C(_0000_),
    .D(_0002_),
    .X(_0003_));
 sky130_fd_sc_hd__a31oi_4 _2059_ (.A1(_0819_),
    .A2(_1255_),
    .A3(_0973_),
    .B1(_0003_),
    .Y(_0004_));
 sky130_fd_sc_hd__xnor2_4 _2060_ (.A(net150),
    .B(_0004_),
    .Y(_0005_));
 sky130_fd_sc_hd__mux2_2 _2061_ (.A0(_1301_),
    .A1(_1304_),
    .S(_0005_),
    .X(_0006_));
 sky130_fd_sc_hd__mux2_2 _2062_ (.A0(\L[28] ),
    .A1(net18),
    .S(_0855_),
    .X(_0007_));
 sky130_fd_sc_hd__xnor2_4 _2063_ (.A(_0006_),
    .B(_0007_),
    .Y(net142));
 sky130_fd_sc_hd__mux2_1 _2064_ (.A0(net81),
    .A1(net72),
    .S(_0670_),
    .X(_0008_));
 sky130_fd_sc_hd__a32o_1 _2065_ (.A1(_0648_),
    .A2(_0667_),
    .A3(_0746_),
    .B1(_0008_),
    .B2(_0687_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _2066_ (.A0(net71),
    .A1(net113),
    .S(_0661_),
    .X(_0010_));
 sky130_fd_sc_hd__a32o_1 _2067_ (.A1(_0683_),
    .A2(_0673_),
    .A3(_0738_),
    .B1(_0010_),
    .B2(_0656_),
    .X(_0011_));
 sky130_fd_sc_hd__mux2_1 _2068_ (.A0(net86),
    .A1(net97),
    .S(_0661_),
    .X(_0012_));
 sky130_fd_sc_hd__a32o_1 _2069_ (.A1(_0748_),
    .A2(_0676_),
    .A3(_0792_),
    .B1(_0012_),
    .B2(_0737_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _2070_ (.A0(net96),
    .A1(net77),
    .S(_0647_),
    .X(_0014_));
 sky130_fd_sc_hd__o21a_1 _2071_ (.A1(_0707_),
    .A2(_0014_),
    .B1(_0706_),
    .X(_0015_));
 sky130_fd_sc_hd__or4_2 _2072_ (.A(_0009_),
    .B(_0011_),
    .C(_0013_),
    .D(_0015_),
    .X(_0016_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(net119),
    .B(_0795_),
    .Y(_0017_));
 sky130_fd_sc_hd__o21ai_1 _2074_ (.A1(_1120_),
    .A2(_0017_),
    .B1(_0751_),
    .Y(_0018_));
 sky130_fd_sc_hd__and3b_1 _2075_ (.A_N(net178),
    .B(_0016_),
    .C(_0018_),
    .X(_0019_));
 sky130_fd_sc_hd__a21boi_2 _2076_ (.A1(_0016_),
    .A2(_0018_),
    .B1_N(net178),
    .Y(_0020_));
 sky130_fd_sc_hd__and3_1 _2077_ (.A(_0642_),
    .B(_0719_),
    .C(_0789_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _2078_ (.A0(net94),
    .A1(net72),
    .S(_0649_),
    .X(_0022_));
 sky130_fd_sc_hd__a32o_1 _2079_ (.A1(_0686_),
    .A2(_0714_),
    .A3(_0833_),
    .B1(_0022_),
    .B2(_0666_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _2080_ (.A0(net119),
    .A1(net103),
    .S(_0649_),
    .X(_0024_));
 sky130_fd_sc_hd__a32o_1 _2081_ (.A1(_0672_),
    .A2(_1118_),
    .A3(_0830_),
    .B1(_0024_),
    .B2(_0695_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _2082_ (.A0(net113),
    .A1(net88),
    .S(_0649_),
    .X(_0026_));
 sky130_fd_sc_hd__a32o_1 _2083_ (.A1(_0655_),
    .A2(_0704_),
    .A3(_0831_),
    .B1(_0026_),
    .B2(_0748_),
    .X(_0027_));
 sky130_fd_sc_hd__or4_1 _2084_ (.A(_0021_),
    .B(_0023_),
    .C(_0025_),
    .D(_0027_),
    .X(_0028_));
 sky130_fd_sc_hd__and3_1 _2085_ (.A(_0662_),
    .B(_0751_),
    .C(_0801_),
    .X(_0029_));
 sky130_fd_sc_hd__o21ai_1 _2086_ (.A1(_0028_),
    .A2(_0029_),
    .B1(net161),
    .Y(_0030_));
 sky130_fd_sc_hd__or3_1 _2087_ (.A(net161),
    .B(_0028_),
    .C(_0029_),
    .X(_0031_));
 sky130_fd_sc_hd__or4bb_1 _2088_ (.A(_0019_),
    .B(_0020_),
    .C_N(_0030_),
    .D_N(_0031_),
    .X(_0032_));
 sky130_fd_sc_hd__inv_2 _2089_ (.A(net169),
    .Y(_0033_));
 sky130_fd_sc_hd__mux2_1 _2090_ (.A0(net81),
    .A1(net90),
    .S(_0675_),
    .X(_0034_));
 sky130_fd_sc_hd__a32o_1 _2091_ (.A1(_0687_),
    .A2(_0766_),
    .A3(_0723_),
    .B1(_0034_),
    .B2(_0667_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2092_ (.A0(net104),
    .A1(net96),
    .S(_0670_),
    .X(_0036_));
 sky130_fd_sc_hd__a32o_1 _2093_ (.A1(_0656_),
    .A2(_0718_),
    .A3(_0835_),
    .B1(_0036_),
    .B2(_0673_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2094_ (.A0(net95),
    .A1(net71),
    .S(_0661_),
    .X(_0038_));
 sky130_fd_sc_hd__a32o_1 _2095_ (.A1(_0737_),
    .A2(_0752_),
    .A3(_0823_),
    .B1(_0038_),
    .B2(_0748_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(net111),
    .A1(net66),
    .S(_0675_),
    .X(_0040_));
 sky130_fd_sc_hd__o21a_1 _2097_ (.A1(_0707_),
    .A2(_0040_),
    .B1(_0706_),
    .X(_0041_));
 sky130_fd_sc_hd__or4_1 _2098_ (.A(_0035_),
    .B(_0037_),
    .C(_0039_),
    .D(_0041_),
    .X(_0042_));
 sky130_fd_sc_hd__a21o_1 _2099_ (.A1(_0677_),
    .A2(_0802_),
    .B1(_0708_),
    .X(_0043_));
 sky130_fd_sc_hd__and3_1 _2100_ (.A(_0033_),
    .B(_0042_),
    .C(_0043_),
    .X(_0044_));
 sky130_fd_sc_hd__a21oi_2 _2101_ (.A1(_0042_),
    .A2(_0043_),
    .B1(_0033_),
    .Y(_0045_));
 sky130_fd_sc_hd__o22a_1 _2102_ (.A1(_0019_),
    .A2(_0020_),
    .B1(_0044_),
    .B2(_0045_),
    .X(_0046_));
 sky130_fd_sc_hd__and3b_1 _2103_ (.A_N(_1120_),
    .B(_0824_),
    .C(_0797_),
    .X(_0047_));
 sky130_fd_sc_hd__a31o_1 _2104_ (.A1(_0821_),
    .A2(_0762_),
    .A3(_0789_),
    .B1(_0047_),
    .X(_0048_));
 sky130_fd_sc_hd__and3_1 _2105_ (.A(_0644_),
    .B(_0766_),
    .C(_0754_),
    .X(_0049_));
 sky130_fd_sc_hd__a31o_1 _2106_ (.A1(_0840_),
    .A2(_1122_),
    .A3(_0833_),
    .B1(_0049_),
    .X(_0050_));
 sky130_fd_sc_hd__and3_1 _2107_ (.A(_0799_),
    .B(_0703_),
    .C(_0835_),
    .X(_0051_));
 sky130_fd_sc_hd__a31o_1 _2108_ (.A1(_0834_),
    .A2(_0823_),
    .A3(_0831_),
    .B1(_0751_),
    .X(_0052_));
 sky130_fd_sc_hd__a311o_1 _2109_ (.A1(_0682_),
    .A2(_0771_),
    .A3(_0830_),
    .B1(_0051_),
    .C1(_0052_),
    .X(_0053_));
 sky130_fd_sc_hd__a21o_1 _2110_ (.A1(_0698_),
    .A2(_0738_),
    .B1(_0709_),
    .X(_0054_));
 sky130_fd_sc_hd__o31a_1 _2111_ (.A1(_0048_),
    .A2(_0050_),
    .A3(_0053_),
    .B1(_0054_),
    .X(_0055_));
 sky130_fd_sc_hd__xor2_2 _2112_ (.A(net152),
    .B(_0055_),
    .X(_0056_));
 sky130_fd_sc_hd__and2b_1 _2113_ (.A_N(_0046_),
    .B(_0056_),
    .X(_0057_));
 sky130_fd_sc_hd__nand2_1 _2114_ (.A(_0032_),
    .B(_0057_),
    .Y(_0058_));
 sky130_fd_sc_hd__and2_1 _2115_ (.A(_0030_),
    .B(_0031_),
    .X(_0059_));
 sky130_fd_sc_hd__clkbuf_2 _2116_ (.A(_0059_),
    .X(_0060_));
 sky130_fd_sc_hd__or4_2 _2117_ (.A(_0019_),
    .B(_0020_),
    .C(_0044_),
    .D(_0045_),
    .X(_0061_));
 sky130_fd_sc_hd__and2b_1 _2118_ (.A_N(_0046_),
    .B(_0061_),
    .X(_0062_));
 sky130_fd_sc_hd__nor2_2 _2119_ (.A(_0044_),
    .B(_0045_),
    .Y(_0063_));
 sky130_fd_sc_hd__buf_2 _2120_ (.A(_0056_),
    .X(_0064_));
 sky130_fd_sc_hd__a21oi_1 _2121_ (.A1(_0060_),
    .A2(_0063_),
    .B1(_0064_),
    .Y(_0065_));
 sky130_fd_sc_hd__o21ai_1 _2122_ (.A1(_0060_),
    .A2(_0062_),
    .B1(_0065_),
    .Y(_0066_));
 sky130_fd_sc_hd__o211a_1 _2123_ (.A1(net95),
    .A2(_0796_),
    .B1(_0981_),
    .C1(_0767_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2124_ (.A0(net66),
    .A1(net109),
    .S(_0753_),
    .X(_0068_));
 sky130_fd_sc_hd__a32o_1 _2125_ (.A1(_0829_),
    .A2(_0752_),
    .A3(_0713_),
    .B1(_0068_),
    .B2(_0832_),
    .X(_0069_));
 sky130_fd_sc_hd__a311o_1 _2126_ (.A1(_0826_),
    .A2(_0718_),
    .A3(_0723_),
    .B1(_0067_),
    .C1(_0069_),
    .X(_0070_));
 sky130_fd_sc_hd__o211a_1 _2127_ (.A1(net94),
    .A2(_0796_),
    .B1(_0839_),
    .C1(_0762_),
    .X(_0071_));
 sky130_fd_sc_hd__a31o_1 _2128_ (.A1(_0668_),
    .A2(_0704_),
    .A3(_1122_),
    .B1(_0788_),
    .X(_0072_));
 sky130_fd_sc_hd__a311o_1 _2129_ (.A1(_0825_),
    .A2(_0766_),
    .A3(_0719_),
    .B1(_0071_),
    .C1(_0072_),
    .X(_0073_));
 sky130_fd_sc_hd__a21o_1 _2130_ (.A1(_0669_),
    .A2(_0740_),
    .B1(_0709_),
    .X(_0074_));
 sky130_fd_sc_hd__o21ai_4 _2131_ (.A1(_0070_),
    .A2(_0073_),
    .B1(_0074_),
    .Y(_0075_));
 sky130_fd_sc_hd__xnor2_4 _2132_ (.A(net187),
    .B(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__a21oi_1 _2133_ (.A1(_0058_),
    .A2(_0066_),
    .B1(_0076_),
    .Y(_0077_));
 sky130_fd_sc_hd__and3_1 _2134_ (.A(_0682_),
    .B(_0831_),
    .C(_0833_),
    .X(_0078_));
 sky130_fd_sc_hd__a31o_1 _2135_ (.A1(_0840_),
    .A2(_0771_),
    .A3(_1123_),
    .B1(_0078_),
    .X(_0079_));
 sky130_fd_sc_hd__o211a_1 _2136_ (.A1(net103),
    .A2(_0838_),
    .B1(_0703_),
    .C1(_0644_),
    .X(_0080_));
 sky130_fd_sc_hd__a31o_1 _2137_ (.A1(_0829_),
    .A2(_0754_),
    .A3(_0789_),
    .B1(_0080_),
    .X(_0081_));
 sky130_fd_sc_hd__and3_1 _2138_ (.A(_0668_),
    .B(_0724_),
    .C(_0835_),
    .X(_0082_));
 sky130_fd_sc_hd__a311o_1 _2139_ (.A1(_0825_),
    .A2(_0823_),
    .A3(_0714_),
    .B1(_0081_),
    .C1(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__a311o_1 _2140_ (.A1(_0981_),
    .A2(_0824_),
    .A3(_0830_),
    .B1(_0079_),
    .C1(_0083_),
    .X(_0084_));
 sky130_fd_sc_hd__a31oi_4 _2141_ (.A1(_0648_),
    .A2(_0819_),
    .A3(_0741_),
    .B1(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__xnor2_4 _2142_ (.A(net143),
    .B(_0085_),
    .Y(_0086_));
 sky130_fd_sc_hd__a31o_1 _2143_ (.A1(_0076_),
    .A2(_0058_),
    .A3(_0066_),
    .B1(_0086_),
    .X(_0087_));
 sky130_fd_sc_hd__and3b_1 _2144_ (.A_N(_0046_),
    .B(_0061_),
    .C(_0060_),
    .X(_0088_));
 sky130_fd_sc_hd__nand2_1 _2145_ (.A(_0030_),
    .B(_0031_),
    .Y(_0089_));
 sky130_fd_sc_hd__and2_1 _2146_ (.A(_0089_),
    .B(_0063_),
    .X(_0090_));
 sky130_fd_sc_hd__o21ai_1 _2147_ (.A1(_0088_),
    .A2(_0090_),
    .B1(_0064_),
    .Y(_0091_));
 sky130_fd_sc_hd__or3_1 _2148_ (.A(_0064_),
    .B(_0088_),
    .C(_0090_),
    .X(_0092_));
 sky130_fd_sc_hd__and3_1 _2149_ (.A(_0076_),
    .B(_0091_),
    .C(_0092_),
    .X(_0093_));
 sky130_fd_sc_hd__or2_2 _2150_ (.A(_0019_),
    .B(_0020_),
    .X(_0094_));
 sky130_fd_sc_hd__nor2_1 _2151_ (.A(_0094_),
    .B(_0089_),
    .Y(_0095_));
 sky130_fd_sc_hd__a2bb2o_1 _2152_ (.A1_N(_0019_),
    .A2_N(_0020_),
    .B1(_0030_),
    .B2(_0031_),
    .X(_0096_));
 sky130_fd_sc_hd__nand2_1 _2153_ (.A(_0064_),
    .B(_0096_),
    .Y(_0097_));
 sky130_fd_sc_hd__o21bai_2 _2154_ (.A1(_0094_),
    .A2(_0060_),
    .B1_N(_0056_),
    .Y(_0098_));
 sky130_fd_sc_hd__o22a_1 _2155_ (.A1(_0095_),
    .A2(_0097_),
    .B1(_0098_),
    .B2(_0088_),
    .X(_0099_));
 sky130_fd_sc_hd__o21ai_1 _2156_ (.A1(_0076_),
    .A2(_0099_),
    .B1(_0086_),
    .Y(_0100_));
 sky130_fd_sc_hd__o22a_1 _2157_ (.A1(_0077_),
    .A2(_0087_),
    .B1(_0093_),
    .B2(_0100_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2158_ (.A0(\L[27] ),
    .A1(net9),
    .S(_0855_),
    .X(_0102_));
 sky130_fd_sc_hd__xnor2_2 _2159_ (.A(_0101_),
    .B(_0102_),
    .Y(net133));
 sky130_fd_sc_hd__o211a_1 _2160_ (.A1(net117),
    .A2(_0838_),
    .B1(_0829_),
    .C1(_0982_),
    .X(_0103_));
 sky130_fd_sc_hd__a31o_1 _2161_ (.A1(_0826_),
    .A2(_0896_),
    .A3(_0979_),
    .B1(_0103_),
    .X(_0104_));
 sky130_fd_sc_hd__and3_1 _2162_ (.A(_0644_),
    .B(_0912_),
    .C(_0971_),
    .X(_0105_));
 sky130_fd_sc_hd__a31o_1 _2163_ (.A1(_0840_),
    .A2(_1039_),
    .A3(_0936_),
    .B1(_0105_),
    .X(_0106_));
 sky130_fd_sc_hd__o211a_1 _2164_ (.A1(net67),
    .A2(_0796_),
    .B1(_0981_),
    .C1(_0978_),
    .X(_0107_));
 sky130_fd_sc_hd__a311o_1 _2165_ (.A1(_0825_),
    .A2(_0857_),
    .A3(_0973_),
    .B1(_0106_),
    .C1(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__a311o_1 _2166_ (.A1(_0821_),
    .A2(_0952_),
    .A3(_0976_),
    .B1(_0104_),
    .C1(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__a31oi_4 _2167_ (.A1(_0819_),
    .A2(_0879_),
    .A3(_1012_),
    .B1(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__xnor2_4 _2168_ (.A(_0627_),
    .B(_0110_),
    .Y(_0111_));
 sky130_fd_sc_hd__and3_1 _2169_ (.A(_0721_),
    .B(_0909_),
    .C(_1019_),
    .X(_0112_));
 sky130_fd_sc_hd__and3_1 _2170_ (.A(_0839_),
    .B(_1255_),
    .C(_0858_),
    .X(_0113_));
 sky130_fd_sc_hd__a311o_1 _2171_ (.A1(_0682_),
    .A2(_0913_),
    .A3(_1026_),
    .B1(_0112_),
    .C1(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__and3_1 _2172_ (.A(_0797_),
    .B(_0935_),
    .C(_0970_),
    .X(_0115_));
 sky130_fd_sc_hd__and3_1 _2173_ (.A(_0799_),
    .B(_1005_),
    .C(_0916_),
    .X(_0116_));
 sky130_fd_sc_hd__and3_1 _2174_ (.A(_0863_),
    .B(_0953_),
    .C(_1021_),
    .X(_0117_));
 sky130_fd_sc_hd__a31o_1 _2175_ (.A1(_0981_),
    .A2(_1226_),
    .A3(_0897_),
    .B1(_0117_),
    .X(_0118_));
 sky130_fd_sc_hd__or4_1 _2176_ (.A(_0114_),
    .B(_0115_),
    .C(_0116_),
    .D(_0118_),
    .X(_0119_));
 sky130_fd_sc_hd__a31o_1 _2177_ (.A1(_0819_),
    .A2(_0883_),
    .A3(_0873_),
    .B1(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__xor2_2 _2178_ (.A(net159),
    .B(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__buf_2 _2179_ (.A(_0121_),
    .X(_0122_));
 sky130_fd_sc_hd__and3_1 _2180_ (.A(_0716_),
    .B(_0868_),
    .C(_0883_),
    .X(_0123_));
 sky130_fd_sc_hd__o211a_1 _2181_ (.A1(net75),
    .A2(_0795_),
    .B1(_0668_),
    .C1(_0904_),
    .X(_0124_));
 sky130_fd_sc_hd__a311o_1 _2182_ (.A1(_0825_),
    .A2(_0954_),
    .A3(_0884_),
    .B1(_0123_),
    .C1(_0124_),
    .X(_0125_));
 sky130_fd_sc_hd__and3_1 _2183_ (.A(_0799_),
    .B(_0872_),
    .C(_0962_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _2184_ (.A0(net76),
    .A1(_0885_),
    .S(_0702_),
    .X(_0127_));
 sky130_fd_sc_hd__a32o_1 _2185_ (.A1(_0834_),
    .A2(_0879_),
    .A3(_0864_),
    .B1(_0127_),
    .B2(_0644_),
    .X(_0128_));
 sky130_fd_sc_hd__a311o_1 _2186_ (.A1(_0840_),
    .A2(_0959_),
    .A3(_0880_),
    .B1(_0126_),
    .C1(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__and3_1 _2187_ (.A(_0788_),
    .B(_0913_),
    .C(_0978_),
    .X(_0130_));
 sky130_fd_sc_hd__nor3_4 _2188_ (.A(_0125_),
    .B(_0129_),
    .C(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__xor2_2 _2189_ (.A(net156),
    .B(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__and3_1 _2190_ (.A(_0643_),
    .B(_0904_),
    .C(_0873_),
    .X(_0133_));
 sky130_fd_sc_hd__and3_1 _2191_ (.A(_0696_),
    .B(_0956_),
    .C(_1009_),
    .X(_0134_));
 sky130_fd_sc_hd__a311o_1 _2192_ (.A1(_0834_),
    .A2(_0959_),
    .A3(_0869_),
    .B1(_0133_),
    .C1(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__and3_1 _2193_ (.A(_0773_),
    .B(_0864_),
    .C(_0930_),
    .X(_0136_));
 sky130_fd_sc_hd__and3_1 _2194_ (.A(_0892_),
    .B(_0955_),
    .C(_1012_),
    .X(_0137_));
 sky130_fd_sc_hd__and3_1 _2195_ (.A(_0681_),
    .B(_0954_),
    .C(_0865_),
    .X(_0138_));
 sky130_fd_sc_hd__and3_1 _2196_ (.A(_0890_),
    .B(_0868_),
    .C(_0929_),
    .X(_0139_));
 sky130_fd_sc_hd__or4_2 _2197_ (.A(_0136_),
    .B(_0137_),
    .C(_0138_),
    .D(_0139_),
    .X(_0140_));
 sky130_fd_sc_hd__and3_1 _2198_ (.A(_0751_),
    .B(_0976_),
    .C(_1021_),
    .X(_0141_));
 sky130_fd_sc_hd__nor3_4 _2199_ (.A(_0135_),
    .B(_0140_),
    .C(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__xor2_2 _2200_ (.A(net165),
    .B(_0142_),
    .X(_0143_));
 sky130_fd_sc_hd__a21o_1 _2201_ (.A1(_1009_),
    .A2(_0884_),
    .B1(_0779_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _2202_ (.A0(net92),
    .A1(net82),
    .S(_0647_),
    .X(_0145_));
 sky130_fd_sc_hd__o21a_1 _2203_ (.A1(_0707_),
    .A2(_0145_),
    .B1(_0706_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2204_ (.A0(net101),
    .A1(net108),
    .S(_0675_),
    .X(_0147_));
 sky130_fd_sc_hd__a32o_1 _2205_ (.A1(_0656_),
    .A2(_0909_),
    .A3(_0979_),
    .B1(_0147_),
    .B2(_0673_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2206_ (.A0(_0885_),
    .A1(net117),
    .S(_0675_),
    .X(_0149_));
 sky130_fd_sc_hd__a32o_1 _2207_ (.A1(_0687_),
    .A2(_0896_),
    .A3(_0857_),
    .B1(_0149_),
    .B2(_0667_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(net107),
    .A1(net67),
    .S(_0647_),
    .X(_0151_));
 sky130_fd_sc_hd__a32o_1 _2209_ (.A1(_0737_),
    .A2(_0935_),
    .A3(_0982_),
    .B1(_0151_),
    .B2(_0748_),
    .X(_0152_));
 sky130_fd_sc_hd__or4_4 _2210_ (.A(_0146_),
    .B(_0148_),
    .C(_0150_),
    .D(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__and3_1 _2211_ (.A(_0623_),
    .B(_0144_),
    .C(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__a21oi_2 _2212_ (.A1(_0144_),
    .A2(_0153_),
    .B1(_0623_),
    .Y(_0155_));
 sky130_fd_sc_hd__a21o_1 _2213_ (.A1(_0912_),
    .A2(_1019_),
    .B1(_0708_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2214_ (.A0(net101),
    .A1(net91),
    .S(_0658_),
    .X(_0157_));
 sky130_fd_sc_hd__o21a_1 _2215_ (.A1(_0707_),
    .A2(_0157_),
    .B1(_0706_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2216_ (.A0(net82),
    .A1(net74),
    .S(_0658_),
    .X(_0159_));
 sky130_fd_sc_hd__a32o_1 _2217_ (.A1(_0656_),
    .A2(_0962_),
    .A3(_0924_),
    .B1(_0159_),
    .B2(_0673_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2218_ (.A0(net85),
    .A1(net106),
    .S(_0646_),
    .X(_0161_));
 sky130_fd_sc_hd__a32o_1 _2219_ (.A1(_0667_),
    .A2(_0883_),
    .A3(_0905_),
    .B1(_0161_),
    .B2(_0687_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2220_ (.A0(net116),
    .A1(net75),
    .S(_0658_),
    .X(_0163_));
 sky130_fd_sc_hd__a32o_1 _2221_ (.A1(_0737_),
    .A2(_0879_),
    .A3(_0888_),
    .B1(_0163_),
    .B2(_0748_),
    .X(_0164_));
 sky130_fd_sc_hd__or4_1 _2222_ (.A(_0158_),
    .B(_0160_),
    .C(_0162_),
    .D(_0164_),
    .X(_0165_));
 sky130_fd_sc_hd__and3_1 _2223_ (.A(net183),
    .B(_0156_),
    .C(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__a21oi_1 _2224_ (.A1(_0156_),
    .A2(_0165_),
    .B1(net183),
    .Y(_0167_));
 sky130_fd_sc_hd__o22a_1 _2225_ (.A1(_0154_),
    .A2(_0155_),
    .B1(_0166_),
    .B2(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__xnor2_1 _2226_ (.A(_0143_),
    .B(_0168_),
    .Y(_0169_));
 sky130_fd_sc_hd__nor2_1 _2227_ (.A(_0132_),
    .B(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__nor2_2 _2228_ (.A(_0154_),
    .B(_0155_),
    .Y(_0171_));
 sky130_fd_sc_hd__or2_1 _2229_ (.A(_0166_),
    .B(_0167_),
    .X(_0172_));
 sky130_fd_sc_hd__buf_2 _2230_ (.A(_0172_),
    .X(_0173_));
 sky130_fd_sc_hd__xor2_1 _2231_ (.A(_0171_),
    .B(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__o21ai_1 _2232_ (.A1(_0171_),
    .A2(_0143_),
    .B1(_0132_),
    .Y(_0175_));
 sky130_fd_sc_hd__a21oi_1 _2233_ (.A1(_0143_),
    .A2(_0174_),
    .B1(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__or3_1 _2234_ (.A(_0122_),
    .B(_0170_),
    .C(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__nand3_1 _2235_ (.A(_0623_),
    .B(_0144_),
    .C(_0153_),
    .Y(_0178_));
 sky130_fd_sc_hd__a21o_1 _2236_ (.A1(_0144_),
    .A2(_0153_),
    .B1(_0623_),
    .X(_0179_));
 sky130_fd_sc_hd__a211o_1 _2237_ (.A1(_0178_),
    .A2(_0179_),
    .B1(_0166_),
    .C1(_0167_),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_1 _2238_ (.A(_0143_),
    .B(_0180_),
    .Y(_0181_));
 sky130_fd_sc_hd__a21oi_1 _2239_ (.A1(_0171_),
    .A2(_0173_),
    .B1(_0132_),
    .Y(_0182_));
 sky130_fd_sc_hd__xnor2_4 _2240_ (.A(net165),
    .B(_0142_),
    .Y(_0183_));
 sky130_fd_sc_hd__xnor2_4 _2241_ (.A(net156),
    .B(_0131_),
    .Y(_0184_));
 sky130_fd_sc_hd__a21oi_1 _2242_ (.A1(_0173_),
    .A2(_0183_),
    .B1(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__a22o_1 _2243_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_0185_),
    .B2(_0180_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_1 _2244_ (.A(_0122_),
    .B(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__or4_2 _2245_ (.A(_0154_),
    .B(_0155_),
    .C(_0166_),
    .D(_0167_),
    .X(_0188_));
 sky130_fd_sc_hd__xnor2_1 _2246_ (.A(_0188_),
    .B(_0183_),
    .Y(_0189_));
 sky130_fd_sc_hd__xnor2_1 _2247_ (.A(_0171_),
    .B(_0173_),
    .Y(_0190_));
 sky130_fd_sc_hd__mux2_1 _2248_ (.A0(_0189_),
    .A1(_0190_),
    .S(_0184_),
    .X(_0191_));
 sky130_fd_sc_hd__a21oi_1 _2249_ (.A1(_0122_),
    .A2(_0191_),
    .B1(_0111_),
    .Y(_0192_));
 sky130_fd_sc_hd__nor2_1 _2250_ (.A(_0188_),
    .B(_0183_),
    .Y(_0193_));
 sky130_fd_sc_hd__nor2_1 _2251_ (.A(_0173_),
    .B(_0183_),
    .Y(_0194_));
 sky130_fd_sc_hd__a21o_1 _2252_ (.A1(_0183_),
    .A2(_0168_),
    .B1(_0184_),
    .X(_0195_));
 sky130_fd_sc_hd__o32a_1 _2253_ (.A1(_0193_),
    .A2(_0132_),
    .A3(_0169_),
    .B1(_0194_),
    .B2(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _2254_ (.A(_0122_),
    .B(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__a32o_1 _2255_ (.A1(_0111_),
    .A2(_0177_),
    .A3(_0187_),
    .B1(_0192_),
    .B2(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2256_ (.A0(\L[26] ),
    .A1(net64),
    .S(_0855_),
    .X(_0199_));
 sky130_fd_sc_hd__xnor2_2 _2257_ (.A(_0198_),
    .B(_0199_),
    .Y(net188));
 sky130_fd_sc_hd__mux2_1 _2258_ (.A0(net94),
    .A1(net103),
    .S(_0702_),
    .X(_0200_));
 sky130_fd_sc_hd__a32o_1 _2259_ (.A1(_0799_),
    .A2(_0714_),
    .A3(_1123_),
    .B1(_0200_),
    .B2(_0834_),
    .X(_0201_));
 sky130_fd_sc_hd__a31o_1 _2260_ (.A1(_0832_),
    .A2(_0704_),
    .A3(_0824_),
    .B1(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2261_ (.A0(net109),
    .A1(net87),
    .S(_0702_),
    .X(_0203_));
 sky130_fd_sc_hd__a32o_1 _2262_ (.A1(_0839_),
    .A2(_0767_),
    .A3(_0789_),
    .B1(_0203_),
    .B2(_0668_),
    .X(_0204_));
 sky130_fd_sc_hd__and3_1 _2263_ (.A(_0716_),
    .B(_0719_),
    .C(_0724_),
    .X(_0205_));
 sky130_fd_sc_hd__a311o_1 _2264_ (.A1(_0797_),
    .A2(_0718_),
    .A3(_0754_),
    .B1(_0204_),
    .C1(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__and3_1 _2265_ (.A(_0652_),
    .B(_0788_),
    .C(_0792_),
    .X(_0207_));
 sky130_fd_sc_hd__nor3_4 _2266_ (.A(_0202_),
    .B(_0206_),
    .C(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__xnor2_1 _2267_ (.A(net159),
    .B(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__buf_2 _2268_ (.A(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2269_ (.A0(net72),
    .A1(net112),
    .S(_0691_),
    .X(_0211_));
 sky130_fd_sc_hd__a32o_1 _2270_ (.A1(_0790_),
    .A2(_0746_),
    .A3(_0801_),
    .B1(_0211_),
    .B2(_0696_),
    .X(_0212_));
 sky130_fd_sc_hd__and3_1 _2271_ (.A(_0648_),
    .B(_0890_),
    .C(_0820_),
    .X(_0213_));
 sky130_fd_sc_hd__a311o_1 _2272_ (.A1(_0660_),
    .A2(_0668_),
    .A3(_0738_),
    .B1(_0212_),
    .C1(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__and3_1 _2273_ (.A(_0737_),
    .B(_0676_),
    .C(_0732_),
    .X(_0215_));
 sky130_fd_sc_hd__and3_1 _2274_ (.A(_0656_),
    .B(_0669_),
    .C(_1116_),
    .X(_0216_));
 sky130_fd_sc_hd__o211a_1 _2275_ (.A1(net97),
    .A2(_0753_),
    .B1(_0748_),
    .C1(_0802_),
    .X(_0217_));
 sky130_fd_sc_hd__or4_1 _2276_ (.A(_0751_),
    .B(_0215_),
    .C(_0216_),
    .D(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__a21o_1 _2277_ (.A1(_0762_),
    .A2(_0714_),
    .B1(_0779_),
    .X(_0219_));
 sky130_fd_sc_hd__o21ai_1 _2278_ (.A1(_0214_),
    .A2(_0218_),
    .B1(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__xnor2_1 _2279_ (.A(net128),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__buf_2 _2280_ (.A(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2281_ (.A0(net79),
    .A1(net103),
    .S(_0670_),
    .X(_0223_));
 sky130_fd_sc_hd__a32o_1 _2282_ (.A1(_0737_),
    .A2(_0778_),
    .A3(_0746_),
    .B1(_0223_),
    .B2(_0748_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _2283_ (.A0(net89),
    .A1(net97),
    .S(_0675_),
    .X(_0225_));
 sky130_fd_sc_hd__a32o_1 _2284_ (.A1(_0687_),
    .A2(_0732_),
    .A3(_0741_),
    .B1(_0225_),
    .B2(_0667_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _2285_ (.A0(net109),
    .A1(net72),
    .S(_0670_),
    .X(_0227_));
 sky130_fd_sc_hd__a32o_1 _2286_ (.A1(_0662_),
    .A2(_0673_),
    .A3(_0792_),
    .B1(_0227_),
    .B2(_0656_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _2287_ (.A0(net119),
    .A1(net88),
    .S(_0647_),
    .X(_0229_));
 sky130_fd_sc_hd__o21a_1 _2288_ (.A1(_0707_),
    .A2(_0229_),
    .B1(_0706_),
    .X(_0230_));
 sky130_fd_sc_hd__or4_1 _2289_ (.A(_0224_),
    .B(_0226_),
    .C(_0228_),
    .D(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__a21o_1 _2290_ (.A1(_0718_),
    .A2(_0830_),
    .B1(_0708_),
    .X(_0232_));
 sky130_fd_sc_hd__and3b_1 _2291_ (.A_N(net136),
    .B(_0231_),
    .C(_0232_),
    .X(_0233_));
 sky130_fd_sc_hd__a21boi_2 _2292_ (.A1(_0231_),
    .A2(_0232_),
    .B1_N(net136),
    .Y(_0234_));
 sky130_fd_sc_hd__mux2_1 _2293_ (.A0(net90),
    .A1(net95),
    .S(_0763_),
    .X(_0235_));
 sky130_fd_sc_hd__a32o_1 _2294_ (.A1(_0737_),
    .A2(_0662_),
    .A3(_0683_),
    .B1(_0235_),
    .B2(_0748_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2295_ (.A0(net66),
    .A1(net120),
    .S(_0763_),
    .X(_0237_));
 sky130_fd_sc_hd__a32o_1 _2296_ (.A1(_0667_),
    .A2(_0677_),
    .A3(_0692_),
    .B1(_0237_),
    .B2(_0687_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _2297_ (.A0(net94),
    .A1(net86),
    .S(_0647_),
    .X(_0239_));
 sky130_fd_sc_hd__a32o_1 _2298_ (.A1(_0648_),
    .A2(_0656_),
    .A3(_1178_),
    .B1(_0239_),
    .B2(_0673_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2299_ (.A0(net105),
    .A1(net80),
    .S(_0763_),
    .X(_0241_));
 sky130_fd_sc_hd__o21a_1 _2300_ (.A1(_0707_),
    .A2(_0241_),
    .B1(_0706_),
    .X(_0242_));
 sky130_fd_sc_hd__or4_1 _2301_ (.A(_0236_),
    .B(_0238_),
    .C(_0240_),
    .D(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__a21o_1 _2302_ (.A1(_0771_),
    .A2(_0719_),
    .B1(_0779_),
    .X(_0244_));
 sky130_fd_sc_hd__and3b_1 _2303_ (.A_N(net145),
    .B(_0243_),
    .C(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__a21boi_1 _2304_ (.A1(_0243_),
    .A2(_0244_),
    .B1_N(net145),
    .Y(_0246_));
 sky130_fd_sc_hd__o22a_2 _2305_ (.A1(_0233_),
    .A2(_0234_),
    .B1(_0245_),
    .B2(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__or4_4 _2306_ (.A(_0233_),
    .B(_0234_),
    .C(_0245_),
    .D(_0246_),
    .X(_0248_));
 sky130_fd_sc_hd__and2b_1 _2307_ (.A_N(_0247_),
    .B(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__xor2_1 _2308_ (.A(_0222_),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_4 _2309_ (.A(_0221_),
    .X(_0251_));
 sky130_fd_sc_hd__and3b_1 _2310_ (.A_N(_0247_),
    .B(_0248_),
    .C(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_1 _2311_ (.A(_0233_),
    .B(_0234_),
    .Y(_0253_));
 sky130_fd_sc_hd__nor2_1 _2312_ (.A(_0222_),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__xor2_4 _2313_ (.A(net159),
    .B(_0208_),
    .X(_0255_));
 sky130_fd_sc_hd__and3_1 _2314_ (.A(_0648_),
    .B(_0981_),
    .C(_0802_),
    .X(_0256_));
 sky130_fd_sc_hd__o211a_1 _2315_ (.A1(net97),
    .A2(_0838_),
    .B1(_0840_),
    .C1(_0699_),
    .X(_0257_));
 sky130_fd_sc_hd__a311o_1 _2316_ (.A1(_0826_),
    .A2(_0669_),
    .A3(_0801_),
    .B1(_0256_),
    .C1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__and3_1 _2317_ (.A(_0660_),
    .B(_0829_),
    .C(_0676_),
    .X(_0259_));
 sky130_fd_sc_hd__o211a_1 _2318_ (.A1(net72),
    .A2(_0796_),
    .B1(_0683_),
    .C1(_0668_),
    .X(_0260_));
 sky130_fd_sc_hd__a31o_1 _2319_ (.A1(_0832_),
    .A2(_0692_),
    .A3(_0792_),
    .B1(_0260_),
    .X(_0261_));
 sky130_fd_sc_hd__a311o_1 _2320_ (.A1(_0698_),
    .A2(_0825_),
    .A3(_0746_),
    .B1(_0259_),
    .C1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__and3_1 _2321_ (.A(_0788_),
    .B(_0723_),
    .C(_0824_),
    .X(_0263_));
 sky130_fd_sc_hd__nor3_4 _2322_ (.A(_0258_),
    .B(_0262_),
    .C(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__xnor2_2 _2323_ (.A(net154),
    .B(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__o31a_1 _2324_ (.A1(_0252_),
    .A2(_0254_),
    .A3(_0255_),
    .B1(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__o21ai_1 _2325_ (.A1(_0210_),
    .A2(_0250_),
    .B1(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__and3_1 _2326_ (.A(_0682_),
    .B(_0677_),
    .C(_0741_),
    .X(_0268_));
 sky130_fd_sc_hd__a31o_1 _2327_ (.A1(_0829_),
    .A2(_0778_),
    .A3(_1178_),
    .B1(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__a31o_1 _2328_ (.A1(_0662_),
    .A2(_0981_),
    .A3(_0740_),
    .B1(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__and3_1 _2329_ (.A(_0644_),
    .B(_0671_),
    .C(_0820_),
    .X(_0271_));
 sky130_fd_sc_hd__a31o_1 _2330_ (.A1(_0840_),
    .A2(_0690_),
    .A3(_0738_),
    .B1(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__and3_1 _2331_ (.A(_0685_),
    .B(_0825_),
    .C(_0732_),
    .X(_0273_));
 sky130_fd_sc_hd__a311o_1 _2332_ (.A1(_0652_),
    .A2(_0821_),
    .A3(_1116_),
    .B1(_0272_),
    .C1(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__o211a_1 _2333_ (.A1(net95),
    .A2(_0796_),
    .B1(_0788_),
    .C1(_0833_),
    .X(_0275_));
 sky130_fd_sc_hd__or3_2 _2334_ (.A(_0270_),
    .B(_0274_),
    .C(_0275_),
    .X(_0276_));
 sky130_fd_sc_hd__xor2_4 _2335_ (.A(net183),
    .B(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__nor2_1 _2336_ (.A(_0245_),
    .B(_0246_),
    .Y(_0278_));
 sky130_fd_sc_hd__buf_2 _2337_ (.A(_0278_),
    .X(_0279_));
 sky130_fd_sc_hd__xor2_1 _2338_ (.A(_0251_),
    .B(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__or2_1 _2339_ (.A(_0233_),
    .B(_0234_),
    .X(_0281_));
 sky130_fd_sc_hd__clkbuf_2 _2340_ (.A(_0281_),
    .X(_0282_));
 sky130_fd_sc_hd__a21o_1 _2341_ (.A1(_0282_),
    .A2(_0279_),
    .B1(_0255_),
    .X(_0283_));
 sky130_fd_sc_hd__nor2_1 _2342_ (.A(_0251_),
    .B(_0279_),
    .Y(_0284_));
 sky130_fd_sc_hd__xor2_4 _2343_ (.A(net154),
    .B(_0264_),
    .X(_0285_));
 sky130_fd_sc_hd__o221ai_2 _2344_ (.A1(_0210_),
    .A2(_0280_),
    .B1(_0283_),
    .B2(_0284_),
    .C1(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__or2_1 _2345_ (.A(_0251_),
    .B(_0253_),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_1 _2346_ (.A(_0282_),
    .B(_0279_),
    .Y(_0288_));
 sky130_fd_sc_hd__and3b_1 _2347_ (.A_N(_0222_),
    .B(_0248_),
    .C(_0255_),
    .X(_0289_));
 sky130_fd_sc_hd__a311o_1 _2348_ (.A1(_0287_),
    .A2(_0210_),
    .A3(_0288_),
    .B1(_0289_),
    .C1(_0265_),
    .X(_0290_));
 sky130_fd_sc_hd__a21o_1 _2349_ (.A1(_0222_),
    .A2(_0279_),
    .B1(_0247_),
    .X(_0291_));
 sky130_fd_sc_hd__a21oi_1 _2350_ (.A1(_0251_),
    .A2(_0279_),
    .B1(_0282_),
    .Y(_0292_));
 sky130_fd_sc_hd__a221o_1 _2351_ (.A1(_0283_),
    .A2(_0291_),
    .B1(_0292_),
    .B2(_0210_),
    .C1(_0285_),
    .X(_0293_));
 sky130_fd_sc_hd__a21oi_1 _2352_ (.A1(_0290_),
    .A2(_0293_),
    .B1(_0277_),
    .Y(_0294_));
 sky130_fd_sc_hd__a31oi_2 _2353_ (.A1(_0267_),
    .A2(_0277_),
    .A3(_0286_),
    .B1(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__mux2_1 _2354_ (.A0(net196),
    .A1(net2),
    .S(_0855_),
    .X(_0296_));
 sky130_fd_sc_hd__xnor2_1 _2355_ (.A(_0295_),
    .B(_0296_),
    .Y(net126));
 sky130_fd_sc_hd__a31o_1 _2356_ (.A1(_1085_),
    .A2(_1107_),
    .A3(_1061_),
    .B1(_1031_),
    .X(_0297_));
 sky130_fd_sc_hd__and3_1 _2357_ (.A(_1073_),
    .B(_1091_),
    .C(_1085_),
    .X(_0298_));
 sky130_fd_sc_hd__a31o_1 _2358_ (.A1(_1060_),
    .A2(_1086_),
    .A3(_1092_),
    .B1(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__a21bo_1 _2359_ (.A1(_1085_),
    .A2(_1062_),
    .B1_N(_1101_),
    .X(_0300_));
 sky130_fd_sc_hd__o22a_1 _2360_ (.A1(_1111_),
    .A2(_0297_),
    .B1(_0299_),
    .B2(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__o211a_1 _2361_ (.A1(_1095_),
    .A2(_1074_),
    .B1(_1098_),
    .C1(_1110_),
    .X(_0302_));
 sky130_fd_sc_hd__a21oi_1 _2362_ (.A1(_1109_),
    .A2(_1110_),
    .B1(_1098_),
    .Y(_0303_));
 sky130_fd_sc_hd__o32ai_1 _2363_ (.A1(_1101_),
    .A2(_1111_),
    .A3(_0302_),
    .B1(_0303_),
    .B2(_0300_),
    .Y(_0304_));
 sky130_fd_sc_hd__mux2_2 _2364_ (.A0(_0301_),
    .A1(_0304_),
    .S(_1017_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_2 _2365_ (.A0(\L[24] ),
    .A1(net55),
    .S(_0855_),
    .X(_0306_));
 sky130_fd_sc_hd__xnor2_4 _2366_ (.A(_0305_),
    .B(_0306_),
    .Y(net179));
 sky130_fd_sc_hd__a311oi_1 _2367_ (.A1(_0944_),
    .A2(_0949_),
    .A3(_0990_),
    .B1(_1000_),
    .C1(_0940_),
    .Y(_0307_));
 sky130_fd_sc_hd__and3_1 _2368_ (.A(_0901_),
    .B(_0940_),
    .C(_0949_),
    .X(_0308_));
 sky130_fd_sc_hd__o21ai_1 _2369_ (.A1(_0307_),
    .A2(_0308_),
    .B1(_0988_),
    .Y(_0309_));
 sky130_fd_sc_hd__and2_1 _2370_ (.A(_0877_),
    .B(_0878_),
    .X(_0310_));
 sky130_fd_sc_hd__o31ai_4 _2371_ (.A1(_0920_),
    .A2(_0921_),
    .A3(_0943_),
    .B1(_0939_),
    .Y(_0311_));
 sky130_fd_sc_hd__a21o_1 _2372_ (.A1(_0310_),
    .A2(_0996_),
    .B1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__a21o_1 _2373_ (.A1(_0946_),
    .A2(_0312_),
    .B1(_0988_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _2374_ (.A(_0944_),
    .B(_0949_),
    .Y(_0314_));
 sky130_fd_sc_hd__or2_1 _2375_ (.A(_0943_),
    .B(_0949_),
    .X(_0315_));
 sky130_fd_sc_hd__and3_1 _2376_ (.A(_0947_),
    .B(_0314_),
    .C(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__nand2_1 _2377_ (.A(_0949_),
    .B(_0990_),
    .Y(_0317_));
 sky130_fd_sc_hd__a211oi_1 _2378_ (.A1(_0944_),
    .A2(_0317_),
    .B1(_1000_),
    .C1(_0947_),
    .Y(_0318_));
 sky130_fd_sc_hd__o21ai_1 _2379_ (.A1(_0316_),
    .A2(_0318_),
    .B1(_0989_),
    .Y(_0319_));
 sky130_fd_sc_hd__o221a_1 _2380_ (.A1(_0940_),
    .A2(_0950_),
    .B1(_0317_),
    .B2(_0311_),
    .C1(_0988_),
    .X(_0320_));
 sky130_fd_sc_hd__nor2_1 _2381_ (.A(_0968_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__a32o_2 _2382_ (.A1(_0968_),
    .A2(_0309_),
    .A3(_0313_),
    .B1(_0319_),
    .B2(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_2 _2383_ (.A0(\L[23] ),
    .A1(net47),
    .S(_1114_),
    .X(_0323_));
 sky130_fd_sc_hd__xor2_4 _2384_ (.A(_0322_),
    .B(_0323_),
    .X(net171));
 sky130_fd_sc_hd__o21a_1 _2385_ (.A1(_0810_),
    .A2(_0849_),
    .B1(_0759_),
    .X(_0324_));
 sky130_fd_sc_hd__and3b_1 _2386_ (.A_N(_0810_),
    .B(_0736_),
    .C(_0785_),
    .X(_0325_));
 sky130_fd_sc_hd__o21ai_1 _2387_ (.A1(_0324_),
    .A2(_0325_),
    .B1(_0712_),
    .Y(_0326_));
 sky130_fd_sc_hd__o21ai_1 _2388_ (.A1(_0850_),
    .A2(_0760_),
    .B1(_0812_),
    .Y(_0327_));
 sky130_fd_sc_hd__a21oi_1 _2389_ (.A1(_0326_),
    .A2(_0327_),
    .B1(_0808_),
    .Y(_0328_));
 sky130_fd_sc_hd__o211ai_1 _2390_ (.A1(_0810_),
    .A2(_0785_),
    .B1(_0783_),
    .C1(_0812_),
    .Y(_0329_));
 sky130_fd_sc_hd__a31o_1 _2391_ (.A1(_0808_),
    .A2(_0326_),
    .A3(_0329_),
    .B1(_0845_),
    .X(_0330_));
 sky130_fd_sc_hd__a21oi_1 _2392_ (.A1(_0783_),
    .A2(_0784_),
    .B1(_0812_),
    .Y(_0331_));
 sky130_fd_sc_hd__and3_1 _2393_ (.A(_0812_),
    .B(_0810_),
    .C(_0849_),
    .X(_0332_));
 sky130_fd_sc_hd__or3_1 _2394_ (.A(_0759_),
    .B(_0331_),
    .C(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__o21ai_1 _2395_ (.A1(_0331_),
    .A2(_0332_),
    .B1(_0759_),
    .Y(_0334_));
 sky130_fd_sc_hd__o21a_1 _2396_ (.A1(_0810_),
    .A2(_0785_),
    .B1(_0736_),
    .X(_0335_));
 sky130_fd_sc_hd__a211o_1 _2397_ (.A1(_0810_),
    .A2(_0759_),
    .B1(_0849_),
    .C1(_0712_),
    .X(_0336_));
 sky130_fd_sc_hd__o211a_1 _2398_ (.A1(_0812_),
    .A2(_0335_),
    .B1(_0336_),
    .C1(_0807_),
    .X(_0337_));
 sky130_fd_sc_hd__a31o_1 _2399_ (.A1(_0808_),
    .A2(_0333_),
    .A3(_0334_),
    .B1(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__a2bb2o_2 _2400_ (.A1_N(_0328_),
    .A2_N(_0330_),
    .B1(_0338_),
    .B2(_0845_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_2 _2401_ (.A0(\L[22] ),
    .A1(net38),
    .S(_0855_),
    .X(_0340_));
 sky130_fd_sc_hd__xnor2_4 _2402_ (.A(_0339_),
    .B(_0340_),
    .Y(net162));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(\L[21] ),
    .A1(net29),
    .S(_1114_),
    .X(_0341_));
 sky130_fd_sc_hd__o211a_1 _2404_ (.A1(_0032_),
    .A2(_0063_),
    .B1(_0056_),
    .C1(_0096_),
    .X(_0342_));
 sky130_fd_sc_hd__o21ba_1 _2405_ (.A1(_0062_),
    .A2(_0098_),
    .B1_N(_0342_),
    .X(_0343_));
 sky130_fd_sc_hd__a21o_1 _2406_ (.A1(_0094_),
    .A2(_0065_),
    .B1(_0342_),
    .X(_0344_));
 sky130_fd_sc_hd__xnor2_1 _2407_ (.A(_0089_),
    .B(_0061_),
    .Y(_0345_));
 sky130_fd_sc_hd__xnor2_1 _2408_ (.A(_0057_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__a22o_1 _2409_ (.A1(_0063_),
    .A2(_0056_),
    .B1(_0061_),
    .B2(_0096_),
    .X(_0347_));
 sky130_fd_sc_hd__a21bo_1 _2410_ (.A1(_0060_),
    .A2(_0057_),
    .B1_N(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__xor2_2 _2411_ (.A(net187),
    .B(_0075_),
    .X(_0349_));
 sky130_fd_sc_hd__mux4_2 _2412_ (.A0(_0343_),
    .A1(_0344_),
    .A2(_0346_),
    .A3(_0348_),
    .S0(_0086_),
    .S1(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__xor2_2 _2413_ (.A(_0341_),
    .B(_0350_),
    .X(net153));
 sky130_fd_sc_hd__inv_2 _2414_ (.A(_0121_),
    .Y(_0351_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(_0196_),
    .A1(_0191_),
    .S(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__o21a_1 _2416_ (.A1(_0170_),
    .A2(_0176_),
    .B1(_0122_),
    .X(_0353_));
 sky130_fd_sc_hd__a21bo_1 _2417_ (.A1(_0351_),
    .A2(_0186_),
    .B1_N(_0111_),
    .X(_0354_));
 sky130_fd_sc_hd__o22a_1 _2418_ (.A1(_0111_),
    .A2(_0352_),
    .B1(_0353_),
    .B2(_0354_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(\L[20] ),
    .A1(net20),
    .S(_1114_),
    .X(_0356_));
 sky130_fd_sc_hd__xor2_2 _2420_ (.A(_0355_),
    .B(_0356_),
    .X(net144));
 sky130_fd_sc_hd__and2_1 _2421_ (.A(_1202_),
    .B(_1205_),
    .X(_0357_));
 sky130_fd_sc_hd__and3_1 _2422_ (.A(_1153_),
    .B(_1154_),
    .C(_1195_),
    .X(_0358_));
 sky130_fd_sc_hd__or3_1 _2423_ (.A(_1194_),
    .B(_0357_),
    .C(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__nand2_2 _2424_ (.A(_1203_),
    .B(_1195_),
    .Y(_0360_));
 sky130_fd_sc_hd__o21ai_1 _2425_ (.A1(_1203_),
    .A2(_1195_),
    .B1(_1193_),
    .Y(_0361_));
 sky130_fd_sc_hd__a21o_1 _2426_ (.A1(_1205_),
    .A2(_0360_),
    .B1(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__a21oi_1 _2427_ (.A1(_0359_),
    .A2(_0362_),
    .B1(_1182_),
    .Y(_0363_));
 sky130_fd_sc_hd__o21ai_1 _2428_ (.A1(_0357_),
    .A2(_0358_),
    .B1(_1194_),
    .Y(_0364_));
 sky130_fd_sc_hd__a31o_1 _2429_ (.A1(_1182_),
    .A2(_0359_),
    .A3(_0364_),
    .B1(_1130_),
    .X(_0365_));
 sky130_fd_sc_hd__nand2_1 _2430_ (.A(_1195_),
    .B(_1182_),
    .Y(_0366_));
 sky130_fd_sc_hd__mux2_1 _2431_ (.A0(_1205_),
    .A1(_1182_),
    .S(_1195_),
    .X(_0367_));
 sky130_fd_sc_hd__a221oi_1 _2432_ (.A1(_1211_),
    .A2(_0366_),
    .B1(_0367_),
    .B2(_1141_),
    .C1(_1194_),
    .Y(_0368_));
 sky130_fd_sc_hd__and3_1 _2433_ (.A(_1167_),
    .B(_1168_),
    .C(_1194_),
    .X(_0369_));
 sky130_fd_sc_hd__or3_1 _2434_ (.A(_1203_),
    .B(_1205_),
    .C(_1182_),
    .X(_0370_));
 sky130_fd_sc_hd__a21bo_1 _2435_ (.A1(_0369_),
    .A2(_0370_),
    .B1_N(_1130_),
    .X(_0371_));
 sky130_fd_sc_hd__o22a_1 _2436_ (.A1(_0363_),
    .A2(_0365_),
    .B1(_0368_),
    .B2(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _2437_ (.A0(net192),
    .A1(net11),
    .S(_0855_),
    .X(_0373_));
 sky130_fd_sc_hd__xnor2_1 _2438_ (.A(_0372_),
    .B(_0373_),
    .Y(net135));
 sky130_fd_sc_hd__nor2_2 _2439_ (.A(_1241_),
    .B(_1242_),
    .Y(_0374_));
 sky130_fd_sc_hd__nor2_1 _2440_ (.A(_1246_),
    .B(_1247_),
    .Y(_0375_));
 sky130_fd_sc_hd__o21a_1 _2441_ (.A1(_0374_),
    .A2(_0375_),
    .B1(_1296_),
    .X(_0376_));
 sky130_fd_sc_hd__nand2_1 _2442_ (.A(_1292_),
    .B(_0375_),
    .Y(_0377_));
 sky130_fd_sc_hd__and3_1 _2443_ (.A(_1243_),
    .B(_1286_),
    .C(_1262_),
    .X(_0378_));
 sky130_fd_sc_hd__a21oi_1 _2444_ (.A1(_0376_),
    .A2(_0377_),
    .B1(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__o21ba_1 _2445_ (.A1(_1298_),
    .A2(_0379_),
    .B1_N(_0005_),
    .X(_0380_));
 sky130_fd_sc_hd__nand2_1 _2446_ (.A(_1295_),
    .B(_0374_),
    .Y(_0381_));
 sky130_fd_sc_hd__a21o_1 _2447_ (.A1(_1286_),
    .A2(_1289_),
    .B1(_0374_),
    .X(_0382_));
 sky130_fd_sc_hd__a21oi_1 _2448_ (.A1(_0381_),
    .A2(_0382_),
    .B1(_1262_),
    .Y(_0383_));
 sky130_fd_sc_hd__a211o_1 _2449_ (.A1(_1294_),
    .A2(_1262_),
    .B1(_1272_),
    .C1(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_1 _2450_ (.A(_1244_),
    .B(_1245_),
    .Y(_0385_));
 sky130_fd_sc_hd__a22o_1 _2451_ (.A1(_0385_),
    .A2(_1262_),
    .B1(_0376_),
    .B2(_1286_),
    .X(_0386_));
 sky130_fd_sc_hd__o21ai_1 _2452_ (.A1(_1272_),
    .A2(_0386_),
    .B1(_0005_),
    .Y(_0387_));
 sky130_fd_sc_hd__nor2_1 _2453_ (.A(_1295_),
    .B(_0374_),
    .Y(_0388_));
 sky130_fd_sc_hd__a211o_1 _2454_ (.A1(_1295_),
    .A2(_1249_),
    .B1(_1296_),
    .C1(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__and3b_1 _2455_ (.A_N(_1291_),
    .B(_0389_),
    .C(_1272_),
    .X(_0390_));
 sky130_fd_sc_hd__o2bb2a_1 _2456_ (.A1_N(_0380_),
    .A2_N(_0384_),
    .B1(_0387_),
    .B2(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__buf_4 _2457_ (.A(_0605_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _2458_ (.A0(\L[18] ),
    .A1(net3),
    .S(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__xnor2_2 _2459_ (.A(_0391_),
    .B(_0393_),
    .Y(net127));
 sky130_fd_sc_hd__nand2_1 _2460_ (.A(_0992_),
    .B(_0996_),
    .Y(_0394_));
 sky130_fd_sc_hd__a211o_1 _2461_ (.A1(_0944_),
    .A2(_0317_),
    .B1(_1000_),
    .C1(_0940_),
    .X(_0395_));
 sky130_fd_sc_hd__o211a_1 _2462_ (.A1(_0947_),
    .A2(_0394_),
    .B1(_0395_),
    .C1(_0967_),
    .X(_0396_));
 sky130_fd_sc_hd__and2b_1 _2463_ (.A_N(_0311_),
    .B(_0902_),
    .X(_0397_));
 sky130_fd_sc_hd__o21a_1 _2464_ (.A1(_0316_),
    .A2(_0397_),
    .B1(_0968_),
    .X(_0398_));
 sky130_fd_sc_hd__a21o_1 _2465_ (.A1(_0945_),
    .A2(_0992_),
    .B1(_0940_),
    .X(_0399_));
 sky130_fd_sc_hd__nand3_1 _2466_ (.A(_0902_),
    .B(_0940_),
    .C(_0990_),
    .Y(_0400_));
 sky130_fd_sc_hd__a21oi_1 _2467_ (.A1(_0399_),
    .A2(_0400_),
    .B1(_0967_),
    .Y(_0401_));
 sky130_fd_sc_hd__nor2_1 _2468_ (.A(_0947_),
    .B(_0950_),
    .Y(_0402_));
 sky130_fd_sc_hd__and3b_1 _2469_ (.A_N(_0948_),
    .B(_0317_),
    .C(_0947_),
    .X(_0403_));
 sky130_fd_sc_hd__o31ai_1 _2470_ (.A1(_0968_),
    .A2(_0402_),
    .A3(_0403_),
    .B1(_0989_),
    .Y(_0404_));
 sky130_fd_sc_hd__o32a_2 _2471_ (.A1(_0989_),
    .A2(_0396_),
    .A3(_0398_),
    .B1(_0401_),
    .B2(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_2 _2472_ (.A0(\L[17] ),
    .A1(net24),
    .S(_0392_),
    .X(_0406_));
 sky130_fd_sc_hd__xnor2_4 _2473_ (.A(_0405_),
    .B(_0406_),
    .Y(net148));
 sky130_fd_sc_hd__a21bo_1 _2474_ (.A1(_1095_),
    .A2(_1091_),
    .B1_N(_1060_),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _2475_ (.A(_1074_),
    .B(_1086_),
    .Y(_0408_));
 sky130_fd_sc_hd__a221o_1 _2476_ (.A1(_1103_),
    .A2(_0407_),
    .B1(_0408_),
    .B2(_1096_),
    .C1(_1032_),
    .X(_0409_));
 sky130_fd_sc_hd__nor2_1 _2477_ (.A(_1098_),
    .B(_0407_),
    .Y(_0410_));
 sky130_fd_sc_hd__a21o_1 _2478_ (.A1(_1085_),
    .A2(_0407_),
    .B1(_1101_),
    .X(_0411_));
 sky130_fd_sc_hd__o21a_1 _2479_ (.A1(_0410_),
    .A2(_0411_),
    .B1(_1017_),
    .X(_0412_));
 sky130_fd_sc_hd__a21o_1 _2480_ (.A1(_1109_),
    .A2(_1075_),
    .B1(_1086_),
    .X(_0413_));
 sky130_fd_sc_hd__and2_1 _2481_ (.A(_1073_),
    .B(_1091_),
    .X(_0414_));
 sky130_fd_sc_hd__nor2_1 _2482_ (.A(_1073_),
    .B(_1074_),
    .Y(_0415_));
 sky130_fd_sc_hd__o31a_1 _2483_ (.A1(_1085_),
    .A2(_0414_),
    .A3(_0415_),
    .B1(_1101_),
    .X(_0416_));
 sky130_fd_sc_hd__and3_1 _2484_ (.A(_1060_),
    .B(_1086_),
    .C(_1075_),
    .X(_0417_));
 sky130_fd_sc_hd__o2bb2a_1 _2485_ (.A1_N(_0413_),
    .A2_N(_0416_),
    .B1(_0411_),
    .B2(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__o2bb2a_1 _2486_ (.A1_N(_0409_),
    .A2_N(_0412_),
    .B1(_0418_),
    .B2(_1017_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _2487_ (.A0(\L[16] ),
    .A1(net58),
    .S(_0392_),
    .X(_0420_));
 sky130_fd_sc_hd__xnor2_2 _2488_ (.A(_0419_),
    .B(_0420_),
    .Y(net182));
 sky130_fd_sc_hd__nor2_1 _2489_ (.A(_0089_),
    .B(_0063_),
    .Y(_0421_));
 sky130_fd_sc_hd__o21bai_1 _2490_ (.A1(_0060_),
    .A2(_0062_),
    .B1_N(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__o31ai_1 _2491_ (.A1(_0064_),
    .A2(_0090_),
    .A3(_0421_),
    .B1(_0349_),
    .Y(_0423_));
 sky130_fd_sc_hd__a21oi_1 _2492_ (.A1(_0064_),
    .A2(_0422_),
    .B1(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__and3_1 _2493_ (.A(_0094_),
    .B(_0060_),
    .C(_0063_),
    .X(_0425_));
 sky130_fd_sc_hd__a21oi_1 _2494_ (.A1(_0094_),
    .A2(_0063_),
    .B1(_0060_),
    .Y(_0426_));
 sky130_fd_sc_hd__nand2_1 _2495_ (.A(_0064_),
    .B(_0061_),
    .Y(_0427_));
 sky130_fd_sc_hd__o32a_1 _2496_ (.A1(_0064_),
    .A2(_0425_),
    .A3(_0426_),
    .B1(_0427_),
    .B2(_0421_),
    .X(_0428_));
 sky130_fd_sc_hd__a21bo_1 _2497_ (.A1(_0076_),
    .A2(_0428_),
    .B1_N(_0086_),
    .X(_0429_));
 sky130_fd_sc_hd__and3_1 _2498_ (.A(_0349_),
    .B(_0094_),
    .C(_0063_),
    .X(_0430_));
 sky130_fd_sc_hd__a211o_1 _2499_ (.A1(_0076_),
    .A2(_0090_),
    .B1(_0430_),
    .C1(_0095_),
    .X(_0431_));
 sky130_fd_sc_hd__a211o_1 _2500_ (.A1(_0094_),
    .A2(_0063_),
    .B1(_0064_),
    .C1(_0095_),
    .X(_0432_));
 sky130_fd_sc_hd__a21boi_1 _2501_ (.A1(_0064_),
    .A2(_0431_),
    .B1_N(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__o22a_2 _2502_ (.A1(_0424_),
    .A2(_0429_),
    .B1(_0433_),
    .B2(_0086_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_2 _2503_ (.A0(\L[15] ),
    .A1(net49),
    .S(_1114_),
    .X(_0435_));
 sky130_fd_sc_hd__xor2_4 _2504_ (.A(_0434_),
    .B(_0435_),
    .X(net173));
 sky130_fd_sc_hd__xnor2_1 _2505_ (.A(_0251_),
    .B(_0247_),
    .Y(_0436_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(_0279_),
    .A1(_0247_),
    .S(_0251_),
    .X(_0437_));
 sky130_fd_sc_hd__nor2_1 _2507_ (.A(_0255_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__a31o_1 _2508_ (.A1(_0248_),
    .A2(_0255_),
    .A3(_0436_),
    .B1(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__nand2_1 _2509_ (.A(_0222_),
    .B(_0279_),
    .Y(_0440_));
 sky130_fd_sc_hd__o21a_1 _2510_ (.A1(_0251_),
    .A2(_0282_),
    .B1(_0255_),
    .X(_0441_));
 sky130_fd_sc_hd__o21bai_1 _2511_ (.A1(_0222_),
    .A2(_0282_),
    .B1_N(_0252_),
    .Y(_0442_));
 sky130_fd_sc_hd__a22oi_1 _2512_ (.A1(_0440_),
    .A2(_0441_),
    .B1(_0442_),
    .B2(_0210_),
    .Y(_0443_));
 sky130_fd_sc_hd__xnor2_1 _2513_ (.A(_0251_),
    .B(_0278_),
    .Y(_0444_));
 sky130_fd_sc_hd__nor2_1 _2514_ (.A(_0253_),
    .B(_0210_),
    .Y(_0445_));
 sky130_fd_sc_hd__xnor2_1 _2515_ (.A(_0444_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__nor2_1 _2516_ (.A(_0254_),
    .B(_0255_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor2_1 _2517_ (.A(_0222_),
    .B(_0248_),
    .Y(_0448_));
 sky130_fd_sc_hd__nor2_1 _2518_ (.A(_0252_),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__a22o_1 _2519_ (.A1(_0249_),
    .A2(_0447_),
    .B1(_0449_),
    .B2(_0255_),
    .X(_0450_));
 sky130_fd_sc_hd__mux4_1 _2520_ (.A0(_0439_),
    .A1(_0443_),
    .A2(_0446_),
    .A3(_0450_),
    .S0(_0277_),
    .S1(_0285_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _2521_ (.A0(\L[14] ),
    .A1(net40),
    .S(_0392_),
    .X(_0452_));
 sky130_fd_sc_hd__xnor2_1 _2522_ (.A(_0451_),
    .B(_0452_),
    .Y(net164));
 sky130_fd_sc_hd__a22o_1 _2523_ (.A1(_1293_),
    .A2(_0375_),
    .B1(_1302_),
    .B2(_1292_),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _2524_ (.A(_0376_),
    .B(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__a21o_1 _2525_ (.A1(_0376_),
    .A2(_0453_),
    .B1(_1298_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(_1249_),
    .A1(_0453_),
    .S(_1262_),
    .X(_0456_));
 sky130_fd_sc_hd__o22a_1 _2527_ (.A1(_0454_),
    .A2(_0455_),
    .B1(_0456_),
    .B2(_1272_),
    .X(_0457_));
 sky130_fd_sc_hd__and3_1 _2528_ (.A(_1249_),
    .B(_1296_),
    .C(_1289_),
    .X(_0458_));
 sky130_fd_sc_hd__nor2_1 _2529_ (.A(_0374_),
    .B(_1261_),
    .Y(_0459_));
 sky130_fd_sc_hd__a21oi_1 _2530_ (.A1(_1248_),
    .A2(_1289_),
    .B1(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__and2_1 _2531_ (.A(_1290_),
    .B(_0459_),
    .X(_0461_));
 sky130_fd_sc_hd__o21ai_1 _2532_ (.A1(_1290_),
    .A2(_0459_),
    .B1(_1298_),
    .Y(_0462_));
 sky130_fd_sc_hd__o32a_1 _2533_ (.A1(_1298_),
    .A2(_0458_),
    .A3(_0460_),
    .B1(_0461_),
    .B2(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_2 _2534_ (.A0(_0457_),
    .A1(_0463_),
    .S(_0005_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_2 _2535_ (.A0(\L[13] ),
    .A1(net31),
    .S(_0392_),
    .X(_0465_));
 sky130_fd_sc_hd__xnor2_4 _2536_ (.A(_0464_),
    .B(_0465_),
    .Y(net155));
 sky130_fd_sc_hd__a21bo_1 _2537_ (.A1(_0810_),
    .A2(_0785_),
    .B1_N(_0786_),
    .X(_0466_));
 sky130_fd_sc_hd__mux4_1 _2538_ (.A0(_0848_),
    .A1(_0852_),
    .A2(_0466_),
    .A3(_0851_),
    .S0(_0808_),
    .S1(_0712_),
    .X(_0467_));
 sky130_fd_sc_hd__xnor2_1 _2539_ (.A(_0809_),
    .B(_0785_),
    .Y(_0468_));
 sky130_fd_sc_hd__a211oi_1 _2540_ (.A1(_0712_),
    .A2(_0468_),
    .B1(_0325_),
    .C1(_0332_),
    .Y(_0469_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(_0816_),
    .A1(_0468_),
    .S(_0712_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _2542_ (.A0(_0469_),
    .A1(_0470_),
    .S(_0808_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _2543_ (.A0(_0467_),
    .A1(_0471_),
    .S(_0845_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_2 _2544_ (.A0(\L[12] ),
    .A1(net22),
    .S(_0392_),
    .X(_0473_));
 sky130_fd_sc_hd__xnor2_2 _2545_ (.A(_0472_),
    .B(_0473_),
    .Y(net146));
 sky130_fd_sc_hd__and3_1 _2546_ (.A(_1169_),
    .B(_1194_),
    .C(_1200_),
    .X(_0474_));
 sky130_fd_sc_hd__o21ai_1 _2547_ (.A1(_1203_),
    .A2(_1205_),
    .B1(_1167_),
    .Y(_0475_));
 sky130_fd_sc_hd__nor2_1 _2548_ (.A(_1194_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__o21ai_1 _2549_ (.A1(_0474_),
    .A2(_0476_),
    .B1(_1182_),
    .Y(_0477_));
 sky130_fd_sc_hd__o211a_1 _2550_ (.A1(_1203_),
    .A2(_1204_),
    .B1(_1196_),
    .C1(_0360_),
    .X(_0478_));
 sky130_fd_sc_hd__a21oi_1 _2551_ (.A1(_1195_),
    .A2(_1209_),
    .B1(_0361_),
    .Y(_0479_));
 sky130_fd_sc_hd__or3_1 _2552_ (.A(_1182_),
    .B(_0478_),
    .C(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__o21ai_1 _2553_ (.A1(_1203_),
    .A2(_1195_),
    .B1(_1169_),
    .Y(_0481_));
 sky130_fd_sc_hd__a211o_1 _2554_ (.A1(_1194_),
    .A2(_0481_),
    .B1(_1201_),
    .C1(_1182_),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _2555_ (.A(_1168_),
    .B(_1196_),
    .Y(_0483_));
 sky130_fd_sc_hd__or2_1 _2556_ (.A(_0475_),
    .B(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__a21oi_1 _2557_ (.A1(_0475_),
    .A2(_0483_),
    .B1(_1212_),
    .Y(_0485_));
 sky130_fd_sc_hd__a21oi_1 _2558_ (.A1(_0484_),
    .A2(_0485_),
    .B1(_1130_),
    .Y(_0486_));
 sky130_fd_sc_hd__a32o_2 _2559_ (.A1(_1130_),
    .A2(_0477_),
    .A3(_0480_),
    .B1(_0482_),
    .B2(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_2 _2560_ (.A0(\L[11] ),
    .A1(net14),
    .S(_0392_),
    .X(_0488_));
 sky130_fd_sc_hd__xnor2_2 _2561_ (.A(_0487_),
    .B(_0488_),
    .Y(net138));
 sky130_fd_sc_hd__inv_2 _2562_ (.A(_0111_),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2_1 _2563_ (.A(_0183_),
    .B(_0168_),
    .Y(_0490_));
 sky130_fd_sc_hd__or2_1 _2564_ (.A(_0188_),
    .B(_0183_),
    .X(_0491_));
 sky130_fd_sc_hd__a32o_1 _2565_ (.A1(_0184_),
    .A2(_0490_),
    .A3(_0189_),
    .B1(_0185_),
    .B2(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _2566_ (.A0(_0169_),
    .A1(_0174_),
    .S(_0184_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(_0492_),
    .A1(_0493_),
    .S(_0121_),
    .X(_0494_));
 sky130_fd_sc_hd__a21bo_1 _2568_ (.A1(_0173_),
    .A2(_0183_),
    .B1_N(_0171_),
    .X(_0495_));
 sky130_fd_sc_hd__a21oi_1 _2569_ (.A1(_0183_),
    .A2(_0168_),
    .B1(_0184_),
    .Y(_0496_));
 sky130_fd_sc_hd__a22o_1 _2570_ (.A1(_0184_),
    .A2(_0189_),
    .B1(_0495_),
    .B2(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__nor2_1 _2571_ (.A(_0122_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(_0143_),
    .A1(_0171_),
    .S(_0173_),
    .X(_0499_));
 sky130_fd_sc_hd__a22o_1 _2573_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_0499_),
    .B2(_0132_),
    .X(_0500_));
 sky130_fd_sc_hd__a21o_1 _2574_ (.A1(_0122_),
    .A2(_0500_),
    .B1(_0111_),
    .X(_0501_));
 sky130_fd_sc_hd__o22a_1 _2575_ (.A1(_0489_),
    .A2(_0494_),
    .B1(_0498_),
    .B2(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(net191),
    .A1(net5),
    .S(_1114_),
    .X(_0503_));
 sky130_fd_sc_hd__xor2_1 _2577_ (.A(_0502_),
    .B(_0503_),
    .X(net129));
 sky130_fd_sc_hd__a21o_1 _2578_ (.A1(_0902_),
    .A2(_0992_),
    .B1(_0940_),
    .X(_0504_));
 sky130_fd_sc_hd__a21o_1 _2579_ (.A1(_0945_),
    .A2(_0992_),
    .B1(_0947_),
    .X(_0505_));
 sky130_fd_sc_hd__a21oi_1 _2580_ (.A1(_0902_),
    .A2(_0991_),
    .B1(_0967_),
    .Y(_0506_));
 sky130_fd_sc_hd__a32o_1 _2581_ (.A1(_0967_),
    .A2(_0400_),
    .A3(_0504_),
    .B1(_0505_),
    .B2(_0506_),
    .X(_0507_));
 sky130_fd_sc_hd__a32o_1 _2582_ (.A1(_0901_),
    .A2(_0940_),
    .A3(_0993_),
    .B1(_0991_),
    .B2(_0315_),
    .X(_0508_));
 sky130_fd_sc_hd__o21bai_1 _2583_ (.A1(_0922_),
    .A2(_0944_),
    .B1_N(_0310_),
    .Y(_0509_));
 sky130_fd_sc_hd__xor2_1 _2584_ (.A(_0311_),
    .B(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _2585_ (.A0(_0508_),
    .A1(_0510_),
    .S(_0968_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(_0507_),
    .A1(_0511_),
    .S(_0989_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(\L[9] ),
    .A1(net46),
    .S(_1114_),
    .X(_0513_));
 sky130_fd_sc_hd__xor2_2 _2588_ (.A(_0512_),
    .B(_0513_),
    .X(net170));
 sky130_fd_sc_hd__or3_1 _2589_ (.A(_0251_),
    .B(_0253_),
    .C(_0278_),
    .X(_0514_));
 sky130_fd_sc_hd__a21oi_1 _2590_ (.A1(_0222_),
    .A2(_0279_),
    .B1(_0209_),
    .Y(_0515_));
 sky130_fd_sc_hd__a2bb2o_1 _2591_ (.A1_N(_0280_),
    .A2_N(_0283_),
    .B1(_0514_),
    .B2(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__a221o_1 _2592_ (.A1(_0210_),
    .A2(_0436_),
    .B1(_0441_),
    .B2(_0288_),
    .C1(_0265_),
    .X(_0517_));
 sky130_fd_sc_hd__o21a_1 _2593_ (.A1(_0285_),
    .A2(_0516_),
    .B1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__a21bo_1 _2594_ (.A1(_0287_),
    .A2(_0283_),
    .B1_N(_0249_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _2595_ (.A(_0249_),
    .B(_0209_),
    .X(_0520_));
 sky130_fd_sc_hd__a21bo_1 _2596_ (.A1(_0248_),
    .A2(_0444_),
    .B1_N(_0441_),
    .X(_0521_));
 sky130_fd_sc_hd__a32o_1 _2597_ (.A1(_0285_),
    .A2(_0519_),
    .A3(_0520_),
    .B1(_0266_),
    .B2(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__inv_2 _2598_ (.A(_0277_),
    .Y(_0523_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(_0518_),
    .A1(_0522_),
    .S(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(\L[8] ),
    .A1(net60),
    .S(_1114_),
    .X(_0525_));
 sky130_fd_sc_hd__xor2_2 _2601_ (.A(_0524_),
    .B(_0525_),
    .X(net184));
 sky130_fd_sc_hd__o211a_1 _2602_ (.A1(_0712_),
    .A2(_0847_),
    .B1(_0807_),
    .C1(_0814_),
    .X(_0526_));
 sky130_fd_sc_hd__a21oi_1 _2603_ (.A1(_0785_),
    .A2(_0784_),
    .B1(_0712_),
    .Y(_0527_));
 sky130_fd_sc_hd__a221o_1 _2604_ (.A1(_0813_),
    .A2(_0784_),
    .B1(_0786_),
    .B2(_0527_),
    .C1(_0807_),
    .X(_0528_));
 sky130_fd_sc_hd__or2b_1 _2605_ (.A(_0845_),
    .B_N(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__o2bb2a_1 _2606_ (.A1_N(_0783_),
    .A2_N(_0784_),
    .B1(_0849_),
    .B2(_0785_),
    .X(_0530_));
 sky130_fd_sc_hd__o2bb2a_1 _2607_ (.A1_N(_0786_),
    .A2_N(_0527_),
    .B1(_0530_),
    .B2(_0812_),
    .X(_0531_));
 sky130_fd_sc_hd__o21ai_1 _2608_ (.A1(_0808_),
    .A2(_0531_),
    .B1(_0528_),
    .Y(_0532_));
 sky130_fd_sc_hd__a2bb2o_1 _2609_ (.A1_N(_0526_),
    .A2_N(_0529_),
    .B1(_0532_),
    .B2(_0845_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_4 _2610_ (.A0(\L[7] ),
    .A1(net51),
    .S(_0392_),
    .X(_0534_));
 sky130_fd_sc_hd__xnor2_2 _2611_ (.A(_0533_),
    .B(_0534_),
    .Y(net175));
 sky130_fd_sc_hd__o21a_1 _2612_ (.A1(_1095_),
    .A2(_1091_),
    .B1(_1061_),
    .X(_0535_));
 sky130_fd_sc_hd__xnor2_1 _2613_ (.A(_1101_),
    .B(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__nor2_1 _2614_ (.A(_1086_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__a21o_1 _2615_ (.A1(_1086_),
    .A2(_0536_),
    .B1(_1017_),
    .X(_0538_));
 sky130_fd_sc_hd__a211oi_1 _2616_ (.A1(_1073_),
    .A2(_1062_),
    .B1(_0415_),
    .C1(_1098_),
    .Y(_0539_));
 sky130_fd_sc_hd__a311oi_1 _2617_ (.A1(_1098_),
    .A2(_1109_),
    .A3(_1110_),
    .B1(_0539_),
    .C1(_1101_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _2618_ (.A(_1098_),
    .B(_1092_),
    .Y(_0541_));
 sky130_fd_sc_hd__nor2_1 _2619_ (.A(_1095_),
    .B(_1074_),
    .Y(_0542_));
 sky130_fd_sc_hd__a211o_1 _2620_ (.A1(_1095_),
    .A2(_1091_),
    .B1(_1098_),
    .C1(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__a31o_1 _2621_ (.A1(_1101_),
    .A2(_0541_),
    .A3(_0543_),
    .B1(_1018_),
    .X(_0544_));
 sky130_fd_sc_hd__o22a_2 _2622_ (.A1(_0537_),
    .A2(_0538_),
    .B1(_0540_),
    .B2(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_2 _2623_ (.A0(\L[6] ),
    .A1(net42),
    .S(_0392_),
    .X(_0546_));
 sky130_fd_sc_hd__xnor2_4 _2624_ (.A(_0545_),
    .B(_0546_),
    .Y(net166));
 sky130_fd_sc_hd__mux2_1 _2625_ (.A0(_0346_),
    .A1(_0348_),
    .S(_0086_),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_1 _2626_ (.A(_0088_),
    .B(_0098_),
    .Y(_0548_));
 sky130_fd_sc_hd__and2b_1 _2627_ (.A_N(_0090_),
    .B(_0342_),
    .X(_0549_));
 sky130_fd_sc_hd__or3_1 _2628_ (.A(_0086_),
    .B(_0548_),
    .C(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__a31oi_1 _2629_ (.A1(_0086_),
    .A2(_0091_),
    .A3(_0432_),
    .B1(_0076_),
    .Y(_0551_));
 sky130_fd_sc_hd__a22o_1 _2630_ (.A1(_0076_),
    .A2(_0547_),
    .B1(_0550_),
    .B2(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_2 _2631_ (.A0(\L[5] ),
    .A1(net33),
    .S(_0392_),
    .X(_0553_));
 sky130_fd_sc_hd__xnor2_2 _2632_ (.A(_0552_),
    .B(_0553_),
    .Y(net157));
 sky130_fd_sc_hd__inv_2 _2633_ (.A(_0360_),
    .Y(_0554_));
 sky130_fd_sc_hd__o22a_1 _2634_ (.A1(_0361_),
    .A2(_0554_),
    .B1(_0483_),
    .B2(_0357_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _2635_ (.A(_1200_),
    .B(_0360_),
    .Y(_0556_));
 sky130_fd_sc_hd__o21a_1 _2636_ (.A1(_1203_),
    .A2(_1205_),
    .B1(_0360_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _2637_ (.A0(_0556_),
    .A1(_0557_),
    .S(_1194_),
    .X(_0558_));
 sky130_fd_sc_hd__nand2_1 _2638_ (.A(_1202_),
    .B(_1193_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand3_1 _2639_ (.A(_1204_),
    .B(_1206_),
    .C(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__o21ai_1 _2640_ (.A1(_0358_),
    .A2(_0559_),
    .B1(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__mux2_1 _2641_ (.A0(_1168_),
    .A1(_1206_),
    .S(_0559_),
    .X(_0562_));
 sky130_fd_sc_hd__and2_1 _2642_ (.A(_0562_),
    .B(_0560_),
    .X(_0563_));
 sky130_fd_sc_hd__mux4_2 _2643_ (.A0(_0555_),
    .A1(_0558_),
    .A2(_0561_),
    .A3(_0563_),
    .S0(_1130_),
    .S1(_1212_),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(\L[4] ),
    .A1(net25),
    .S(_0605_),
    .X(_0565_));
 sky130_fd_sc_hd__xnor2_2 _2645_ (.A(_0564_),
    .B(_0565_),
    .Y(net149));
 sky130_fd_sc_hd__or3_1 _2646_ (.A(_0255_),
    .B(_0284_),
    .C(_0292_),
    .X(_0566_));
 sky130_fd_sc_hd__o311a_1 _2647_ (.A1(_0252_),
    .A2(_0254_),
    .A3(_0210_),
    .B1(_0566_),
    .C1(_0285_),
    .X(_0567_));
 sky130_fd_sc_hd__or2_1 _2648_ (.A(_0222_),
    .B(_0279_),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_1 _2649_ (.A(_0222_),
    .B(_0282_),
    .Y(_0569_));
 sky130_fd_sc_hd__a21o_1 _2650_ (.A1(_0568_),
    .A2(_0569_),
    .B1(_0255_),
    .X(_0570_));
 sky130_fd_sc_hd__a21oi_1 _2651_ (.A1(_0520_),
    .A2(_0570_),
    .B1(_0285_),
    .Y(_0571_));
 sky130_fd_sc_hd__o21a_1 _2652_ (.A1(_0252_),
    .A2(_0448_),
    .B1(_0210_),
    .X(_0572_));
 sky130_fd_sc_hd__a211oi_1 _2653_ (.A1(_0514_),
    .A2(_0515_),
    .B1(_0572_),
    .C1(_0265_),
    .Y(_0573_));
 sky130_fd_sc_hd__a21o_1 _2654_ (.A1(_0248_),
    .A2(_0287_),
    .B1(_0210_),
    .X(_0574_));
 sky130_fd_sc_hd__a31o_1 _2655_ (.A1(_0265_),
    .A2(_0570_),
    .A3(_0574_),
    .B1(_0277_),
    .X(_0575_));
 sky130_fd_sc_hd__o32a_2 _2656_ (.A1(_0523_),
    .A2(_0567_),
    .A3(_0571_),
    .B1(_0573_),
    .B2(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_2 _2657_ (.A0(\L[3] ),
    .A1(net16),
    .S(_1114_),
    .X(_0577_));
 sky130_fd_sc_hd__xor2_4 _2658_ (.A(_0576_),
    .B(_0577_),
    .X(net140));
 sky130_fd_sc_hd__and3_1 _2659_ (.A(_1249_),
    .B(_1262_),
    .C(_0377_),
    .X(_0578_));
 sky130_fd_sc_hd__o211a_1 _2660_ (.A1(_1292_),
    .A2(_1248_),
    .B1(_1296_),
    .C1(_1289_),
    .X(_0579_));
 sky130_fd_sc_hd__and4_1 _2661_ (.A(_1284_),
    .B(_1285_),
    .C(_1228_),
    .D(_1229_),
    .X(_0580_));
 sky130_fd_sc_hd__a32o_1 _2662_ (.A1(_1295_),
    .A2(_1243_),
    .A3(_1248_),
    .B1(_0580_),
    .B2(_0385_),
    .X(_0581_));
 sky130_fd_sc_hd__nor2_1 _2663_ (.A(_1262_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__a21o_1 _2664_ (.A1(_1262_),
    .A2(_0581_),
    .B1(_1272_),
    .X(_0583_));
 sky130_fd_sc_hd__o32a_1 _2665_ (.A1(_1298_),
    .A2(_0578_),
    .A3(_0579_),
    .B1(_0582_),
    .B2(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__a21oi_1 _2666_ (.A1(_0381_),
    .A2(_0382_),
    .B1(_1296_),
    .Y(_0585_));
 sky130_fd_sc_hd__a21o_1 _2667_ (.A1(_0381_),
    .A2(_0376_),
    .B1(_1298_),
    .X(_0586_));
 sky130_fd_sc_hd__nand2_1 _2668_ (.A(_1292_),
    .B(_1243_),
    .Y(_0587_));
 sky130_fd_sc_hd__or2_1 _2669_ (.A(_1292_),
    .B(_1243_),
    .X(_0588_));
 sky130_fd_sc_hd__a21oi_1 _2670_ (.A1(_0587_),
    .A2(_0588_),
    .B1(_1296_),
    .Y(_0589_));
 sky130_fd_sc_hd__a31o_1 _2671_ (.A1(_1248_),
    .A2(_1296_),
    .A3(_0587_),
    .B1(_1272_),
    .X(_0590_));
 sky130_fd_sc_hd__o22a_1 _2672_ (.A1(_0585_),
    .A2(_0586_),
    .B1(_0589_),
    .B2(_0590_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_2 _2673_ (.A0(_0584_),
    .A1(_0591_),
    .S(_0005_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_2 _2674_ (.A0(\L[2] ),
    .A1(net7),
    .S(_0605_),
    .X(_0593_));
 sky130_fd_sc_hd__xnor2_4 _2675_ (.A(_0592_),
    .B(_0593_),
    .Y(net131));
 sky130_fd_sc_hd__mux2_1 _2676_ (.A0(_0500_),
    .A1(_0497_),
    .S(_0122_),
    .X(_0594_));
 sky130_fd_sc_hd__o21ai_1 _2677_ (.A1(_0122_),
    .A2(_0493_),
    .B1(_0111_),
    .Y(_0595_));
 sky130_fd_sc_hd__and2_1 _2678_ (.A(_0122_),
    .B(_0492_),
    .X(_0596_));
 sky130_fd_sc_hd__o2bb2a_2 _2679_ (.A1_N(_0489_),
    .A2_N(_0594_),
    .B1(_0595_),
    .B2(_0596_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _2680_ (.A0(\L[1] ),
    .A1(net62),
    .S(_1114_),
    .X(_0598_));
 sky130_fd_sc_hd__xor2_2 _2681_ (.A(_0597_),
    .B(_0598_),
    .X(net186));
 sky130_fd_sc_hd__dfxtp_1 _2682_ (.CLK(clknet_3_4__leaf_clk),
    .D(net178),
    .Q(\L[32] ));
 sky130_fd_sc_hd__dfxtp_1 _2683_ (.CLK(clknet_3_6__leaf_clk),
    .D(net169),
    .Q(\L[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2684_ (.CLK(clknet_3_5__leaf_clk),
    .D(net161),
    .Q(\L[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2685_ (.CLK(clknet_3_0__leaf_clk),
    .D(net152),
    .Q(\L[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2686_ (.CLK(clknet_3_3__leaf_clk),
    .D(net143),
    .Q(\L[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2687_ (.CLK(clknet_3_4__leaf_clk),
    .D(net134),
    .Q(\L[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2688_ (.CLK(clknet_3_5__leaf_clk),
    .D(net189),
    .Q(\L[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2689_ (.CLK(clknet_3_4__leaf_clk),
    .D(net137),
    .Q(\L[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2690_ (.CLK(clknet_3_2__leaf_clk),
    .D(net180),
    .Q(\L[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2691_ (.CLK(clknet_3_5__leaf_clk),
    .D(net172),
    .Q(\L[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2692_ (.CLK(clknet_3_6__leaf_clk),
    .D(net163),
    .Q(\L[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2693_ (.CLK(clknet_3_4__leaf_clk),
    .D(net154),
    .Q(\L[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2694_ (.CLK(clknet_3_6__leaf_clk),
    .D(net145),
    .Q(\L[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2695_ (.CLK(clknet_3_1__leaf_clk),
    .D(net136),
    .Q(\L[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2696_ (.CLK(clknet_3_3__leaf_clk),
    .D(net128),
    .Q(\L[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2697_ (.CLK(clknet_3_7__leaf_clk),
    .D(net159),
    .Q(\L[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2698_ (.CLK(clknet_3_3__leaf_clk),
    .D(net183),
    .Q(\L[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2699_ (.CLK(clknet_3_4__leaf_clk),
    .D(net174),
    .Q(\L[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2700_ (.CLK(clknet_3_0__leaf_clk),
    .D(net165),
    .Q(\L[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2701_ (.CLK(clknet_3_2__leaf_clk),
    .D(net156),
    .Q(\L[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2702_ (.CLK(clknet_3_0__leaf_clk),
    .D(net147),
    .Q(\L[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2703_ (.CLK(clknet_3_7__leaf_clk),
    .D(net139),
    .Q(\L[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2704_ (.CLK(clknet_3_2__leaf_clk),
    .D(net130),
    .Q(\L[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2705_ (.CLK(clknet_3_3__leaf_clk),
    .D(net181),
    .Q(\L[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2706_ (.CLK(clknet_3_1__leaf_clk),
    .D(net185),
    .Q(\L[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2707_ (.CLK(clknet_3_3__leaf_clk),
    .D(net176),
    .Q(\L[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2708_ (.CLK(clknet_3_2__leaf_clk),
    .D(net167),
    .Q(\L[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2709_ (.CLK(clknet_3_7__leaf_clk),
    .D(net158),
    .Q(\L[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2710_ (.CLK(clknet_3_2__leaf_clk),
    .D(net150),
    .Q(\L[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2711_ (.CLK(clknet_3_5__leaf_clk),
    .D(net141),
    .Q(\L[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2712_ (.CLK(clknet_3_6__leaf_clk),
    .D(net132),
    .Q(\L[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2713_ (.CLK(clknet_3_4__leaf_clk),
    .D(net187),
    .Q(\L[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2714_ (.CLK(clknet_3_4__leaf_clk),
    .D(net177),
    .Q(\R[32] ));
 sky130_fd_sc_hd__dfxtp_1 _2715_ (.CLK(clknet_3_6__leaf_clk),
    .D(net168),
    .Q(\R[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2716_ (.CLK(clknet_3_7__leaf_clk),
    .D(net160),
    .Q(\R[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2717_ (.CLK(clknet_3_1__leaf_clk),
    .D(net151),
    .Q(\R[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2718_ (.CLK(clknet_3_2__leaf_clk),
    .D(net142),
    .Q(\R[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2719_ (.CLK(clknet_3_7__leaf_clk),
    .D(net133),
    .Q(\R[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2720_ (.CLK(clknet_3_7__leaf_clk),
    .D(net188),
    .Q(\R[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2721_ (.CLK(clknet_3_4__leaf_clk),
    .D(net126),
    .Q(\R[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2722_ (.CLK(clknet_3_2__leaf_clk),
    .D(net179),
    .Q(\R[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2723_ (.CLK(clknet_3_7__leaf_clk),
    .D(net171),
    .Q(\R[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2724_ (.CLK(clknet_3_7__leaf_clk),
    .D(net162),
    .Q(\R[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2725_ (.CLK(clknet_3_4__leaf_clk),
    .D(net153),
    .Q(\R[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2726_ (.CLK(clknet_3_6__leaf_clk),
    .D(net144),
    .Q(\R[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2727_ (.CLK(clknet_3_1__leaf_clk),
    .D(net135),
    .Q(\R[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2728_ (.CLK(clknet_3_7__leaf_clk),
    .D(net127),
    .Q(\R[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2729_ (.CLK(clknet_3_7__leaf_clk),
    .D(net148),
    .Q(\R[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2730_ (.CLK(clknet_3_6__leaf_clk),
    .D(net182),
    .Q(\R[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2731_ (.CLK(clknet_3_3__leaf_clk),
    .D(net173),
    .Q(\R[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2732_ (.CLK(clknet_3_1__leaf_clk),
    .D(net164),
    .Q(\R[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2733_ (.CLK(clknet_3_1__leaf_clk),
    .D(net155),
    .Q(\R[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2734_ (.CLK(clknet_3_7__leaf_clk),
    .D(net146),
    .Q(\R[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2735_ (.CLK(clknet_3_4__leaf_clk),
    .D(net138),
    .Q(\R[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2736_ (.CLK(clknet_3_3__leaf_clk),
    .D(net129),
    .Q(\R[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2737_ (.CLK(clknet_3_7__leaf_clk),
    .D(net170),
    .Q(\R[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2738_ (.CLK(clknet_3_2__leaf_clk),
    .D(net184),
    .Q(\R[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2739_ (.CLK(clknet_3_0__leaf_clk),
    .D(net175),
    .Q(\R[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2740_ (.CLK(clknet_3_0__leaf_clk),
    .D(net166),
    .Q(\R[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2741_ (.CLK(clknet_3_5__leaf_clk),
    .D(net157),
    .Q(\R[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2742_ (.CLK(clknet_3_6__leaf_clk),
    .D(net149),
    .Q(\R[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2743_ (.CLK(clknet_3_5__leaf_clk),
    .D(net140),
    .Q(\R[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2744_ (.CLK(clknet_3_6__leaf_clk),
    .D(net131),
    .Q(\R[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2745_ (.CLK(clknet_3_4__leaf_clk),
    .D(net186),
    .Q(\R[1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\L[10] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\L[19] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\R[15] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\L[32] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\L[29] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\L[25] ),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(decrypt),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(desIn[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input100 (.A(key[40]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(key[41]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 input102 (.A(key[42]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(key[43]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(key[44]),
    .X(net104));
 sky130_fd_sc_hd__buf_2 input105 (.A(key[45]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(key[46]),
    .X(net106));
 sky130_fd_sc_hd__buf_2 input107 (.A(key[47]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(key[48]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(key[49]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(desIn[18]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input110 (.A(key[4]),
    .X(net110));
 sky130_fd_sc_hd__buf_2 input111 (.A(key[50]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 input112 (.A(key[51]),
    .X(net112));
 sky130_fd_sc_hd__buf_2 input113 (.A(key[52]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(key[53]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(key[54]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 input116 (.A(key[55]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 input117 (.A(key[5]),
    .X(net117));
 sky130_fd_sc_hd__buf_2 input118 (.A(key[6]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(key[7]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(desIn[19]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input120 (.A(key[8]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(key[9]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 input122 (.A(roundSel[0]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 input123 (.A(roundSel[1]),
    .X(net123));
 sky130_fd_sc_hd__buf_4 input124 (.A(roundSel[2]),
    .X(net124));
 sky130_fd_sc_hd__buf_1 input125 (.A(roundSel[3]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input13 (.A(desIn[1]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(desIn[20]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(desIn[21]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(desIn[22]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(desIn[23]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(desIn[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(desIn[25]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(desIn[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(desIn[26]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(desIn[27]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(desIn[28]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(desIn[29]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(desIn[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(desIn[30]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(desIn[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(desIn[32]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(desIn[33]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(desIn[34]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(desIn[10]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(desIn[35]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(desIn[36]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(desIn[37]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(desIn[38]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(desIn[39]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(desIn[3]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(desIn[40]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(desIn[41]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(desIn[42]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(desIn[43]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(desIn[11]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(desIn[44]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(desIn[45]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(desIn[46]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(desIn[47]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(desIn[48]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(desIn[49]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(desIn[4]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(desIn[50]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(desIn[51]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(desIn[52]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(desIn[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(desIn[53]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(desIn[54]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(desIn[55]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(desIn[56]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(desIn[57]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(desIn[58]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(desIn[59]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(desIn[5]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input58 (.A(desIn[60]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(desIn[61]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(desIn[13]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(desIn[62]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(desIn[63]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(desIn[6]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(desIn[7]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(desIn[8]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(desIn[9]),
    .X(net65));
 sky130_fd_sc_hd__buf_2 input66 (.A(key[0]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(key[10]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(key[11]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(key[12]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(desIn[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(key[13]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(key[14]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 input72 (.A(key[15]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(key[16]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 input74 (.A(key[17]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_4 input75 (.A(key[18]),
    .X(net75));
 sky130_fd_sc_hd__buf_2 input76 (.A(key[19]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 input77 (.A(key[1]),
    .X(net77));
 sky130_fd_sc_hd__buf_2 input78 (.A(key[20]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(key[21]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input8 (.A(desIn[15]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input80 (.A(key[22]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(key[23]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 input82 (.A(key[24]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(key[25]),
    .X(net83));
 sky130_fd_sc_hd__buf_2 input84 (.A(key[26]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(key[27]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input86 (.A(key[28]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(key[29]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(key[2]),
    .X(net88));
 sky130_fd_sc_hd__buf_2 input89 (.A(key[30]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(desIn[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input90 (.A(key[31]),
    .X(net90));
 sky130_fd_sc_hd__buf_2 input91 (.A(key[32]),
    .X(net91));
 sky130_fd_sc_hd__buf_2 input92 (.A(key[33]),
    .X(net92));
 sky130_fd_sc_hd__buf_2 input93 (.A(key[34]),
    .X(net93));
 sky130_fd_sc_hd__buf_4 input94 (.A(key[35]),
    .X(net94));
 sky130_fd_sc_hd__buf_4 input95 (.A(key[36]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 input96 (.A(key[37]),
    .X(net96));
 sky130_fd_sc_hd__buf_2 input97 (.A(key[38]),
    .X(net97));
 sky130_fd_sc_hd__buf_2 input98 (.A(key[39]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input99 (.A(key[3]),
    .X(net99));
 sky130_fd_sc_hd__buf_4 max_cap190 (.A(_0600_),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net126),
    .X(desOut[0]));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net127),
    .X(desOut[10]));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net128),
    .X(desOut[11]));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net129),
    .X(desOut[12]));
 sky130_fd_sc_hd__clkbuf_4 output130 (.A(net130),
    .X(desOut[13]));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net131),
    .X(desOut[14]));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net132),
    .X(desOut[15]));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net133),
    .X(desOut[16]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(desOut[17]));
 sky130_fd_sc_hd__clkbuf_4 output135 (.A(net135),
    .X(desOut[18]));
 sky130_fd_sc_hd__clkbuf_4 output136 (.A(net136),
    .X(desOut[19]));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net137),
    .X(desOut[1]));
 sky130_fd_sc_hd__clkbuf_4 output138 (.A(net138),
    .X(desOut[20]));
 sky130_fd_sc_hd__clkbuf_4 output139 (.A(net139),
    .X(desOut[21]));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net140),
    .X(desOut[22]));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net141),
    .X(desOut[23]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(desOut[24]));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net143),
    .X(desOut[25]));
 sky130_fd_sc_hd__clkbuf_4 output144 (.A(net144),
    .X(desOut[26]));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net145),
    .X(desOut[27]));
 sky130_fd_sc_hd__clkbuf_4 output146 (.A(net146),
    .X(desOut[28]));
 sky130_fd_sc_hd__clkbuf_4 output147 (.A(net147),
    .X(desOut[29]));
 sky130_fd_sc_hd__clkbuf_4 output148 (.A(net148),
    .X(desOut[2]));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net149),
    .X(desOut[30]));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net150),
    .X(desOut[31]));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net151),
    .X(desOut[32]));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net152),
    .X(desOut[33]));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net153),
    .X(desOut[34]));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net154),
    .X(desOut[35]));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net155),
    .X(desOut[36]));
 sky130_fd_sc_hd__clkbuf_4 output156 (.A(net156),
    .X(desOut[37]));
 sky130_fd_sc_hd__clkbuf_4 output157 (.A(net157),
    .X(desOut[38]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(desOut[39]));
 sky130_fd_sc_hd__clkbuf_4 output159 (.A(net159),
    .X(desOut[3]));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net160),
    .X(desOut[40]));
 sky130_fd_sc_hd__clkbuf_4 output161 (.A(net161),
    .X(desOut[41]));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net162),
    .X(desOut[42]));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net163),
    .X(desOut[43]));
 sky130_fd_sc_hd__clkbuf_4 output164 (.A(net164),
    .X(desOut[44]));
 sky130_fd_sc_hd__clkbuf_4 output165 (.A(net165),
    .X(desOut[45]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(desOut[46]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(desOut[47]));
 sky130_fd_sc_hd__clkbuf_4 output168 (.A(net168),
    .X(desOut[48]));
 sky130_fd_sc_hd__clkbuf_4 output169 (.A(net169),
    .X(desOut[49]));
 sky130_fd_sc_hd__clkbuf_4 output170 (.A(net170),
    .X(desOut[4]));
 sky130_fd_sc_hd__clkbuf_4 output171 (.A(net171),
    .X(desOut[50]));
 sky130_fd_sc_hd__clkbuf_4 output172 (.A(net172),
    .X(desOut[51]));
 sky130_fd_sc_hd__clkbuf_4 output173 (.A(net173),
    .X(desOut[52]));
 sky130_fd_sc_hd__clkbuf_4 output174 (.A(net174),
    .X(desOut[53]));
 sky130_fd_sc_hd__clkbuf_4 output175 (.A(net175),
    .X(desOut[54]));
 sky130_fd_sc_hd__clkbuf_4 output176 (.A(net176),
    .X(desOut[55]));
 sky130_fd_sc_hd__clkbuf_4 output177 (.A(net177),
    .X(desOut[56]));
 sky130_fd_sc_hd__clkbuf_4 output178 (.A(net178),
    .X(desOut[57]));
 sky130_fd_sc_hd__clkbuf_4 output179 (.A(net179),
    .X(desOut[58]));
 sky130_fd_sc_hd__clkbuf_4 output180 (.A(net180),
    .X(desOut[59]));
 sky130_fd_sc_hd__clkbuf_4 output181 (.A(net181),
    .X(desOut[5]));
 sky130_fd_sc_hd__clkbuf_4 output182 (.A(net182),
    .X(desOut[60]));
 sky130_fd_sc_hd__clkbuf_4 output183 (.A(net183),
    .X(desOut[61]));
 sky130_fd_sc_hd__clkbuf_4 output184 (.A(net184),
    .X(desOut[62]));
 sky130_fd_sc_hd__clkbuf_4 output185 (.A(net185),
    .X(desOut[63]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(desOut[6]));
 sky130_fd_sc_hd__clkbuf_4 output187 (.A(net187),
    .X(desOut[7]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(desOut[8]));
 sky130_fd_sc_hd__clkbuf_4 output189 (.A(net189),
    .X(desOut[9]));
endmodule

