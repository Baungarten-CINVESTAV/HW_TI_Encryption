VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO des_Trojan
  CLASS BLOCK ;
  FOREIGN des_Trojan ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 496.000 210.840 500.000 211.440 ;
    END
  END clk
  PIN decrypt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END decrypt
  PIN desIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END desIn[0]
  PIN desIn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END desIn[10]
  PIN desIn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 360.440 500.000 361.040 ;
    END
  END desIn[11]
  PIN desIn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END desIn[12]
  PIN desIn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END desIn[13]
  PIN desIn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END desIn[14]
  PIN desIn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 142.840 500.000 143.440 ;
    END
  END desIn[15]
  PIN desIn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 421.910 496.000 422.190 500.000 ;
    END
  END desIn[16]
  PIN desIn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END desIn[17]
  PIN desIn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END desIn[18]
  PIN desIn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 122.440 500.000 123.040 ;
    END
  END desIn[19]
  PIN desIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END desIn[1]
  PIN desIn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END desIn[20]
  PIN desIn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END desIn[21]
  PIN desIn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 496.000 42.230 500.000 ;
    END
  END desIn[22]
  PIN desIn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 496.000 103.410 500.000 ;
    END
  END desIn[23]
  PIN desIn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 374.040 500.000 374.640 ;
    END
  END desIn[24]
  PIN desIn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 267.350 496.000 267.630 500.000 ;
    END
  END desIn[25]
  PIN desIn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 295.840 500.000 296.440 ;
    END
  END desIn[26]
  PIN desIn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END desIn[27]
  PIN desIn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 289.890 496.000 290.170 500.000 ;
    END
  END desIn[28]
  PIN desIn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END desIn[29]
  PIN desIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END desIn[2]
  PIN desIn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 384.240 500.000 384.840 ;
    END
  END desIn[30]
  PIN desIn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 68.040 500.000 68.640 ;
    END
  END desIn[31]
  PIN desIn[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END desIn[32]
  PIN desIn[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 318.870 496.000 319.150 500.000 ;
    END
  END desIn[33]
  PIN desIn[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 496.000 71.210 500.000 ;
    END
  END desIn[34]
  PIN desIn[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END desIn[35]
  PIN desIn[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END desIn[36]
  PIN desIn[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END desIn[37]
  PIN desIn[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END desIn[38]
  PIN desIn[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 438.640 500.000 439.240 ;
    END
  END desIn[39]
  PIN desIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 493.040 500.000 493.640 ;
    END
  END desIn[3]
  PIN desIn[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 265.240 500.000 265.840 ;
    END
  END desIn[40]
  PIN desIn[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 257.690 496.000 257.970 500.000 ;
    END
  END desIn[41]
  PIN desIn[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 434.790 496.000 435.070 500.000 ;
    END
  END desIn[42]
  PIN desIn[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END desIn[43]
  PIN desIn[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END desIn[44]
  PIN desIn[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END desIn[45]
  PIN desIn[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 463.770 496.000 464.050 500.000 ;
    END
  END desIn[46]
  PIN desIn[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 57.840 500.000 58.440 ;
    END
  END desIn[47]
  PIN desIn[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 23.840 500.000 24.440 ;
    END
  END desIn[48]
  PIN desIn[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END desIn[49]
  PIN desIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END desIn[4]
  PIN desIn[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END desIn[50]
  PIN desIn[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 156.440 500.000 157.040 ;
    END
  END desIn[51]
  PIN desIn[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 496.000 174.250 500.000 ;
    END
  END desIn[52]
  PIN desIn[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 392.930 496.000 393.210 500.000 ;
    END
  END desIn[53]
  PIN desIn[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END desIn[54]
  PIN desIn[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 496.000 154.930 500.000 ;
    END
  END desIn[55]
  PIN desIn[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 496.000 187.130 500.000 ;
    END
  END desIn[56]
  PIN desIn[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END desIn[57]
  PIN desIn[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 88.440 500.000 89.040 ;
    END
  END desIn[58]
  PIN desIn[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 196.510 496.000 196.790 500.000 ;
    END
  END desIn[59]
  PIN desIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 448.840 500.000 449.440 ;
    END
  END desIn[5]
  PIN desIn[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END desIn[60]
  PIN desIn[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END desIn[61]
  PIN desIn[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END desIn[62]
  PIN desIn[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 241.440 500.000 242.040 ;
    END
  END desIn[63]
  PIN desIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END desIn[6]
  PIN desIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END desIn[7]
  PIN desIn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 44.240 500.000 44.840 ;
    END
  END desIn[8]
  PIN desIn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 238.370 496.000 238.650 500.000 ;
    END
  END desIn[9]
  PIN desOut_ff[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 454.110 496.000 454.390 500.000 ;
    END
  END desOut_ff[0]
  PIN desOut_ff[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 469.240 500.000 469.840 ;
    END
  END desOut_ff[10]
  PIN desOut_ff[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 444.450 496.000 444.730 500.000 ;
    END
  END desOut_ff[11]
  PIN desOut_ff[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END desOut_ff[12]
  PIN desOut_ff[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END desOut_ff[13]
  PIN desOut_ff[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 496.000 93.750 500.000 ;
    END
  END desOut_ff[14]
  PIN desOut_ff[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 402.590 496.000 402.870 500.000 ;
    END
  END desOut_ff[15]
  PIN desOut_ff[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END desOut_ff[16]
  PIN desOut_ff[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END desOut_ff[17]
  PIN desOut_ff[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END desOut_ff[18]
  PIN desOut_ff[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.330 496.000 135.610 500.000 ;
    END
  END desOut_ff[19]
  PIN desOut_ff[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END desOut_ff[1]
  PIN desOut_ff[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 251.640 500.000 252.240 ;
    END
  END desOut_ff[20]
  PIN desOut_ff[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END desOut_ff[21]
  PIN desOut_ff[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END desOut_ff[22]
  PIN desOut_ff[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 51.610 496.000 51.890 500.000 ;
    END
  END desOut_ff[23]
  PIN desOut_ff[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.310 496.000 164.590 500.000 ;
    END
  END desOut_ff[24]
  PIN desOut_ff[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 19.410 496.000 19.690 500.000 ;
    END
  END desOut_ff[25]
  PIN desOut_ff[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 329.840 500.000 330.440 ;
    END
  END desOut_ff[26]
  PIN desOut_ff[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END desOut_ff[27]
  PIN desOut_ff[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END desOut_ff[28]
  PIN desOut_ff[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END desOut_ff[29]
  PIN desOut_ff[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 404.640 500.000 405.240 ;
    END
  END desOut_ff[2]
  PIN desOut_ff[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END desOut_ff[30]
  PIN desOut_ff[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END desOut_ff[31]
  PIN desOut_ff[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 383.270 496.000 383.550 500.000 ;
    END
  END desOut_ff[32]
  PIN desOut_ff[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 13.640 500.000 14.240 ;
    END
  END desOut_ff[33]
  PIN desOut_ff[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END desOut_ff[34]
  PIN desOut_ff[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 496.000 3.440 500.000 4.040 ;
    END
  END desOut_ff[35]
  PIN desOut_ff[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END desOut_ff[36]
  PIN desOut_ff[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END desOut_ff[37]
  PIN desOut_ff[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 496.000 275.440 500.000 276.040 ;
    END
  END desOut_ff[38]
  PIN desOut_ff[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 370.390 496.000 370.670 500.000 ;
    END
  END desOut_ff[39]
  PIN desOut_ff[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END desOut_ff[3]
  PIN desOut_ff[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.990 496.000 145.270 500.000 ;
    END
  END desOut_ff[40]
  PIN desOut_ff[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END desOut_ff[41]
  PIN desOut_ff[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 496.000 482.840 500.000 483.440 ;
    END
  END desOut_ff[42]
  PIN desOut_ff[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END desOut_ff[43]
  PIN desOut_ff[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END desOut_ff[44]
  PIN desOut_ff[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 428.440 500.000 429.040 ;
    END
  END desOut_ff[45]
  PIN desOut_ff[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END desOut_ff[46]
  PIN desOut_ff[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 176.840 500.000 177.440 ;
    END
  END desOut_ff[47]
  PIN desOut_ff[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END desOut_ff[48]
  PIN desOut_ff[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 285.640 500.000 286.240 ;
    END
  END desOut_ff[49]
  PIN desOut_ff[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END desOut_ff[4]
  PIN desOut_ff[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 309.210 496.000 309.490 500.000 ;
    END
  END desOut_ff[50]
  PIN desOut_ff[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 306.040 500.000 306.640 ;
    END
  END desOut_ff[51]
  PIN desOut_ff[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END desOut_ff[52]
  PIN desOut_ff[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END desOut_ff[53]
  PIN desOut_ff[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 206.170 496.000 206.450 500.000 ;
    END
  END desOut_ff[54]
  PIN desOut_ff[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END desOut_ff[55]
  PIN desOut_ff[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 4.000 ;
    END
  END desOut_ff[56]
  PIN desOut_ff[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 486.310 496.000 486.590 500.000 ;
    END
  END desOut_ff[57]
  PIN desOut_ff[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 197.240 500.000 197.840 ;
    END
  END desOut_ff[58]
  PIN desOut_ff[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 215.830 496.000 216.110 500.000 ;
    END
  END desOut_ff[59]
  PIN desOut_ff[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 299.550 496.000 299.830 500.000 ;
    END
  END desOut_ff[5]
  PIN desOut_ff[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 280.230 496.000 280.510 500.000 ;
    END
  END desOut_ff[60]
  PIN desOut_ff[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END desOut_ff[61]
  PIN desOut_ff[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END desOut_ff[62]
  PIN desOut_ff[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 78.240 500.000 78.840 ;
    END
  END desOut_ff[63]
  PIN desOut_ff[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END desOut_ff[6]
  PIN desOut_ff[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 414.840 500.000 415.440 ;
    END
  END desOut_ff[7]
  PIN desOut_ff[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 112.790 496.000 113.070 500.000 ;
    END
  END desOut_ff[8]
  PIN desOut_ff[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 331.750 496.000 332.030 500.000 ;
    END
  END desOut_ff[9]
  PIN finish
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END finish
  PIN init
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 132.640 500.000 133.240 ;
    END
  END init
  PIN key[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END key[0]
  PIN key[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 496.000 122.730 500.000 ;
    END
  END key[10]
  PIN key[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 221.040 500.000 221.640 ;
    END
  END key[11]
  PIN key[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 9.750 496.000 10.030 500.000 ;
    END
  END key[12]
  PIN key[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END key[13]
  PIN key[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 394.440 500.000 395.040 ;
    END
  END key[14]
  PIN key[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END key[15]
  PIN key[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END key[16]
  PIN key[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 166.640 500.000 167.240 ;
    END
  END key[17]
  PIN key[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END key[18]
  PIN key[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 34.040 500.000 34.640 ;
    END
  END key[19]
  PIN key[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 496.000 32.570 500.000 ;
    END
  END key[1]
  PIN key[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END key[20]
  PIN key[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END key[21]
  PIN key[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END key[22]
  PIN key[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 112.240 500.000 112.840 ;
    END
  END key[23]
  PIN key[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 459.040 500.000 459.640 ;
    END
  END key[24]
  PIN key[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 319.640 500.000 320.240 ;
    END
  END key[25]
  PIN key[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END key[26]
  PIN key[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END key[27]
  PIN key[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 187.040 500.000 187.640 ;
    END
  END key[28]
  PIN key[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END key[29]
  PIN key[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 350.240 500.000 350.840 ;
    END
  END key[2]
  PIN key[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 495.970 496.000 496.250 500.000 ;
    END
  END key[30]
  PIN key[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END key[31]
  PIN key[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 473.430 496.000 473.710 500.000 ;
    END
  END key[32]
  PIN key[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END key[33]
  PIN key[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END key[34]
  PIN key[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END key[35]
  PIN key[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END key[36]
  PIN key[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END key[37]
  PIN key[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END key[38]
  PIN key[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 496.000 61.550 500.000 ;
    END
  END key[39]
  PIN key[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 248.030 496.000 248.310 500.000 ;
    END
  END key[3]
  PIN key[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END key[40]
  PIN key[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END key[41]
  PIN key[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END key[42]
  PIN key[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 341.410 496.000 341.690 500.000 ;
    END
  END key[43]
  PIN key[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 228.710 496.000 228.990 500.000 ;
    END
  END key[44]
  PIN key[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END key[45]
  PIN key[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 412.250 496.000 412.530 500.000 ;
    END
  END key[46]
  PIN key[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 98.640 500.000 99.240 ;
    END
  END key[47]
  PIN key[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END key[48]
  PIN key[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END key[49]
  PIN key[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END key[4]
  PIN key[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END key[50]
  PIN key[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END key[51]
  PIN key[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 496.000 340.040 500.000 340.640 ;
    END
  END key[52]
  PIN key[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END key[53]
  PIN key[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 360.730 496.000 361.010 500.000 ;
    END
  END key[54]
  PIN key[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 351.070 496.000 351.350 500.000 ;
    END
  END key[55]
  PIN key[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 496.000 0.370 500.000 ;
    END
  END key[5]
  PIN key[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 496.000 84.090 500.000 ;
    END
  END key[6]
  PIN key[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END key[7]
  PIN key[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END key[8]
  PIN key[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END key[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 496.000 231.240 500.000 231.840 ;
    END
  END reset
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.720 10.640 191.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 369.720 10.640 371.320 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 99.720 10.640 101.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.720 10.640 281.320 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 459.720 10.640 461.320 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 0.070 10.640 496.270 487.120 ;
      LAYER met2 ;
        RECT 0.650 495.720 9.470 496.810 ;
        RECT 10.310 495.720 19.130 496.810 ;
        RECT 19.970 495.720 32.010 496.810 ;
        RECT 32.850 495.720 41.670 496.810 ;
        RECT 42.510 495.720 51.330 496.810 ;
        RECT 52.170 495.720 60.990 496.810 ;
        RECT 61.830 495.720 70.650 496.810 ;
        RECT 71.490 495.720 83.530 496.810 ;
        RECT 84.370 495.720 93.190 496.810 ;
        RECT 94.030 495.720 102.850 496.810 ;
        RECT 103.690 495.720 112.510 496.810 ;
        RECT 113.350 495.720 122.170 496.810 ;
        RECT 123.010 495.720 135.050 496.810 ;
        RECT 135.890 495.720 144.710 496.810 ;
        RECT 145.550 495.720 154.370 496.810 ;
        RECT 155.210 495.720 164.030 496.810 ;
        RECT 164.870 495.720 173.690 496.810 ;
        RECT 174.530 495.720 186.570 496.810 ;
        RECT 187.410 495.720 196.230 496.810 ;
        RECT 197.070 495.720 205.890 496.810 ;
        RECT 206.730 495.720 215.550 496.810 ;
        RECT 216.390 495.720 228.430 496.810 ;
        RECT 229.270 495.720 238.090 496.810 ;
        RECT 238.930 495.720 247.750 496.810 ;
        RECT 248.590 495.720 257.410 496.810 ;
        RECT 258.250 495.720 267.070 496.810 ;
        RECT 267.910 495.720 279.950 496.810 ;
        RECT 280.790 495.720 289.610 496.810 ;
        RECT 290.450 495.720 299.270 496.810 ;
        RECT 300.110 495.720 308.930 496.810 ;
        RECT 309.770 495.720 318.590 496.810 ;
        RECT 319.430 495.720 331.470 496.810 ;
        RECT 332.310 495.720 341.130 496.810 ;
        RECT 341.970 495.720 350.790 496.810 ;
        RECT 351.630 495.720 360.450 496.810 ;
        RECT 361.290 495.720 370.110 496.810 ;
        RECT 370.950 495.720 382.990 496.810 ;
        RECT 383.830 495.720 392.650 496.810 ;
        RECT 393.490 495.720 402.310 496.810 ;
        RECT 403.150 495.720 411.970 496.810 ;
        RECT 412.810 495.720 421.630 496.810 ;
        RECT 422.470 495.720 434.510 496.810 ;
        RECT 435.350 495.720 444.170 496.810 ;
        RECT 445.010 495.720 453.830 496.810 ;
        RECT 454.670 495.720 463.490 496.810 ;
        RECT 464.330 495.720 473.150 496.810 ;
        RECT 473.990 495.720 486.030 496.810 ;
        RECT 486.870 495.720 495.690 496.810 ;
        RECT 0.100 4.280 496.240 495.720 ;
        RECT 0.650 3.555 9.470 4.280 ;
        RECT 10.310 3.555 19.130 4.280 ;
        RECT 19.970 3.555 28.790 4.280 ;
        RECT 29.630 3.555 38.450 4.280 ;
        RECT 39.290 3.555 51.330 4.280 ;
        RECT 52.170 3.555 60.990 4.280 ;
        RECT 61.830 3.555 70.650 4.280 ;
        RECT 71.490 3.555 80.310 4.280 ;
        RECT 81.150 3.555 89.970 4.280 ;
        RECT 90.810 3.555 102.850 4.280 ;
        RECT 103.690 3.555 112.510 4.280 ;
        RECT 113.350 3.555 122.170 4.280 ;
        RECT 123.010 3.555 131.830 4.280 ;
        RECT 132.670 3.555 141.490 4.280 ;
        RECT 142.330 3.555 154.370 4.280 ;
        RECT 155.210 3.555 164.030 4.280 ;
        RECT 164.870 3.555 173.690 4.280 ;
        RECT 174.530 3.555 183.350 4.280 ;
        RECT 184.190 3.555 193.010 4.280 ;
        RECT 193.850 3.555 205.890 4.280 ;
        RECT 206.730 3.555 215.550 4.280 ;
        RECT 216.390 3.555 225.210 4.280 ;
        RECT 226.050 3.555 234.870 4.280 ;
        RECT 235.710 3.555 244.530 4.280 ;
        RECT 245.370 3.555 257.410 4.280 ;
        RECT 258.250 3.555 267.070 4.280 ;
        RECT 267.910 3.555 276.730 4.280 ;
        RECT 277.570 3.555 286.390 4.280 ;
        RECT 287.230 3.555 296.050 4.280 ;
        RECT 296.890 3.555 308.930 4.280 ;
        RECT 309.770 3.555 318.590 4.280 ;
        RECT 319.430 3.555 328.250 4.280 ;
        RECT 329.090 3.555 337.910 4.280 ;
        RECT 338.750 3.555 350.790 4.280 ;
        RECT 351.630 3.555 360.450 4.280 ;
        RECT 361.290 3.555 370.110 4.280 ;
        RECT 370.950 3.555 379.770 4.280 ;
        RECT 380.610 3.555 389.430 4.280 ;
        RECT 390.270 3.555 402.310 4.280 ;
        RECT 403.150 3.555 411.970 4.280 ;
        RECT 412.810 3.555 421.630 4.280 ;
        RECT 422.470 3.555 431.290 4.280 ;
        RECT 432.130 3.555 440.950 4.280 ;
        RECT 441.790 3.555 453.830 4.280 ;
        RECT 454.670 3.555 463.490 4.280 ;
        RECT 464.330 3.555 473.150 4.280 ;
        RECT 473.990 3.555 482.810 4.280 ;
        RECT 483.650 3.555 492.470 4.280 ;
        RECT 493.310 3.555 496.240 4.280 ;
      LAYER met3 ;
        RECT 3.990 492.640 495.600 493.505 ;
        RECT 3.990 490.640 496.000 492.640 ;
        RECT 4.400 489.240 496.000 490.640 ;
        RECT 3.990 483.840 496.000 489.240 ;
        RECT 3.990 482.440 495.600 483.840 ;
        RECT 3.990 480.440 496.000 482.440 ;
        RECT 4.400 479.040 496.000 480.440 ;
        RECT 3.990 470.240 496.000 479.040 ;
        RECT 3.990 468.840 495.600 470.240 ;
        RECT 3.990 466.840 496.000 468.840 ;
        RECT 4.400 465.440 496.000 466.840 ;
        RECT 3.990 460.040 496.000 465.440 ;
        RECT 3.990 458.640 495.600 460.040 ;
        RECT 3.990 456.640 496.000 458.640 ;
        RECT 4.400 455.240 496.000 456.640 ;
        RECT 3.990 449.840 496.000 455.240 ;
        RECT 3.990 448.440 495.600 449.840 ;
        RECT 3.990 446.440 496.000 448.440 ;
        RECT 4.400 445.040 496.000 446.440 ;
        RECT 3.990 439.640 496.000 445.040 ;
        RECT 3.990 438.240 495.600 439.640 ;
        RECT 3.990 436.240 496.000 438.240 ;
        RECT 4.400 434.840 496.000 436.240 ;
        RECT 3.990 429.440 496.000 434.840 ;
        RECT 3.990 428.040 495.600 429.440 ;
        RECT 3.990 426.040 496.000 428.040 ;
        RECT 4.400 424.640 496.000 426.040 ;
        RECT 3.990 415.840 496.000 424.640 ;
        RECT 3.990 414.440 495.600 415.840 ;
        RECT 3.990 412.440 496.000 414.440 ;
        RECT 4.400 411.040 496.000 412.440 ;
        RECT 3.990 405.640 496.000 411.040 ;
        RECT 3.990 404.240 495.600 405.640 ;
        RECT 3.990 402.240 496.000 404.240 ;
        RECT 4.400 400.840 496.000 402.240 ;
        RECT 3.990 395.440 496.000 400.840 ;
        RECT 3.990 394.040 495.600 395.440 ;
        RECT 3.990 392.040 496.000 394.040 ;
        RECT 4.400 390.640 496.000 392.040 ;
        RECT 3.990 385.240 496.000 390.640 ;
        RECT 3.990 383.840 495.600 385.240 ;
        RECT 3.990 381.840 496.000 383.840 ;
        RECT 4.400 380.440 496.000 381.840 ;
        RECT 3.990 375.040 496.000 380.440 ;
        RECT 3.990 373.640 495.600 375.040 ;
        RECT 3.990 371.640 496.000 373.640 ;
        RECT 4.400 370.240 496.000 371.640 ;
        RECT 3.990 361.440 496.000 370.240 ;
        RECT 3.990 360.040 495.600 361.440 ;
        RECT 3.990 358.040 496.000 360.040 ;
        RECT 4.400 356.640 496.000 358.040 ;
        RECT 3.990 351.240 496.000 356.640 ;
        RECT 3.990 349.840 495.600 351.240 ;
        RECT 3.990 347.840 496.000 349.840 ;
        RECT 4.400 346.440 496.000 347.840 ;
        RECT 3.990 341.040 496.000 346.440 ;
        RECT 3.990 339.640 495.600 341.040 ;
        RECT 3.990 337.640 496.000 339.640 ;
        RECT 4.400 336.240 496.000 337.640 ;
        RECT 3.990 330.840 496.000 336.240 ;
        RECT 3.990 329.440 495.600 330.840 ;
        RECT 3.990 327.440 496.000 329.440 ;
        RECT 4.400 326.040 496.000 327.440 ;
        RECT 3.990 320.640 496.000 326.040 ;
        RECT 3.990 319.240 495.600 320.640 ;
        RECT 3.990 313.840 496.000 319.240 ;
        RECT 4.400 312.440 496.000 313.840 ;
        RECT 3.990 307.040 496.000 312.440 ;
        RECT 3.990 305.640 495.600 307.040 ;
        RECT 3.990 303.640 496.000 305.640 ;
        RECT 4.400 302.240 496.000 303.640 ;
        RECT 3.990 296.840 496.000 302.240 ;
        RECT 3.990 295.440 495.600 296.840 ;
        RECT 3.990 293.440 496.000 295.440 ;
        RECT 4.400 292.040 496.000 293.440 ;
        RECT 3.990 286.640 496.000 292.040 ;
        RECT 3.990 285.240 495.600 286.640 ;
        RECT 3.990 283.240 496.000 285.240 ;
        RECT 4.400 281.840 496.000 283.240 ;
        RECT 3.990 276.440 496.000 281.840 ;
        RECT 3.990 275.040 495.600 276.440 ;
        RECT 3.990 273.040 496.000 275.040 ;
        RECT 4.400 271.640 496.000 273.040 ;
        RECT 3.990 266.240 496.000 271.640 ;
        RECT 3.990 264.840 495.600 266.240 ;
        RECT 3.990 259.440 496.000 264.840 ;
        RECT 4.400 258.040 496.000 259.440 ;
        RECT 3.990 252.640 496.000 258.040 ;
        RECT 3.990 251.240 495.600 252.640 ;
        RECT 3.990 249.240 496.000 251.240 ;
        RECT 4.400 247.840 496.000 249.240 ;
        RECT 3.990 242.440 496.000 247.840 ;
        RECT 3.990 241.040 495.600 242.440 ;
        RECT 3.990 239.040 496.000 241.040 ;
        RECT 4.400 237.640 496.000 239.040 ;
        RECT 3.990 232.240 496.000 237.640 ;
        RECT 3.990 230.840 495.600 232.240 ;
        RECT 3.990 228.840 496.000 230.840 ;
        RECT 4.400 227.440 496.000 228.840 ;
        RECT 3.990 222.040 496.000 227.440 ;
        RECT 3.990 220.640 495.600 222.040 ;
        RECT 3.990 218.640 496.000 220.640 ;
        RECT 4.400 217.240 496.000 218.640 ;
        RECT 3.990 211.840 496.000 217.240 ;
        RECT 3.990 210.440 495.600 211.840 ;
        RECT 3.990 205.040 496.000 210.440 ;
        RECT 4.400 203.640 496.000 205.040 ;
        RECT 3.990 198.240 496.000 203.640 ;
        RECT 3.990 196.840 495.600 198.240 ;
        RECT 3.990 194.840 496.000 196.840 ;
        RECT 4.400 193.440 496.000 194.840 ;
        RECT 3.990 188.040 496.000 193.440 ;
        RECT 3.990 186.640 495.600 188.040 ;
        RECT 3.990 184.640 496.000 186.640 ;
        RECT 4.400 183.240 496.000 184.640 ;
        RECT 3.990 177.840 496.000 183.240 ;
        RECT 3.990 176.440 495.600 177.840 ;
        RECT 3.990 174.440 496.000 176.440 ;
        RECT 4.400 173.040 496.000 174.440 ;
        RECT 3.990 167.640 496.000 173.040 ;
        RECT 3.990 166.240 495.600 167.640 ;
        RECT 3.990 164.240 496.000 166.240 ;
        RECT 4.400 162.840 496.000 164.240 ;
        RECT 3.990 157.440 496.000 162.840 ;
        RECT 3.990 156.040 495.600 157.440 ;
        RECT 3.990 150.640 496.000 156.040 ;
        RECT 4.400 149.240 496.000 150.640 ;
        RECT 3.990 143.840 496.000 149.240 ;
        RECT 3.990 142.440 495.600 143.840 ;
        RECT 3.990 140.440 496.000 142.440 ;
        RECT 4.400 139.040 496.000 140.440 ;
        RECT 3.990 133.640 496.000 139.040 ;
        RECT 3.990 132.240 495.600 133.640 ;
        RECT 3.990 130.240 496.000 132.240 ;
        RECT 4.400 128.840 496.000 130.240 ;
        RECT 3.990 123.440 496.000 128.840 ;
        RECT 3.990 122.040 495.600 123.440 ;
        RECT 3.990 120.040 496.000 122.040 ;
        RECT 4.400 118.640 496.000 120.040 ;
        RECT 3.990 113.240 496.000 118.640 ;
        RECT 3.990 111.840 495.600 113.240 ;
        RECT 3.990 109.840 496.000 111.840 ;
        RECT 4.400 108.440 496.000 109.840 ;
        RECT 3.990 99.640 496.000 108.440 ;
        RECT 3.990 98.240 495.600 99.640 ;
        RECT 3.990 96.240 496.000 98.240 ;
        RECT 4.400 94.840 496.000 96.240 ;
        RECT 3.990 89.440 496.000 94.840 ;
        RECT 3.990 88.040 495.600 89.440 ;
        RECT 3.990 86.040 496.000 88.040 ;
        RECT 4.400 84.640 496.000 86.040 ;
        RECT 3.990 79.240 496.000 84.640 ;
        RECT 3.990 77.840 495.600 79.240 ;
        RECT 3.990 75.840 496.000 77.840 ;
        RECT 4.400 74.440 496.000 75.840 ;
        RECT 3.990 69.040 496.000 74.440 ;
        RECT 3.990 67.640 495.600 69.040 ;
        RECT 3.990 65.640 496.000 67.640 ;
        RECT 4.400 64.240 496.000 65.640 ;
        RECT 3.990 58.840 496.000 64.240 ;
        RECT 3.990 57.440 495.600 58.840 ;
        RECT 3.990 55.440 496.000 57.440 ;
        RECT 4.400 54.040 496.000 55.440 ;
        RECT 3.990 45.240 496.000 54.040 ;
        RECT 3.990 43.840 495.600 45.240 ;
        RECT 3.990 41.840 496.000 43.840 ;
        RECT 4.400 40.440 496.000 41.840 ;
        RECT 3.990 35.040 496.000 40.440 ;
        RECT 3.990 33.640 495.600 35.040 ;
        RECT 3.990 31.640 496.000 33.640 ;
        RECT 4.400 30.240 496.000 31.640 ;
        RECT 3.990 24.840 496.000 30.240 ;
        RECT 3.990 23.440 495.600 24.840 ;
        RECT 3.990 21.440 496.000 23.440 ;
        RECT 4.400 20.040 496.000 21.440 ;
        RECT 3.990 14.640 496.000 20.040 ;
        RECT 3.990 13.240 495.600 14.640 ;
        RECT 3.990 11.240 496.000 13.240 ;
        RECT 4.400 9.840 496.000 11.240 ;
        RECT 3.990 4.440 496.000 9.840 ;
        RECT 3.990 3.575 495.600 4.440 ;
      LAYER met4 ;
        RECT 98.735 11.735 99.320 485.345 ;
        RECT 101.720 11.735 189.320 485.345 ;
        RECT 191.720 11.735 279.320 485.345 ;
        RECT 281.720 11.735 355.745 485.345 ;
  END
END des_Trojan
END LIBRARY

