magic
tech sky130A
magscale 1 2
timestamp 1698778774
<< obsli1 >>
rect 1104 2159 128892 127313
<< obsm1 >>
rect 14 1844 129798 127696
<< metal2 >>
rect 18 129200 74 130000
rect 1306 129200 1362 130000
rect 2594 129200 2650 130000
rect 4526 129200 4582 130000
rect 5814 129200 5870 130000
rect 7102 129200 7158 130000
rect 8390 129200 8446 130000
rect 9678 129200 9734 130000
rect 10966 129200 11022 130000
rect 12254 129200 12310 130000
rect 13542 129200 13598 130000
rect 14830 129200 14886 130000
rect 16118 129200 16174 130000
rect 17406 129200 17462 130000
rect 18694 129200 18750 130000
rect 19982 129200 20038 130000
rect 21270 129200 21326 130000
rect 22558 129200 22614 130000
rect 23846 129200 23902 130000
rect 25134 129200 25190 130000
rect 26422 129200 26478 130000
rect 27710 129200 27766 130000
rect 28998 129200 29054 130000
rect 30286 129200 30342 130000
rect 31574 129200 31630 130000
rect 32862 129200 32918 130000
rect 34150 129200 34206 130000
rect 35438 129200 35494 130000
rect 36726 129200 36782 130000
rect 38014 129200 38070 130000
rect 39302 129200 39358 130000
rect 40590 129200 40646 130000
rect 41878 129200 41934 130000
rect 43166 129200 43222 130000
rect 44454 129200 44510 130000
rect 45742 129200 45798 130000
rect 47030 129200 47086 130000
rect 48318 129200 48374 130000
rect 49606 129200 49662 130000
rect 50894 129200 50950 130000
rect 52182 129200 52238 130000
rect 53470 129200 53526 130000
rect 54758 129200 54814 130000
rect 56046 129200 56102 130000
rect 57334 129200 57390 130000
rect 58622 129200 58678 130000
rect 59910 129200 59966 130000
rect 61198 129200 61254 130000
rect 62486 129200 62542 130000
rect 63774 129200 63830 130000
rect 65062 129200 65118 130000
rect 66994 129200 67050 130000
rect 68282 129200 68338 130000
rect 69570 129200 69626 130000
rect 70858 129200 70914 130000
rect 72146 129200 72202 130000
rect 73434 129200 73490 130000
rect 74722 129200 74778 130000
rect 76010 129200 76066 130000
rect 77298 129200 77354 130000
rect 78586 129200 78642 130000
rect 79874 129200 79930 130000
rect 81162 129200 81218 130000
rect 82450 129200 82506 130000
rect 83738 129200 83794 130000
rect 85026 129200 85082 130000
rect 86314 129200 86370 130000
rect 87602 129200 87658 130000
rect 88890 129200 88946 130000
rect 90178 129200 90234 130000
rect 91466 129200 91522 130000
rect 92754 129200 92810 130000
rect 94042 129200 94098 130000
rect 95330 129200 95386 130000
rect 96618 129200 96674 130000
rect 97906 129200 97962 130000
rect 99194 129200 99250 130000
rect 100482 129200 100538 130000
rect 101770 129200 101826 130000
rect 103058 129200 103114 130000
rect 104346 129200 104402 130000
rect 105634 129200 105690 130000
rect 106922 129200 106978 130000
rect 108210 129200 108266 130000
rect 109498 129200 109554 130000
rect 110786 129200 110842 130000
rect 112074 129200 112130 130000
rect 113362 129200 113418 130000
rect 114650 129200 114706 130000
rect 115938 129200 115994 130000
rect 117226 129200 117282 130000
rect 118514 129200 118570 130000
rect 119802 129200 119858 130000
rect 121090 129200 121146 130000
rect 122378 129200 122434 130000
rect 123666 129200 123722 130000
rect 124954 129200 125010 130000
rect 126242 129200 126298 130000
rect 127530 129200 127586 130000
rect 128818 129200 128874 130000
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 32218 0 32274 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 47674 0 47730 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 51538 0 51594 800
rect 52826 0 52882 800
rect 54114 0 54170 800
rect 55402 0 55458 800
rect 56690 0 56746 800
rect 57978 0 58034 800
rect 59266 0 59322 800
rect 60554 0 60610 800
rect 61842 0 61898 800
rect 63774 0 63830 800
rect 65062 0 65118 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68926 0 68982 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 77942 0 77998 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 84382 0 84438 800
rect 85670 0 85726 800
rect 86958 0 87014 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 90822 0 90878 800
rect 92110 0 92166 800
rect 93398 0 93454 800
rect 94686 0 94742 800
rect 95974 0 96030 800
rect 97262 0 97318 800
rect 98550 0 98606 800
rect 99838 0 99894 800
rect 101126 0 101182 800
rect 102414 0 102470 800
rect 103702 0 103758 800
rect 104990 0 105046 800
rect 106278 0 106334 800
rect 107566 0 107622 800
rect 108854 0 108910 800
rect 110142 0 110198 800
rect 111430 0 111486 800
rect 112718 0 112774 800
rect 114006 0 114062 800
rect 115294 0 115350 800
rect 116582 0 116638 800
rect 117870 0 117926 800
rect 119158 0 119214 800
rect 120446 0 120502 800
rect 121734 0 121790 800
rect 123022 0 123078 800
rect 124310 0 124366 800
rect 125598 0 125654 800
rect 127530 0 127586 800
rect 128818 0 128874 800
<< obsm2 >>
rect 130 129144 1250 129282
rect 1418 129144 2538 129282
rect 2706 129144 4470 129282
rect 4638 129144 5758 129282
rect 5926 129144 7046 129282
rect 7214 129144 8334 129282
rect 8502 129144 9622 129282
rect 9790 129144 10910 129282
rect 11078 129144 12198 129282
rect 12366 129144 13486 129282
rect 13654 129144 14774 129282
rect 14942 129144 16062 129282
rect 16230 129144 17350 129282
rect 17518 129144 18638 129282
rect 18806 129144 19926 129282
rect 20094 129144 21214 129282
rect 21382 129144 22502 129282
rect 22670 129144 23790 129282
rect 23958 129144 25078 129282
rect 25246 129144 26366 129282
rect 26534 129144 27654 129282
rect 27822 129144 28942 129282
rect 29110 129144 30230 129282
rect 30398 129144 31518 129282
rect 31686 129144 32806 129282
rect 32974 129144 34094 129282
rect 34262 129144 35382 129282
rect 35550 129144 36670 129282
rect 36838 129144 37958 129282
rect 38126 129144 39246 129282
rect 39414 129144 40534 129282
rect 40702 129144 41822 129282
rect 41990 129144 43110 129282
rect 43278 129144 44398 129282
rect 44566 129144 45686 129282
rect 45854 129144 46974 129282
rect 47142 129144 48262 129282
rect 48430 129144 49550 129282
rect 49718 129144 50838 129282
rect 51006 129144 52126 129282
rect 52294 129144 53414 129282
rect 53582 129144 54702 129282
rect 54870 129144 55990 129282
rect 56158 129144 57278 129282
rect 57446 129144 58566 129282
rect 58734 129144 59854 129282
rect 60022 129144 61142 129282
rect 61310 129144 62430 129282
rect 62598 129144 63718 129282
rect 63886 129144 65006 129282
rect 65174 129144 66938 129282
rect 67106 129144 68226 129282
rect 68394 129144 69514 129282
rect 69682 129144 70802 129282
rect 70970 129144 72090 129282
rect 72258 129144 73378 129282
rect 73546 129144 74666 129282
rect 74834 129144 75954 129282
rect 76122 129144 77242 129282
rect 77410 129144 78530 129282
rect 78698 129144 79818 129282
rect 79986 129144 81106 129282
rect 81274 129144 82394 129282
rect 82562 129144 83682 129282
rect 83850 129144 84970 129282
rect 85138 129144 86258 129282
rect 86426 129144 87546 129282
rect 87714 129144 88834 129282
rect 89002 129144 90122 129282
rect 90290 129144 91410 129282
rect 91578 129144 92698 129282
rect 92866 129144 93986 129282
rect 94154 129144 95274 129282
rect 95442 129144 96562 129282
rect 96730 129144 97850 129282
rect 98018 129144 99138 129282
rect 99306 129144 100426 129282
rect 100594 129144 101714 129282
rect 101882 129144 103002 129282
rect 103170 129144 104290 129282
rect 104458 129144 105578 129282
rect 105746 129144 106866 129282
rect 107034 129144 108154 129282
rect 108322 129144 109442 129282
rect 109610 129144 110730 129282
rect 110898 129144 112018 129282
rect 112186 129144 113306 129282
rect 113474 129144 114594 129282
rect 114762 129144 115882 129282
rect 116050 129144 117170 129282
rect 117338 129144 118458 129282
rect 118626 129144 119746 129282
rect 119914 129144 121034 129282
rect 121202 129144 122322 129282
rect 122490 129144 123610 129282
rect 123778 129144 124898 129282
rect 125066 129144 126186 129282
rect 126354 129144 127474 129282
rect 127642 129144 128762 129282
rect 128930 129144 129794 129282
rect 20 856 129794 129144
rect 130 31 1250 856
rect 1418 31 2538 856
rect 2706 31 3826 856
rect 3994 31 5114 856
rect 5282 31 6402 856
rect 6570 31 7690 856
rect 7858 31 8978 856
rect 9146 31 10266 856
rect 10434 31 11554 856
rect 11722 31 12842 856
rect 13010 31 14130 856
rect 14298 31 15418 856
rect 15586 31 16706 856
rect 16874 31 17994 856
rect 18162 31 19282 856
rect 19450 31 20570 856
rect 20738 31 21858 856
rect 22026 31 23146 856
rect 23314 31 24434 856
rect 24602 31 25722 856
rect 25890 31 27010 856
rect 27178 31 28298 856
rect 28466 31 29586 856
rect 29754 31 30874 856
rect 31042 31 32162 856
rect 32330 31 33450 856
rect 33618 31 34738 856
rect 34906 31 36026 856
rect 36194 31 37314 856
rect 37482 31 38602 856
rect 38770 31 39890 856
rect 40058 31 41178 856
rect 41346 31 42466 856
rect 42634 31 43754 856
rect 43922 31 45042 856
rect 45210 31 46330 856
rect 46498 31 47618 856
rect 47786 31 48906 856
rect 49074 31 50194 856
rect 50362 31 51482 856
rect 51650 31 52770 856
rect 52938 31 54058 856
rect 54226 31 55346 856
rect 55514 31 56634 856
rect 56802 31 57922 856
rect 58090 31 59210 856
rect 59378 31 60498 856
rect 60666 31 61786 856
rect 61954 31 63718 856
rect 63886 31 65006 856
rect 65174 31 66294 856
rect 66462 31 67582 856
rect 67750 31 68870 856
rect 69038 31 70158 856
rect 70326 31 71446 856
rect 71614 31 72734 856
rect 72902 31 74022 856
rect 74190 31 75310 856
rect 75478 31 76598 856
rect 76766 31 77886 856
rect 78054 31 79174 856
rect 79342 31 80462 856
rect 80630 31 81750 856
rect 81918 31 83038 856
rect 83206 31 84326 856
rect 84494 31 85614 856
rect 85782 31 86902 856
rect 87070 31 88190 856
rect 88358 31 89478 856
rect 89646 31 90766 856
rect 90934 31 92054 856
rect 92222 31 93342 856
rect 93510 31 94630 856
rect 94798 31 95918 856
rect 96086 31 97206 856
rect 97374 31 98494 856
rect 98662 31 99782 856
rect 99950 31 101070 856
rect 101238 31 102358 856
rect 102526 31 103646 856
rect 103814 31 104934 856
rect 105102 31 106222 856
rect 106390 31 107510 856
rect 107678 31 108798 856
rect 108966 31 110086 856
rect 110254 31 111374 856
rect 111542 31 112662 856
rect 112830 31 113950 856
rect 114118 31 115238 856
rect 115406 31 116526 856
rect 116694 31 117814 856
rect 117982 31 119102 856
rect 119270 31 120390 856
rect 120558 31 121678 856
rect 121846 31 122966 856
rect 123134 31 124254 856
rect 124422 31 125542 856
rect 125710 31 127474 856
rect 127642 31 128762 856
rect 128930 31 129794 856
<< metal3 >>
rect 0 128528 800 128648
rect 129200 128528 130000 128648
rect 0 127168 800 127288
rect 129200 127168 130000 127288
rect 0 125808 800 125928
rect 129200 125808 130000 125928
rect 0 124448 800 124568
rect 129200 124448 130000 124568
rect 0 123088 800 123208
rect 129200 123088 130000 123208
rect 0 121728 800 121848
rect 129200 121728 130000 121848
rect 0 120368 800 120488
rect 129200 120368 130000 120488
rect 0 119008 800 119128
rect 129200 119008 130000 119128
rect 0 117648 800 117768
rect 129200 117648 130000 117768
rect 0 116288 800 116408
rect 129200 116288 130000 116408
rect 0 114928 800 115048
rect 129200 114928 130000 115048
rect 0 113568 800 113688
rect 129200 113568 130000 113688
rect 0 112208 800 112328
rect 129200 112208 130000 112328
rect 0 110848 800 110968
rect 129200 110848 130000 110968
rect 0 109488 800 109608
rect 129200 109488 130000 109608
rect 0 108128 800 108248
rect 129200 108128 130000 108248
rect 0 106768 800 106888
rect 129200 106768 130000 106888
rect 0 105408 800 105528
rect 129200 105408 130000 105528
rect 0 104048 800 104168
rect 129200 104048 130000 104168
rect 0 102688 800 102808
rect 129200 102688 130000 102808
rect 0 101328 800 101448
rect 129200 101328 130000 101448
rect 0 99968 800 100088
rect 129200 99968 130000 100088
rect 0 98608 800 98728
rect 129200 98608 130000 98728
rect 0 97248 800 97368
rect 129200 97248 130000 97368
rect 0 95888 800 96008
rect 129200 95888 130000 96008
rect 0 94528 800 94648
rect 129200 94528 130000 94648
rect 0 93168 800 93288
rect 129200 93168 130000 93288
rect 0 91808 800 91928
rect 129200 91808 130000 91928
rect 0 90448 800 90568
rect 129200 90448 130000 90568
rect 0 89088 800 89208
rect 129200 89088 130000 89208
rect 0 87728 800 87848
rect 129200 87728 130000 87848
rect 0 86368 800 86488
rect 129200 86368 130000 86488
rect 0 85008 800 85128
rect 129200 85008 130000 85128
rect 0 83648 800 83768
rect 129200 83648 130000 83768
rect 0 82288 800 82408
rect 129200 82288 130000 82408
rect 0 80928 800 81048
rect 129200 80928 130000 81048
rect 0 79568 800 79688
rect 129200 79568 130000 79688
rect 0 78208 800 78328
rect 129200 78208 130000 78328
rect 0 76848 800 76968
rect 129200 76848 130000 76968
rect 0 75488 800 75608
rect 129200 75488 130000 75608
rect 0 74128 800 74248
rect 129200 74128 130000 74248
rect 0 72768 800 72888
rect 129200 72768 130000 72888
rect 0 71408 800 71528
rect 129200 71408 130000 71528
rect 0 70048 800 70168
rect 129200 70048 130000 70168
rect 0 68688 800 68808
rect 129200 68688 130000 68808
rect 0 67328 800 67448
rect 129200 67328 130000 67448
rect 129200 65968 130000 66088
rect 0 65288 800 65408
rect 129200 64608 130000 64728
rect 0 63928 800 64048
rect 129200 63248 130000 63368
rect 0 62568 800 62688
rect 0 61208 800 61328
rect 129200 61208 130000 61328
rect 0 59848 800 59968
rect 129200 59848 130000 59968
rect 0 58488 800 58608
rect 129200 58488 130000 58608
rect 0 57128 800 57248
rect 129200 57128 130000 57248
rect 0 55768 800 55888
rect 129200 55768 130000 55888
rect 0 54408 800 54528
rect 129200 54408 130000 54528
rect 0 53048 800 53168
rect 129200 53048 130000 53168
rect 0 51688 800 51808
rect 129200 51688 130000 51808
rect 0 50328 800 50448
rect 129200 50328 130000 50448
rect 0 48968 800 49088
rect 129200 48968 130000 49088
rect 0 47608 800 47728
rect 129200 47608 130000 47728
rect 0 46248 800 46368
rect 129200 46248 130000 46368
rect 0 44888 800 45008
rect 129200 44888 130000 45008
rect 0 43528 800 43648
rect 129200 43528 130000 43648
rect 0 42168 800 42288
rect 129200 42168 130000 42288
rect 0 40808 800 40928
rect 129200 40808 130000 40928
rect 0 39448 800 39568
rect 129200 39448 130000 39568
rect 0 38088 800 38208
rect 129200 38088 130000 38208
rect 0 36728 800 36848
rect 129200 36728 130000 36848
rect 0 35368 800 35488
rect 129200 35368 130000 35488
rect 0 34008 800 34128
rect 129200 34008 130000 34128
rect 0 32648 800 32768
rect 129200 32648 130000 32768
rect 0 31288 800 31408
rect 129200 31288 130000 31408
rect 0 29928 800 30048
rect 129200 29928 130000 30048
rect 0 28568 800 28688
rect 129200 28568 130000 28688
rect 0 27208 800 27328
rect 129200 27208 130000 27328
rect 0 25848 800 25968
rect 129200 25848 130000 25968
rect 0 24488 800 24608
rect 129200 24488 130000 24608
rect 0 23128 800 23248
rect 129200 23128 130000 23248
rect 0 21768 800 21888
rect 129200 21768 130000 21888
rect 0 20408 800 20528
rect 129200 20408 130000 20528
rect 0 19048 800 19168
rect 129200 19048 130000 19168
rect 0 17688 800 17808
rect 129200 17688 130000 17808
rect 0 16328 800 16448
rect 129200 16328 130000 16448
rect 0 14968 800 15088
rect 129200 14968 130000 15088
rect 0 13608 800 13728
rect 129200 13608 130000 13728
rect 0 12248 800 12368
rect 129200 12248 130000 12368
rect 0 10888 800 11008
rect 129200 10888 130000 11008
rect 0 9528 800 9648
rect 129200 9528 130000 9648
rect 0 8168 800 8288
rect 129200 8168 130000 8288
rect 0 6808 800 6928
rect 129200 6808 130000 6928
rect 0 5448 800 5568
rect 129200 5448 130000 5568
rect 0 4088 800 4208
rect 129200 4088 130000 4208
rect 0 2728 800 2848
rect 129200 2728 130000 2848
rect 0 1368 800 1488
rect 129200 1368 130000 1488
rect 129200 8 130000 128
<< obsm3 >>
rect 880 128448 129120 128621
rect 798 127368 129799 128448
rect 880 127088 129120 127368
rect 798 126008 129799 127088
rect 880 125728 129120 126008
rect 798 124648 129799 125728
rect 880 124368 129120 124648
rect 798 123288 129799 124368
rect 880 123008 129120 123288
rect 798 121928 129799 123008
rect 880 121648 129120 121928
rect 798 120568 129799 121648
rect 880 120288 129120 120568
rect 798 119208 129799 120288
rect 880 118928 129120 119208
rect 798 117848 129799 118928
rect 880 117568 129120 117848
rect 798 116488 129799 117568
rect 880 116208 129120 116488
rect 798 115128 129799 116208
rect 880 114848 129120 115128
rect 798 113768 129799 114848
rect 880 113488 129120 113768
rect 798 112408 129799 113488
rect 880 112128 129120 112408
rect 798 111048 129799 112128
rect 880 110768 129120 111048
rect 798 109688 129799 110768
rect 880 109408 129120 109688
rect 798 108328 129799 109408
rect 880 108048 129120 108328
rect 798 106968 129799 108048
rect 880 106688 129120 106968
rect 798 105608 129799 106688
rect 880 105328 129120 105608
rect 798 104248 129799 105328
rect 880 103968 129120 104248
rect 798 102888 129799 103968
rect 880 102608 129120 102888
rect 798 101528 129799 102608
rect 880 101248 129120 101528
rect 798 100168 129799 101248
rect 880 99888 129120 100168
rect 798 98808 129799 99888
rect 880 98528 129120 98808
rect 798 97448 129799 98528
rect 880 97168 129120 97448
rect 798 96088 129799 97168
rect 880 95808 129120 96088
rect 798 94728 129799 95808
rect 880 94448 129120 94728
rect 798 93368 129799 94448
rect 880 93088 129120 93368
rect 798 92008 129799 93088
rect 880 91728 129120 92008
rect 798 90648 129799 91728
rect 880 90368 129120 90648
rect 798 89288 129799 90368
rect 880 89008 129120 89288
rect 798 87928 129799 89008
rect 880 87648 129120 87928
rect 798 86568 129799 87648
rect 880 86288 129120 86568
rect 798 85208 129799 86288
rect 880 84928 129120 85208
rect 798 83848 129799 84928
rect 880 83568 129120 83848
rect 798 82488 129799 83568
rect 880 82208 129120 82488
rect 798 81128 129799 82208
rect 880 80848 129120 81128
rect 798 79768 129799 80848
rect 880 79488 129120 79768
rect 798 78408 129799 79488
rect 880 78128 129120 78408
rect 798 77048 129799 78128
rect 880 76768 129120 77048
rect 798 75688 129799 76768
rect 880 75408 129120 75688
rect 798 74328 129799 75408
rect 880 74048 129120 74328
rect 798 72968 129799 74048
rect 880 72688 129120 72968
rect 798 71608 129799 72688
rect 880 71328 129120 71608
rect 798 70248 129799 71328
rect 880 69968 129120 70248
rect 798 68888 129799 69968
rect 880 68608 129120 68888
rect 798 67528 129799 68608
rect 880 67248 129120 67528
rect 798 66168 129799 67248
rect 798 65888 129120 66168
rect 798 65488 129799 65888
rect 880 65208 129799 65488
rect 798 64808 129799 65208
rect 798 64528 129120 64808
rect 798 64128 129799 64528
rect 880 63848 129799 64128
rect 798 63448 129799 63848
rect 798 63168 129120 63448
rect 798 62768 129799 63168
rect 880 62488 129799 62768
rect 798 61408 129799 62488
rect 880 61128 129120 61408
rect 798 60048 129799 61128
rect 880 59768 129120 60048
rect 798 58688 129799 59768
rect 880 58408 129120 58688
rect 798 57328 129799 58408
rect 880 57048 129120 57328
rect 798 55968 129799 57048
rect 880 55688 129120 55968
rect 798 54608 129799 55688
rect 880 54328 129120 54608
rect 798 53248 129799 54328
rect 880 52968 129120 53248
rect 798 51888 129799 52968
rect 880 51608 129120 51888
rect 798 50528 129799 51608
rect 880 50248 129120 50528
rect 798 49168 129799 50248
rect 880 48888 129120 49168
rect 798 47808 129799 48888
rect 880 47528 129120 47808
rect 798 46448 129799 47528
rect 880 46168 129120 46448
rect 798 45088 129799 46168
rect 880 44808 129120 45088
rect 798 43728 129799 44808
rect 880 43448 129120 43728
rect 798 42368 129799 43448
rect 880 42088 129120 42368
rect 798 41008 129799 42088
rect 880 40728 129120 41008
rect 798 39648 129799 40728
rect 880 39368 129120 39648
rect 798 38288 129799 39368
rect 880 38008 129120 38288
rect 798 36928 129799 38008
rect 880 36648 129120 36928
rect 798 35568 129799 36648
rect 880 35288 129120 35568
rect 798 34208 129799 35288
rect 880 33928 129120 34208
rect 798 32848 129799 33928
rect 880 32568 129120 32848
rect 798 31488 129799 32568
rect 880 31208 129120 31488
rect 798 30128 129799 31208
rect 880 29848 129120 30128
rect 798 28768 129799 29848
rect 880 28488 129120 28768
rect 798 27408 129799 28488
rect 880 27128 129120 27408
rect 798 26048 129799 27128
rect 880 25768 129120 26048
rect 798 24688 129799 25768
rect 880 24408 129120 24688
rect 798 23328 129799 24408
rect 880 23048 129120 23328
rect 798 21968 129799 23048
rect 880 21688 129120 21968
rect 798 20608 129799 21688
rect 880 20328 129120 20608
rect 798 19248 129799 20328
rect 880 18968 129120 19248
rect 798 17888 129799 18968
rect 880 17608 129120 17888
rect 798 16528 129799 17608
rect 880 16248 129120 16528
rect 798 15168 129799 16248
rect 880 14888 129120 15168
rect 798 13808 129799 14888
rect 880 13528 129120 13808
rect 798 12448 129799 13528
rect 880 12168 129120 12448
rect 798 11088 129799 12168
rect 880 10808 129120 11088
rect 798 9728 129799 10808
rect 880 9448 129120 9728
rect 798 8368 129799 9448
rect 880 8088 129120 8368
rect 798 7008 129799 8088
rect 880 6728 129120 7008
rect 798 5648 129799 6728
rect 880 5368 129120 5648
rect 798 4288 129799 5368
rect 880 4008 129120 4288
rect 798 2928 129799 4008
rect 880 2648 129120 2928
rect 798 1568 129799 2648
rect 880 1288 129120 1568
rect 798 208 129799 1288
rect 798 35 129120 208
<< metal4 >>
rect 1944 2128 2264 127344
rect 19944 2128 20264 127344
rect 37944 2128 38264 127344
rect 55944 2128 56264 127344
rect 73944 2128 74264 127344
rect 91944 2128 92264 127344
rect 109944 2128 110264 127344
rect 127944 2128 128264 127344
<< obsm4 >>
rect 23979 127424 117885 127805
rect 23979 2048 37864 127424
rect 38344 2048 55864 127424
rect 56344 2048 73864 127424
rect 74344 2048 91864 127424
rect 92344 2048 109864 127424
rect 110344 2048 117885 127424
rect 23979 1531 117885 2048
<< labels >>
rlabel metal3 s 0 99968 800 100088 6 clk
port 1 nsew signal input
rlabel metal2 s 12254 129200 12310 130000 6 data_i[0]
port 2 nsew signal input
rlabel metal2 s 65062 129200 65118 130000 6 data_i[100]
port 3 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 data_i[101]
port 4 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 data_i[102]
port 5 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 data_i[103]
port 6 nsew signal input
rlabel metal3 s 129200 39448 130000 39568 6 data_i[104]
port 7 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 data_i[105]
port 8 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 data_i[106]
port 9 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 data_i[107]
port 10 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 data_i[108]
port 11 nsew signal input
rlabel metal3 s 129200 67328 130000 67448 6 data_i[109]
port 12 nsew signal input
rlabel metal3 s 129200 102688 130000 102808 6 data_i[10]
port 13 nsew signal input
rlabel metal3 s 129200 14968 130000 15088 6 data_i[110]
port 14 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 data_i[111]
port 15 nsew signal input
rlabel metal2 s 4526 129200 4582 130000 6 data_i[112]
port 16 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 data_i[113]
port 17 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 data_i[114]
port 18 nsew signal input
rlabel metal2 s 112074 129200 112130 130000 6 data_i[115]
port 19 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 data_i[116]
port 20 nsew signal input
rlabel metal3 s 129200 68688 130000 68808 6 data_i[117]
port 21 nsew signal input
rlabel metal2 s 2594 129200 2650 130000 6 data_i[118]
port 22 nsew signal input
rlabel metal2 s 58622 129200 58678 130000 6 data_i[119]
port 23 nsew signal input
rlabel metal3 s 129200 124448 130000 124568 6 data_i[11]
port 24 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 data_i[120]
port 25 nsew signal input
rlabel metal2 s 82450 129200 82506 130000 6 data_i[121]
port 26 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 data_i[122]
port 27 nsew signal input
rlabel metal3 s 129200 28568 130000 28688 6 data_i[123]
port 28 nsew signal input
rlabel metal2 s 77298 129200 77354 130000 6 data_i[124]
port 29 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 data_i[125]
port 30 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 data_i[126]
port 31 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 data_i[127]
port 32 nsew signal input
rlabel metal2 s 1306 129200 1362 130000 6 data_i[12]
port 33 nsew signal input
rlabel metal2 s 99194 129200 99250 130000 6 data_i[13]
port 34 nsew signal input
rlabel metal2 s 72146 129200 72202 130000 6 data_i[14]
port 35 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 data_i[15]
port 36 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 data_i[16]
port 37 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 data_i[17]
port 38 nsew signal input
rlabel metal2 s 50894 129200 50950 130000 6 data_i[18]
port 39 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 data_i[19]
port 40 nsew signal input
rlabel metal2 s 57334 129200 57390 130000 6 data_i[1]
port 41 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 data_i[20]
port 42 nsew signal input
rlabel metal2 s 7102 129200 7158 130000 6 data_i[21]
port 43 nsew signal input
rlabel metal3 s 129200 99968 130000 100088 6 data_i[22]
port 44 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 data_i[23]
port 45 nsew signal input
rlabel metal2 s 47030 129200 47086 130000 6 data_i[24]
port 46 nsew signal input
rlabel metal2 s 115938 129200 115994 130000 6 data_i[25]
port 47 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 data_i[26]
port 48 nsew signal input
rlabel metal2 s 103058 129200 103114 130000 6 data_i[27]
port 49 nsew signal input
rlabel metal3 s 129200 80928 130000 81048 6 data_i[28]
port 50 nsew signal input
rlabel metal3 s 129200 86368 130000 86488 6 data_i[29]
port 51 nsew signal input
rlabel metal3 s 129200 116288 130000 116408 6 data_i[2]
port 52 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 data_i[30]
port 53 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 data_i[31]
port 54 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 data_i[32]
port 55 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 data_i[33]
port 56 nsew signal input
rlabel metal2 s 19982 129200 20038 130000 6 data_i[34]
port 57 nsew signal input
rlabel metal2 s 32862 129200 32918 130000 6 data_i[35]
port 58 nsew signal input
rlabel metal2 s 62486 129200 62542 130000 6 data_i[36]
port 59 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 data_i[37]
port 60 nsew signal input
rlabel metal2 s 106922 129200 106978 130000 6 data_i[38]
port 61 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 data_i[39]
port 62 nsew signal input
rlabel metal3 s 129200 31288 130000 31408 6 data_i[3]
port 63 nsew signal input
rlabel metal2 s 96618 129200 96674 130000 6 data_i[40]
port 64 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 data_i[41]
port 65 nsew signal input
rlabel metal3 s 129200 20408 130000 20528 6 data_i[42]
port 66 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 data_i[43]
port 67 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 data_i[44]
port 68 nsew signal input
rlabel metal2 s 128818 129200 128874 130000 6 data_i[45]
port 69 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 data_i[46]
port 70 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 data_i[47]
port 71 nsew signal input
rlabel metal2 s 45742 129200 45798 130000 6 data_i[48]
port 72 nsew signal input
rlabel metal2 s 78586 129200 78642 130000 6 data_i[49]
port 73 nsew signal input
rlabel metal3 s 129200 12248 130000 12368 6 data_i[4]
port 74 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 data_i[50]
port 75 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 data_i[51]
port 76 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 data_i[52]
port 77 nsew signal input
rlabel metal2 s 113362 129200 113418 130000 6 data_i[53]
port 78 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 data_i[54]
port 79 nsew signal input
rlabel metal3 s 129200 128528 130000 128648 6 data_i[55]
port 80 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 data_i[56]
port 81 nsew signal input
rlabel metal2 s 49606 129200 49662 130000 6 data_i[57]
port 82 nsew signal input
rlabel metal3 s 129200 44888 130000 45008 6 data_i[58]
port 83 nsew signal input
rlabel metal3 s 129200 106768 130000 106888 6 data_i[59]
port 84 nsew signal input
rlabel metal2 s 28998 129200 29054 130000 6 data_i[5]
port 85 nsew signal input
rlabel metal3 s 129200 114928 130000 115048 6 data_i[60]
port 86 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 data_i[61]
port 87 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 data_i[62]
port 88 nsew signal input
rlabel metal3 s 129200 65968 130000 66088 6 data_i[63]
port 89 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 data_i[64]
port 90 nsew signal input
rlabel metal3 s 129200 23128 130000 23248 6 data_i[65]
port 91 nsew signal input
rlabel metal2 s 9678 129200 9734 130000 6 data_i[66]
port 92 nsew signal input
rlabel metal2 s 59910 129200 59966 130000 6 data_i[67]
port 93 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 data_i[68]
port 94 nsew signal input
rlabel metal3 s 129200 47608 130000 47728 6 data_i[69]
port 95 nsew signal input
rlabel metal2 s 76010 129200 76066 130000 6 data_i[6]
port 96 nsew signal input
rlabel metal2 s 79874 129200 79930 130000 6 data_i[70]
port 97 nsew signal input
rlabel metal3 s 129200 8168 130000 8288 6 data_i[71]
port 98 nsew signal input
rlabel metal2 s 66994 129200 67050 130000 6 data_i[72]
port 99 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 data_i[73]
port 100 nsew signal input
rlabel metal3 s 129200 76848 130000 76968 6 data_i[74]
port 101 nsew signal input
rlabel metal2 s 27710 129200 27766 130000 6 data_i[75]
port 102 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 data_i[76]
port 103 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 data_i[77]
port 104 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 data_i[78]
port 105 nsew signal input
rlabel metal2 s 44454 129200 44510 130000 6 data_i[79]
port 106 nsew signal input
rlabel metal3 s 129200 13608 130000 13728 6 data_i[7]
port 107 nsew signal input
rlabel metal3 s 129200 90448 130000 90568 6 data_i[80]
port 108 nsew signal input
rlabel metal2 s 34150 129200 34206 130000 6 data_i[81]
port 109 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 data_i[82]
port 110 nsew signal input
rlabel metal3 s 129200 105408 130000 105528 6 data_i[83]
port 111 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 data_i[84]
port 112 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 data_i[85]
port 113 nsew signal input
rlabel metal3 s 129200 59848 130000 59968 6 data_i[86]
port 114 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 data_i[87]
port 115 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 data_i[88]
port 116 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 data_i[89]
port 117 nsew signal input
rlabel metal3 s 129200 108128 130000 108248 6 data_i[8]
port 118 nsew signal input
rlabel metal2 s 88890 129200 88946 130000 6 data_i[90]
port 119 nsew signal input
rlabel metal3 s 129200 123088 130000 123208 6 data_i[91]
port 120 nsew signal input
rlabel metal3 s 129200 19048 130000 19168 6 data_i[92]
port 121 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 data_i[93]
port 122 nsew signal input
rlabel metal2 s 16118 129200 16174 130000 6 data_i[94]
port 123 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 data_i[95]
port 124 nsew signal input
rlabel metal2 s 10966 129200 11022 130000 6 data_i[96]
port 125 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 data_i[97]
port 126 nsew signal input
rlabel metal2 s 13542 129200 13598 130000 6 data_i[98]
port 127 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 data_i[99]
port 128 nsew signal input
rlabel metal2 s 26422 129200 26478 130000 6 data_i[9]
port 129 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 data_o[0]
port 130 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 data_o[100]
port 131 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 data_o[101]
port 132 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 data_o[102]
port 133 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 data_o[103]
port 134 nsew signal output
rlabel metal3 s 129200 91808 130000 91928 6 data_o[104]
port 135 nsew signal output
rlabel metal3 s 129200 83648 130000 83768 6 data_o[105]
port 136 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 data_o[106]
port 137 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 data_o[107]
port 138 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 data_o[108]
port 139 nsew signal output
rlabel metal2 s 22558 129200 22614 130000 6 data_o[109]
port 140 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 data_o[10]
port 141 nsew signal output
rlabel metal3 s 129200 121728 130000 121848 6 data_o[110]
port 142 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 data_o[111]
port 143 nsew signal output
rlabel metal3 s 129200 40808 130000 40928 6 data_o[112]
port 144 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 data_o[113]
port 145 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 data_o[114]
port 146 nsew signal output
rlabel metal3 s 129200 97248 130000 97368 6 data_o[115]
port 147 nsew signal output
rlabel metal2 s 30286 129200 30342 130000 6 data_o[116]
port 148 nsew signal output
rlabel metal3 s 129200 27208 130000 27328 6 data_o[117]
port 149 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 data_o[118]
port 150 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 data_o[119]
port 151 nsew signal output
rlabel metal3 s 129200 46248 130000 46368 6 data_o[11]
port 152 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 data_o[120]
port 153 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 data_o[121]
port 154 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 data_o[122]
port 155 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 data_o[123]
port 156 nsew signal output
rlabel metal3 s 129200 110848 130000 110968 6 data_o[124]
port 157 nsew signal output
rlabel metal3 s 129200 104048 130000 104168 6 data_o[125]
port 158 nsew signal output
rlabel metal3 s 129200 51688 130000 51808 6 data_o[126]
port 159 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 data_o[127]
port 160 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 data_o[12]
port 161 nsew signal output
rlabel metal2 s 121090 129200 121146 130000 6 data_o[13]
port 162 nsew signal output
rlabel metal3 s 129200 42168 130000 42288 6 data_o[14]
port 163 nsew signal output
rlabel metal2 s 127530 129200 127586 130000 6 data_o[15]
port 164 nsew signal output
rlabel metal2 s 18 129200 74 130000 6 data_o[16]
port 165 nsew signal output
rlabel metal3 s 0 87728 800 87848 6 data_o[17]
port 166 nsew signal output
rlabel metal2 s 83738 129200 83794 130000 6 data_o[18]
port 167 nsew signal output
rlabel metal3 s 129200 21768 130000 21888 6 data_o[19]
port 168 nsew signal output
rlabel metal2 s 69570 129200 69626 130000 6 data_o[1]
port 169 nsew signal output
rlabel metal3 s 0 125808 800 125928 6 data_o[20]
port 170 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 data_o[21]
port 171 nsew signal output
rlabel metal3 s 129200 85008 130000 85128 6 data_o[22]
port 172 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 data_o[23]
port 173 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 data_o[24]
port 174 nsew signal output
rlabel metal3 s 129200 43528 130000 43648 6 data_o[25]
port 175 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 data_o[26]
port 176 nsew signal output
rlabel metal2 s 63774 129200 63830 130000 6 data_o[27]
port 177 nsew signal output
rlabel metal3 s 129200 9528 130000 9648 6 data_o[28]
port 178 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 data_o[29]
port 179 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 data_o[2]
port 180 nsew signal output
rlabel metal3 s 129200 87728 130000 87848 6 data_o[30]
port 181 nsew signal output
rlabel metal3 s 129200 35368 130000 35488 6 data_o[31]
port 182 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 data_o[32]
port 183 nsew signal output
rlabel metal3 s 129200 4088 130000 4208 6 data_o[33]
port 184 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 data_o[34]
port 185 nsew signal output
rlabel metal2 s 31574 129200 31630 130000 6 data_o[35]
port 186 nsew signal output
rlabel metal3 s 129200 25848 130000 25968 6 data_o[36]
port 187 nsew signal output
rlabel metal2 s 8390 129200 8446 130000 6 data_o[37]
port 188 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 data_o[38]
port 189 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 data_o[39]
port 190 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 data_o[3]
port 191 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 data_o[40]
port 192 nsew signal output
rlabel metal3 s 0 90448 800 90568 6 data_o[41]
port 193 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 data_o[42]
port 194 nsew signal output
rlabel metal2 s 81162 129200 81218 130000 6 data_o[43]
port 195 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 data_o[44]
port 196 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 data_o[45]
port 197 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 data_o[46]
port 198 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 data_o[47]
port 199 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 data_o[48]
port 200 nsew signal output
rlabel metal2 s 40590 129200 40646 130000 6 data_o[49]
port 201 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 data_o[4]
port 202 nsew signal output
rlabel metal3 s 129200 17688 130000 17808 6 data_o[50]
port 203 nsew signal output
rlabel metal2 s 114650 129200 114706 130000 6 data_o[51]
port 204 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 data_o[52]
port 205 nsew signal output
rlabel metal2 s 73434 129200 73490 130000 6 data_o[53]
port 206 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 data_o[54]
port 207 nsew signal output
rlabel metal2 s 119802 129200 119858 130000 6 data_o[55]
port 208 nsew signal output
rlabel metal2 s 23846 129200 23902 130000 6 data_o[56]
port 209 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 data_o[57]
port 210 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 data_o[58]
port 211 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 data_o[59]
port 212 nsew signal output
rlabel metal2 s 74722 129200 74778 130000 6 data_o[5]
port 213 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 data_o[60]
port 214 nsew signal output
rlabel metal3 s 129200 50328 130000 50448 6 data_o[61]
port 215 nsew signal output
rlabel metal3 s 129200 36728 130000 36848 6 data_o[62]
port 216 nsew signal output
rlabel metal3 s 129200 79568 130000 79688 6 data_o[63]
port 217 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 data_o[64]
port 218 nsew signal output
rlabel metal2 s 21270 129200 21326 130000 6 data_o[65]
port 219 nsew signal output
rlabel metal3 s 129200 64608 130000 64728 6 data_o[66]
port 220 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 data_o[67]
port 221 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 data_o[68]
port 222 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 data_o[69]
port 223 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 data_o[6]
port 224 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 data_o[70]
port 225 nsew signal output
rlabel metal3 s 129200 1368 130000 1488 6 data_o[71]
port 226 nsew signal output
rlabel metal3 s 129200 55768 130000 55888 6 data_o[72]
port 227 nsew signal output
rlabel metal3 s 129200 127168 130000 127288 6 data_o[73]
port 228 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 data_o[74]
port 229 nsew signal output
rlabel metal2 s 109498 129200 109554 130000 6 data_o[75]
port 230 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 data_o[76]
port 231 nsew signal output
rlabel metal3 s 129200 70048 130000 70168 6 data_o[77]
port 232 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 data_o[78]
port 233 nsew signal output
rlabel metal2 s 101770 129200 101826 130000 6 data_o[79]
port 234 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 data_o[7]
port 235 nsew signal output
rlabel metal2 s 38014 129200 38070 130000 6 data_o[80]
port 236 nsew signal output
rlabel metal3 s 129200 112208 130000 112328 6 data_o[81]
port 237 nsew signal output
rlabel metal3 s 129200 120368 130000 120488 6 data_o[82]
port 238 nsew signal output
rlabel metal3 s 129200 101328 130000 101448 6 data_o[83]
port 239 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 data_o[84]
port 240 nsew signal output
rlabel metal3 s 129200 95888 130000 96008 6 data_o[85]
port 241 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 data_o[86]
port 242 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 data_o[87]
port 243 nsew signal output
rlabel metal2 s 56046 129200 56102 130000 6 data_o[88]
port 244 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 data_o[89]
port 245 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 data_o[8]
port 246 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 data_o[90]
port 247 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 data_o[91]
port 248 nsew signal output
rlabel metal3 s 129200 125808 130000 125928 6 data_o[92]
port 249 nsew signal output
rlabel metal3 s 129200 6808 130000 6928 6 data_o[93]
port 250 nsew signal output
rlabel metal2 s 61198 129200 61254 130000 6 data_o[94]
port 251 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 data_o[95]
port 252 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 data_o[96]
port 253 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 data_o[97]
port 254 nsew signal output
rlabel metal2 s 117226 129200 117282 130000 6 data_o[98]
port 255 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 data_o[99]
port 256 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 data_o[9]
port 257 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 decrypt_i
port 258 nsew signal input
rlabel metal3 s 129200 54408 130000 54528 6 key_i[0]
port 259 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 key_i[100]
port 260 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 key_i[101]
port 261 nsew signal input
rlabel metal2 s 54758 129200 54814 130000 6 key_i[102]
port 262 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 key_i[103]
port 263 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 key_i[104]
port 264 nsew signal input
rlabel metal2 s 97906 129200 97962 130000 6 key_i[105]
port 265 nsew signal input
rlabel metal3 s 129200 58488 130000 58608 6 key_i[106]
port 266 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 key_i[107]
port 267 nsew signal input
rlabel metal2 s 122378 129200 122434 130000 6 key_i[108]
port 268 nsew signal input
rlabel metal3 s 129200 5448 130000 5568 6 key_i[109]
port 269 nsew signal input
rlabel metal2 s 86314 129200 86370 130000 6 key_i[10]
port 270 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 key_i[110]
port 271 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 key_i[111]
port 272 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 key_i[112]
port 273 nsew signal input
rlabel metal3 s 129200 57128 130000 57248 6 key_i[113]
port 274 nsew signal input
rlabel metal2 s 5814 129200 5870 130000 6 key_i[114]
port 275 nsew signal input
rlabel metal3 s 129200 78208 130000 78328 6 key_i[115]
port 276 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 key_i[116]
port 277 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 key_i[117]
port 278 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 key_i[118]
port 279 nsew signal input
rlabel metal2 s 118514 129200 118570 130000 6 key_i[119]
port 280 nsew signal input
rlabel metal3 s 129200 93168 130000 93288 6 key_i[11]
port 281 nsew signal input
rlabel metal2 s 43166 129200 43222 130000 6 key_i[120]
port 282 nsew signal input
rlabel metal2 s 53470 129200 53526 130000 6 key_i[121]
port 283 nsew signal input
rlabel metal3 s 129200 16328 130000 16448 6 key_i[122]
port 284 nsew signal input
rlabel metal2 s 35438 129200 35494 130000 6 key_i[123]
port 285 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 key_i[124]
port 286 nsew signal input
rlabel metal2 s 94042 129200 94098 130000 6 key_i[125]
port 287 nsew signal input
rlabel metal2 s 68282 129200 68338 130000 6 key_i[126]
port 288 nsew signal input
rlabel metal2 s 18694 129200 18750 130000 6 key_i[127]
port 289 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 key_i[12]
port 290 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 key_i[13]
port 291 nsew signal input
rlabel metal3 s 129200 89088 130000 89208 6 key_i[14]
port 292 nsew signal input
rlabel metal3 s 129200 82288 130000 82408 6 key_i[15]
port 293 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 key_i[16]
port 294 nsew signal input
rlabel metal3 s 129200 72768 130000 72888 6 key_i[17]
port 295 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 key_i[18]
port 296 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 key_i[19]
port 297 nsew signal input
rlabel metal2 s 90178 129200 90234 130000 6 key_i[1]
port 298 nsew signal input
rlabel metal2 s 124954 129200 125010 130000 6 key_i[20]
port 299 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 key_i[21]
port 300 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 key_i[22]
port 301 nsew signal input
rlabel metal3 s 129200 24488 130000 24608 6 key_i[23]
port 302 nsew signal input
rlabel metal2 s 25134 129200 25190 130000 6 key_i[24]
port 303 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 key_i[25]
port 304 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 key_i[26]
port 305 nsew signal input
rlabel metal2 s 52182 129200 52238 130000 6 key_i[27]
port 306 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 key_i[28]
port 307 nsew signal input
rlabel metal3 s 129200 119008 130000 119128 6 key_i[29]
port 308 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 key_i[2]
port 309 nsew signal input
rlabel metal2 s 108210 129200 108266 130000 6 key_i[30]
port 310 nsew signal input
rlabel metal3 s 129200 48968 130000 49088 6 key_i[31]
port 311 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 key_i[32]
port 312 nsew signal input
rlabel metal2 s 104346 129200 104402 130000 6 key_i[33]
port 313 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 key_i[34]
port 314 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 key_i[35]
port 315 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 key_i[36]
port 316 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 key_i[37]
port 317 nsew signal input
rlabel metal3 s 129200 29928 130000 30048 6 key_i[38]
port 318 nsew signal input
rlabel metal2 s 48318 129200 48374 130000 6 key_i[39]
port 319 nsew signal input
rlabel metal3 s 129200 109488 130000 109608 6 key_i[3]
port 320 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 key_i[40]
port 321 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 key_i[41]
port 322 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 key_i[42]
port 323 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 key_i[43]
port 324 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 key_i[44]
port 325 nsew signal input
rlabel metal3 s 129200 63248 130000 63368 6 key_i[45]
port 326 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 key_i[46]
port 327 nsew signal input
rlabel metal2 s 92754 129200 92810 130000 6 key_i[47]
port 328 nsew signal input
rlabel metal2 s 123666 129200 123722 130000 6 key_i[48]
port 329 nsew signal input
rlabel metal2 s 14830 129200 14886 130000 6 key_i[49]
port 330 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 key_i[4]
port 331 nsew signal input
rlabel metal3 s 129200 74128 130000 74248 6 key_i[50]
port 332 nsew signal input
rlabel metal2 s 126242 129200 126298 130000 6 key_i[51]
port 333 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 key_i[52]
port 334 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 key_i[53]
port 335 nsew signal input
rlabel metal3 s 129200 38088 130000 38208 6 key_i[54]
port 336 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 key_i[55]
port 337 nsew signal input
rlabel metal2 s 110786 129200 110842 130000 6 key_i[56]
port 338 nsew signal input
rlabel metal2 s 36726 129200 36782 130000 6 key_i[57]
port 339 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 key_i[58]
port 340 nsew signal input
rlabel metal3 s 129200 75488 130000 75608 6 key_i[59]
port 341 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 key_i[5]
port 342 nsew signal input
rlabel metal3 s 129200 34008 130000 34128 6 key_i[60]
port 343 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 key_i[61]
port 344 nsew signal input
rlabel metal3 s 129200 8 130000 128 6 key_i[62]
port 345 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 key_i[63]
port 346 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 key_i[64]
port 347 nsew signal input
rlabel metal3 s 129200 53048 130000 53168 6 key_i[65]
port 348 nsew signal input
rlabel metal2 s 105634 129200 105690 130000 6 key_i[66]
port 349 nsew signal input
rlabel metal3 s 129200 113568 130000 113688 6 key_i[67]
port 350 nsew signal input
rlabel metal3 s 129200 2728 130000 2848 6 key_i[68]
port 351 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 key_i[69]
port 352 nsew signal input
rlabel metal3 s 129200 71408 130000 71528 6 key_i[6]
port 353 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 key_i[70]
port 354 nsew signal input
rlabel metal3 s 129200 117648 130000 117768 6 key_i[71]
port 355 nsew signal input
rlabel metal2 s 100482 129200 100538 130000 6 key_i[72]
port 356 nsew signal input
rlabel metal3 s 129200 10888 130000 11008 6 key_i[73]
port 357 nsew signal input
rlabel metal2 s 95330 129200 95386 130000 6 key_i[74]
port 358 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 key_i[75]
port 359 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 key_i[76]
port 360 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 key_i[77]
port 361 nsew signal input
rlabel metal2 s 18 0 74 800 6 key_i[78]
port 362 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 key_i[79]
port 363 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 key_i[7]
port 364 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 key_i[80]
port 365 nsew signal input
rlabel metal2 s 39302 129200 39358 130000 6 key_i[81]
port 366 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 key_i[82]
port 367 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 key_i[83]
port 368 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 key_i[84]
port 369 nsew signal input
rlabel metal2 s 70858 129200 70914 130000 6 key_i[85]
port 370 nsew signal input
rlabel metal2 s 41878 129200 41934 130000 6 key_i[86]
port 371 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 key_i[87]
port 372 nsew signal input
rlabel metal2 s 91466 129200 91522 130000 6 key_i[88]
port 373 nsew signal input
rlabel metal3 s 129200 32648 130000 32768 6 key_i[89]
port 374 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 key_i[8]
port 375 nsew signal input
rlabel metal3 s 129200 98608 130000 98728 6 key_i[90]
port 376 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 key_i[91]
port 377 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 key_i[92]
port 378 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 key_i[93]
port 379 nsew signal input
rlabel metal3 s 129200 94528 130000 94648 6 key_i[94]
port 380 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 key_i[95]
port 381 nsew signal input
rlabel metal2 s 87602 129200 87658 130000 6 key_i[96]
port 382 nsew signal input
rlabel metal2 s 85026 129200 85082 130000 6 key_i[97]
port 383 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 key_i[98]
port 384 nsew signal input
rlabel metal2 s 17406 129200 17462 130000 6 key_i[99]
port 385 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 key_i[9]
port 386 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 load_i
port 387 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 ready_o
port 388 nsew signal output
rlabel metal3 s 129200 61208 130000 61328 6 reset
port 389 nsew signal input
rlabel metal4 s 1944 2128 2264 127344 6 vccd1
port 390 nsew power bidirectional
rlabel metal4 s 37944 2128 38264 127344 6 vccd1
port 390 nsew power bidirectional
rlabel metal4 s 73944 2128 74264 127344 6 vccd1
port 390 nsew power bidirectional
rlabel metal4 s 109944 2128 110264 127344 6 vccd1
port 390 nsew power bidirectional
rlabel metal4 s 19944 2128 20264 127344 6 vssd1
port 391 nsew ground bidirectional
rlabel metal4 s 55944 2128 56264 127344 6 vssd1
port 391 nsew ground bidirectional
rlabel metal4 s 91944 2128 92264 127344 6 vssd1
port 391 nsew ground bidirectional
rlabel metal4 s 127944 2128 128264 127344 6 vssd1
port 391 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 130000 130000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32010330
string GDS_FILE /home/baungarten/Desktop/HW_TI_Encryption/openlane/AES_Trojan/runs/23_10_31_12_51/results/signoff/aes_Trojan.magic.gds
string GDS_START 937450
<< end >>

