// This is the unpowered netlist.
module aes_Trojan (clk,
    decrypt_i,
    load_i,
    ready_o,
    reset,
    data_i,
    data_o,
    key_i);
 input clk;
 input decrypt_i;
 input load_i;
 output ready_o;
 input reset;
 input [127:0] data_i;
 output [127:0] data_o;
 input [127:0] key_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire \addroundkey_data_o[0] ;
 wire \addroundkey_data_o[100] ;
 wire \addroundkey_data_o[101] ;
 wire \addroundkey_data_o[102] ;
 wire \addroundkey_data_o[103] ;
 wire \addroundkey_data_o[104] ;
 wire \addroundkey_data_o[105] ;
 wire \addroundkey_data_o[106] ;
 wire \addroundkey_data_o[107] ;
 wire \addroundkey_data_o[108] ;
 wire \addroundkey_data_o[109] ;
 wire \addroundkey_data_o[10] ;
 wire \addroundkey_data_o[110] ;
 wire \addroundkey_data_o[111] ;
 wire \addroundkey_data_o[112] ;
 wire \addroundkey_data_o[113] ;
 wire \addroundkey_data_o[114] ;
 wire \addroundkey_data_o[115] ;
 wire \addroundkey_data_o[116] ;
 wire \addroundkey_data_o[117] ;
 wire \addroundkey_data_o[118] ;
 wire \addroundkey_data_o[119] ;
 wire \addroundkey_data_o[11] ;
 wire \addroundkey_data_o[120] ;
 wire \addroundkey_data_o[121] ;
 wire \addroundkey_data_o[122] ;
 wire \addroundkey_data_o[123] ;
 wire \addroundkey_data_o[124] ;
 wire \addroundkey_data_o[125] ;
 wire \addroundkey_data_o[126] ;
 wire \addroundkey_data_o[127] ;
 wire \addroundkey_data_o[12] ;
 wire \addroundkey_data_o[13] ;
 wire \addroundkey_data_o[14] ;
 wire \addroundkey_data_o[15] ;
 wire \addroundkey_data_o[16] ;
 wire \addroundkey_data_o[17] ;
 wire \addroundkey_data_o[18] ;
 wire \addroundkey_data_o[19] ;
 wire \addroundkey_data_o[1] ;
 wire \addroundkey_data_o[20] ;
 wire \addroundkey_data_o[21] ;
 wire \addroundkey_data_o[22] ;
 wire \addroundkey_data_o[23] ;
 wire \addroundkey_data_o[24] ;
 wire \addroundkey_data_o[25] ;
 wire \addroundkey_data_o[26] ;
 wire \addroundkey_data_o[27] ;
 wire \addroundkey_data_o[28] ;
 wire \addroundkey_data_o[29] ;
 wire \addroundkey_data_o[2] ;
 wire \addroundkey_data_o[30] ;
 wire \addroundkey_data_o[31] ;
 wire \addroundkey_data_o[32] ;
 wire \addroundkey_data_o[33] ;
 wire \addroundkey_data_o[34] ;
 wire \addroundkey_data_o[35] ;
 wire \addroundkey_data_o[36] ;
 wire \addroundkey_data_o[37] ;
 wire \addroundkey_data_o[38] ;
 wire \addroundkey_data_o[39] ;
 wire \addroundkey_data_o[3] ;
 wire \addroundkey_data_o[40] ;
 wire \addroundkey_data_o[41] ;
 wire \addroundkey_data_o[42] ;
 wire \addroundkey_data_o[43] ;
 wire \addroundkey_data_o[44] ;
 wire \addroundkey_data_o[45] ;
 wire \addroundkey_data_o[46] ;
 wire \addroundkey_data_o[47] ;
 wire \addroundkey_data_o[48] ;
 wire \addroundkey_data_o[49] ;
 wire \addroundkey_data_o[4] ;
 wire \addroundkey_data_o[50] ;
 wire \addroundkey_data_o[51] ;
 wire \addroundkey_data_o[52] ;
 wire \addroundkey_data_o[53] ;
 wire \addroundkey_data_o[54] ;
 wire \addroundkey_data_o[55] ;
 wire \addroundkey_data_o[56] ;
 wire \addroundkey_data_o[57] ;
 wire \addroundkey_data_o[58] ;
 wire \addroundkey_data_o[59] ;
 wire \addroundkey_data_o[5] ;
 wire \addroundkey_data_o[60] ;
 wire \addroundkey_data_o[61] ;
 wire \addroundkey_data_o[62] ;
 wire \addroundkey_data_o[63] ;
 wire \addroundkey_data_o[64] ;
 wire \addroundkey_data_o[65] ;
 wire \addroundkey_data_o[66] ;
 wire \addroundkey_data_o[67] ;
 wire \addroundkey_data_o[68] ;
 wire \addroundkey_data_o[69] ;
 wire \addroundkey_data_o[6] ;
 wire \addroundkey_data_o[70] ;
 wire \addroundkey_data_o[71] ;
 wire \addroundkey_data_o[72] ;
 wire \addroundkey_data_o[73] ;
 wire \addroundkey_data_o[74] ;
 wire \addroundkey_data_o[75] ;
 wire \addroundkey_data_o[76] ;
 wire \addroundkey_data_o[77] ;
 wire \addroundkey_data_o[78] ;
 wire \addroundkey_data_o[79] ;
 wire \addroundkey_data_o[7] ;
 wire \addroundkey_data_o[80] ;
 wire \addroundkey_data_o[81] ;
 wire \addroundkey_data_o[82] ;
 wire \addroundkey_data_o[83] ;
 wire \addroundkey_data_o[84] ;
 wire \addroundkey_data_o[85] ;
 wire \addroundkey_data_o[86] ;
 wire \addroundkey_data_o[87] ;
 wire \addroundkey_data_o[88] ;
 wire \addroundkey_data_o[89] ;
 wire \addroundkey_data_o[8] ;
 wire \addroundkey_data_o[90] ;
 wire \addroundkey_data_o[91] ;
 wire \addroundkey_data_o[92] ;
 wire \addroundkey_data_o[93] ;
 wire \addroundkey_data_o[94] ;
 wire \addroundkey_data_o[95] ;
 wire \addroundkey_data_o[96] ;
 wire \addroundkey_data_o[97] ;
 wire \addroundkey_data_o[98] ;
 wire \addroundkey_data_o[99] ;
 wire \addroundkey_data_o[9] ;
 wire addroundkey_ready_o;
 wire \addroundkey_round[0] ;
 wire \addroundkey_round[1] ;
 wire \addroundkey_round[2] ;
 wire \addroundkey_round[3] ;
 wire addroundkey_start_i;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire \fifo_bank_register.bank[0][0] ;
 wire \fifo_bank_register.bank[0][100] ;
 wire \fifo_bank_register.bank[0][101] ;
 wire \fifo_bank_register.bank[0][102] ;
 wire \fifo_bank_register.bank[0][103] ;
 wire \fifo_bank_register.bank[0][104] ;
 wire \fifo_bank_register.bank[0][105] ;
 wire \fifo_bank_register.bank[0][106] ;
 wire \fifo_bank_register.bank[0][107] ;
 wire \fifo_bank_register.bank[0][108] ;
 wire \fifo_bank_register.bank[0][109] ;
 wire \fifo_bank_register.bank[0][10] ;
 wire \fifo_bank_register.bank[0][110] ;
 wire \fifo_bank_register.bank[0][111] ;
 wire \fifo_bank_register.bank[0][112] ;
 wire \fifo_bank_register.bank[0][113] ;
 wire \fifo_bank_register.bank[0][114] ;
 wire \fifo_bank_register.bank[0][115] ;
 wire \fifo_bank_register.bank[0][116] ;
 wire \fifo_bank_register.bank[0][117] ;
 wire \fifo_bank_register.bank[0][118] ;
 wire \fifo_bank_register.bank[0][119] ;
 wire \fifo_bank_register.bank[0][11] ;
 wire \fifo_bank_register.bank[0][120] ;
 wire \fifo_bank_register.bank[0][121] ;
 wire \fifo_bank_register.bank[0][122] ;
 wire \fifo_bank_register.bank[0][123] ;
 wire \fifo_bank_register.bank[0][124] ;
 wire \fifo_bank_register.bank[0][125] ;
 wire \fifo_bank_register.bank[0][126] ;
 wire \fifo_bank_register.bank[0][127] ;
 wire \fifo_bank_register.bank[0][12] ;
 wire \fifo_bank_register.bank[0][13] ;
 wire \fifo_bank_register.bank[0][14] ;
 wire \fifo_bank_register.bank[0][15] ;
 wire \fifo_bank_register.bank[0][16] ;
 wire \fifo_bank_register.bank[0][17] ;
 wire \fifo_bank_register.bank[0][18] ;
 wire \fifo_bank_register.bank[0][19] ;
 wire \fifo_bank_register.bank[0][1] ;
 wire \fifo_bank_register.bank[0][20] ;
 wire \fifo_bank_register.bank[0][21] ;
 wire \fifo_bank_register.bank[0][22] ;
 wire \fifo_bank_register.bank[0][23] ;
 wire \fifo_bank_register.bank[0][24] ;
 wire \fifo_bank_register.bank[0][25] ;
 wire \fifo_bank_register.bank[0][26] ;
 wire \fifo_bank_register.bank[0][27] ;
 wire \fifo_bank_register.bank[0][28] ;
 wire \fifo_bank_register.bank[0][29] ;
 wire \fifo_bank_register.bank[0][2] ;
 wire \fifo_bank_register.bank[0][30] ;
 wire \fifo_bank_register.bank[0][31] ;
 wire \fifo_bank_register.bank[0][32] ;
 wire \fifo_bank_register.bank[0][33] ;
 wire \fifo_bank_register.bank[0][34] ;
 wire \fifo_bank_register.bank[0][35] ;
 wire \fifo_bank_register.bank[0][36] ;
 wire \fifo_bank_register.bank[0][37] ;
 wire \fifo_bank_register.bank[0][38] ;
 wire \fifo_bank_register.bank[0][39] ;
 wire \fifo_bank_register.bank[0][3] ;
 wire \fifo_bank_register.bank[0][40] ;
 wire \fifo_bank_register.bank[0][41] ;
 wire \fifo_bank_register.bank[0][42] ;
 wire \fifo_bank_register.bank[0][43] ;
 wire \fifo_bank_register.bank[0][44] ;
 wire \fifo_bank_register.bank[0][45] ;
 wire \fifo_bank_register.bank[0][46] ;
 wire \fifo_bank_register.bank[0][47] ;
 wire \fifo_bank_register.bank[0][48] ;
 wire \fifo_bank_register.bank[0][49] ;
 wire \fifo_bank_register.bank[0][4] ;
 wire \fifo_bank_register.bank[0][50] ;
 wire \fifo_bank_register.bank[0][51] ;
 wire \fifo_bank_register.bank[0][52] ;
 wire \fifo_bank_register.bank[0][53] ;
 wire \fifo_bank_register.bank[0][54] ;
 wire \fifo_bank_register.bank[0][55] ;
 wire \fifo_bank_register.bank[0][56] ;
 wire \fifo_bank_register.bank[0][57] ;
 wire \fifo_bank_register.bank[0][58] ;
 wire \fifo_bank_register.bank[0][59] ;
 wire \fifo_bank_register.bank[0][5] ;
 wire \fifo_bank_register.bank[0][60] ;
 wire \fifo_bank_register.bank[0][61] ;
 wire \fifo_bank_register.bank[0][62] ;
 wire \fifo_bank_register.bank[0][63] ;
 wire \fifo_bank_register.bank[0][64] ;
 wire \fifo_bank_register.bank[0][65] ;
 wire \fifo_bank_register.bank[0][66] ;
 wire \fifo_bank_register.bank[0][67] ;
 wire \fifo_bank_register.bank[0][68] ;
 wire \fifo_bank_register.bank[0][69] ;
 wire \fifo_bank_register.bank[0][6] ;
 wire \fifo_bank_register.bank[0][70] ;
 wire \fifo_bank_register.bank[0][71] ;
 wire \fifo_bank_register.bank[0][72] ;
 wire \fifo_bank_register.bank[0][73] ;
 wire \fifo_bank_register.bank[0][74] ;
 wire \fifo_bank_register.bank[0][75] ;
 wire \fifo_bank_register.bank[0][76] ;
 wire \fifo_bank_register.bank[0][77] ;
 wire \fifo_bank_register.bank[0][78] ;
 wire \fifo_bank_register.bank[0][79] ;
 wire \fifo_bank_register.bank[0][7] ;
 wire \fifo_bank_register.bank[0][80] ;
 wire \fifo_bank_register.bank[0][81] ;
 wire \fifo_bank_register.bank[0][82] ;
 wire \fifo_bank_register.bank[0][83] ;
 wire \fifo_bank_register.bank[0][84] ;
 wire \fifo_bank_register.bank[0][85] ;
 wire \fifo_bank_register.bank[0][86] ;
 wire \fifo_bank_register.bank[0][87] ;
 wire \fifo_bank_register.bank[0][88] ;
 wire \fifo_bank_register.bank[0][89] ;
 wire \fifo_bank_register.bank[0][8] ;
 wire \fifo_bank_register.bank[0][90] ;
 wire \fifo_bank_register.bank[0][91] ;
 wire \fifo_bank_register.bank[0][92] ;
 wire \fifo_bank_register.bank[0][93] ;
 wire \fifo_bank_register.bank[0][94] ;
 wire \fifo_bank_register.bank[0][95] ;
 wire \fifo_bank_register.bank[0][96] ;
 wire \fifo_bank_register.bank[0][97] ;
 wire \fifo_bank_register.bank[0][98] ;
 wire \fifo_bank_register.bank[0][99] ;
 wire \fifo_bank_register.bank[0][9] ;
 wire \fifo_bank_register.bank[1][0] ;
 wire \fifo_bank_register.bank[1][100] ;
 wire \fifo_bank_register.bank[1][101] ;
 wire \fifo_bank_register.bank[1][102] ;
 wire \fifo_bank_register.bank[1][103] ;
 wire \fifo_bank_register.bank[1][104] ;
 wire \fifo_bank_register.bank[1][105] ;
 wire \fifo_bank_register.bank[1][106] ;
 wire \fifo_bank_register.bank[1][107] ;
 wire \fifo_bank_register.bank[1][108] ;
 wire \fifo_bank_register.bank[1][109] ;
 wire \fifo_bank_register.bank[1][10] ;
 wire \fifo_bank_register.bank[1][110] ;
 wire \fifo_bank_register.bank[1][111] ;
 wire \fifo_bank_register.bank[1][112] ;
 wire \fifo_bank_register.bank[1][113] ;
 wire \fifo_bank_register.bank[1][114] ;
 wire \fifo_bank_register.bank[1][115] ;
 wire \fifo_bank_register.bank[1][116] ;
 wire \fifo_bank_register.bank[1][117] ;
 wire \fifo_bank_register.bank[1][118] ;
 wire \fifo_bank_register.bank[1][119] ;
 wire \fifo_bank_register.bank[1][11] ;
 wire \fifo_bank_register.bank[1][120] ;
 wire \fifo_bank_register.bank[1][121] ;
 wire \fifo_bank_register.bank[1][122] ;
 wire \fifo_bank_register.bank[1][123] ;
 wire \fifo_bank_register.bank[1][124] ;
 wire \fifo_bank_register.bank[1][125] ;
 wire \fifo_bank_register.bank[1][126] ;
 wire \fifo_bank_register.bank[1][127] ;
 wire \fifo_bank_register.bank[1][12] ;
 wire \fifo_bank_register.bank[1][13] ;
 wire \fifo_bank_register.bank[1][14] ;
 wire \fifo_bank_register.bank[1][15] ;
 wire \fifo_bank_register.bank[1][16] ;
 wire \fifo_bank_register.bank[1][17] ;
 wire \fifo_bank_register.bank[1][18] ;
 wire \fifo_bank_register.bank[1][19] ;
 wire \fifo_bank_register.bank[1][1] ;
 wire \fifo_bank_register.bank[1][20] ;
 wire \fifo_bank_register.bank[1][21] ;
 wire \fifo_bank_register.bank[1][22] ;
 wire \fifo_bank_register.bank[1][23] ;
 wire \fifo_bank_register.bank[1][24] ;
 wire \fifo_bank_register.bank[1][25] ;
 wire \fifo_bank_register.bank[1][26] ;
 wire \fifo_bank_register.bank[1][27] ;
 wire \fifo_bank_register.bank[1][28] ;
 wire \fifo_bank_register.bank[1][29] ;
 wire \fifo_bank_register.bank[1][2] ;
 wire \fifo_bank_register.bank[1][30] ;
 wire \fifo_bank_register.bank[1][31] ;
 wire \fifo_bank_register.bank[1][32] ;
 wire \fifo_bank_register.bank[1][33] ;
 wire \fifo_bank_register.bank[1][34] ;
 wire \fifo_bank_register.bank[1][35] ;
 wire \fifo_bank_register.bank[1][36] ;
 wire \fifo_bank_register.bank[1][37] ;
 wire \fifo_bank_register.bank[1][38] ;
 wire \fifo_bank_register.bank[1][39] ;
 wire \fifo_bank_register.bank[1][3] ;
 wire \fifo_bank_register.bank[1][40] ;
 wire \fifo_bank_register.bank[1][41] ;
 wire \fifo_bank_register.bank[1][42] ;
 wire \fifo_bank_register.bank[1][43] ;
 wire \fifo_bank_register.bank[1][44] ;
 wire \fifo_bank_register.bank[1][45] ;
 wire \fifo_bank_register.bank[1][46] ;
 wire \fifo_bank_register.bank[1][47] ;
 wire \fifo_bank_register.bank[1][48] ;
 wire \fifo_bank_register.bank[1][49] ;
 wire \fifo_bank_register.bank[1][4] ;
 wire \fifo_bank_register.bank[1][50] ;
 wire \fifo_bank_register.bank[1][51] ;
 wire \fifo_bank_register.bank[1][52] ;
 wire \fifo_bank_register.bank[1][53] ;
 wire \fifo_bank_register.bank[1][54] ;
 wire \fifo_bank_register.bank[1][55] ;
 wire \fifo_bank_register.bank[1][56] ;
 wire \fifo_bank_register.bank[1][57] ;
 wire \fifo_bank_register.bank[1][58] ;
 wire \fifo_bank_register.bank[1][59] ;
 wire \fifo_bank_register.bank[1][5] ;
 wire \fifo_bank_register.bank[1][60] ;
 wire \fifo_bank_register.bank[1][61] ;
 wire \fifo_bank_register.bank[1][62] ;
 wire \fifo_bank_register.bank[1][63] ;
 wire \fifo_bank_register.bank[1][64] ;
 wire \fifo_bank_register.bank[1][65] ;
 wire \fifo_bank_register.bank[1][66] ;
 wire \fifo_bank_register.bank[1][67] ;
 wire \fifo_bank_register.bank[1][68] ;
 wire \fifo_bank_register.bank[1][69] ;
 wire \fifo_bank_register.bank[1][6] ;
 wire \fifo_bank_register.bank[1][70] ;
 wire \fifo_bank_register.bank[1][71] ;
 wire \fifo_bank_register.bank[1][72] ;
 wire \fifo_bank_register.bank[1][73] ;
 wire \fifo_bank_register.bank[1][74] ;
 wire \fifo_bank_register.bank[1][75] ;
 wire \fifo_bank_register.bank[1][76] ;
 wire \fifo_bank_register.bank[1][77] ;
 wire \fifo_bank_register.bank[1][78] ;
 wire \fifo_bank_register.bank[1][79] ;
 wire \fifo_bank_register.bank[1][7] ;
 wire \fifo_bank_register.bank[1][80] ;
 wire \fifo_bank_register.bank[1][81] ;
 wire \fifo_bank_register.bank[1][82] ;
 wire \fifo_bank_register.bank[1][83] ;
 wire \fifo_bank_register.bank[1][84] ;
 wire \fifo_bank_register.bank[1][85] ;
 wire \fifo_bank_register.bank[1][86] ;
 wire \fifo_bank_register.bank[1][87] ;
 wire \fifo_bank_register.bank[1][88] ;
 wire \fifo_bank_register.bank[1][89] ;
 wire \fifo_bank_register.bank[1][8] ;
 wire \fifo_bank_register.bank[1][90] ;
 wire \fifo_bank_register.bank[1][91] ;
 wire \fifo_bank_register.bank[1][92] ;
 wire \fifo_bank_register.bank[1][93] ;
 wire \fifo_bank_register.bank[1][94] ;
 wire \fifo_bank_register.bank[1][95] ;
 wire \fifo_bank_register.bank[1][96] ;
 wire \fifo_bank_register.bank[1][97] ;
 wire \fifo_bank_register.bank[1][98] ;
 wire \fifo_bank_register.bank[1][99] ;
 wire \fifo_bank_register.bank[1][9] ;
 wire \fifo_bank_register.bank[2][0] ;
 wire \fifo_bank_register.bank[2][100] ;
 wire \fifo_bank_register.bank[2][101] ;
 wire \fifo_bank_register.bank[2][102] ;
 wire \fifo_bank_register.bank[2][103] ;
 wire \fifo_bank_register.bank[2][104] ;
 wire \fifo_bank_register.bank[2][105] ;
 wire \fifo_bank_register.bank[2][106] ;
 wire \fifo_bank_register.bank[2][107] ;
 wire \fifo_bank_register.bank[2][108] ;
 wire \fifo_bank_register.bank[2][109] ;
 wire \fifo_bank_register.bank[2][10] ;
 wire \fifo_bank_register.bank[2][110] ;
 wire \fifo_bank_register.bank[2][111] ;
 wire \fifo_bank_register.bank[2][112] ;
 wire \fifo_bank_register.bank[2][113] ;
 wire \fifo_bank_register.bank[2][114] ;
 wire \fifo_bank_register.bank[2][115] ;
 wire \fifo_bank_register.bank[2][116] ;
 wire \fifo_bank_register.bank[2][117] ;
 wire \fifo_bank_register.bank[2][118] ;
 wire \fifo_bank_register.bank[2][119] ;
 wire \fifo_bank_register.bank[2][11] ;
 wire \fifo_bank_register.bank[2][120] ;
 wire \fifo_bank_register.bank[2][121] ;
 wire \fifo_bank_register.bank[2][122] ;
 wire \fifo_bank_register.bank[2][123] ;
 wire \fifo_bank_register.bank[2][124] ;
 wire \fifo_bank_register.bank[2][125] ;
 wire \fifo_bank_register.bank[2][126] ;
 wire \fifo_bank_register.bank[2][127] ;
 wire \fifo_bank_register.bank[2][12] ;
 wire \fifo_bank_register.bank[2][13] ;
 wire \fifo_bank_register.bank[2][14] ;
 wire \fifo_bank_register.bank[2][15] ;
 wire \fifo_bank_register.bank[2][16] ;
 wire \fifo_bank_register.bank[2][17] ;
 wire \fifo_bank_register.bank[2][18] ;
 wire \fifo_bank_register.bank[2][19] ;
 wire \fifo_bank_register.bank[2][1] ;
 wire \fifo_bank_register.bank[2][20] ;
 wire \fifo_bank_register.bank[2][21] ;
 wire \fifo_bank_register.bank[2][22] ;
 wire \fifo_bank_register.bank[2][23] ;
 wire \fifo_bank_register.bank[2][24] ;
 wire \fifo_bank_register.bank[2][25] ;
 wire \fifo_bank_register.bank[2][26] ;
 wire \fifo_bank_register.bank[2][27] ;
 wire \fifo_bank_register.bank[2][28] ;
 wire \fifo_bank_register.bank[2][29] ;
 wire \fifo_bank_register.bank[2][2] ;
 wire \fifo_bank_register.bank[2][30] ;
 wire \fifo_bank_register.bank[2][31] ;
 wire \fifo_bank_register.bank[2][32] ;
 wire \fifo_bank_register.bank[2][33] ;
 wire \fifo_bank_register.bank[2][34] ;
 wire \fifo_bank_register.bank[2][35] ;
 wire \fifo_bank_register.bank[2][36] ;
 wire \fifo_bank_register.bank[2][37] ;
 wire \fifo_bank_register.bank[2][38] ;
 wire \fifo_bank_register.bank[2][39] ;
 wire \fifo_bank_register.bank[2][3] ;
 wire \fifo_bank_register.bank[2][40] ;
 wire \fifo_bank_register.bank[2][41] ;
 wire \fifo_bank_register.bank[2][42] ;
 wire \fifo_bank_register.bank[2][43] ;
 wire \fifo_bank_register.bank[2][44] ;
 wire \fifo_bank_register.bank[2][45] ;
 wire \fifo_bank_register.bank[2][46] ;
 wire \fifo_bank_register.bank[2][47] ;
 wire \fifo_bank_register.bank[2][48] ;
 wire \fifo_bank_register.bank[2][49] ;
 wire \fifo_bank_register.bank[2][4] ;
 wire \fifo_bank_register.bank[2][50] ;
 wire \fifo_bank_register.bank[2][51] ;
 wire \fifo_bank_register.bank[2][52] ;
 wire \fifo_bank_register.bank[2][53] ;
 wire \fifo_bank_register.bank[2][54] ;
 wire \fifo_bank_register.bank[2][55] ;
 wire \fifo_bank_register.bank[2][56] ;
 wire \fifo_bank_register.bank[2][57] ;
 wire \fifo_bank_register.bank[2][58] ;
 wire \fifo_bank_register.bank[2][59] ;
 wire \fifo_bank_register.bank[2][5] ;
 wire \fifo_bank_register.bank[2][60] ;
 wire \fifo_bank_register.bank[2][61] ;
 wire \fifo_bank_register.bank[2][62] ;
 wire \fifo_bank_register.bank[2][63] ;
 wire \fifo_bank_register.bank[2][64] ;
 wire \fifo_bank_register.bank[2][65] ;
 wire \fifo_bank_register.bank[2][66] ;
 wire \fifo_bank_register.bank[2][67] ;
 wire \fifo_bank_register.bank[2][68] ;
 wire \fifo_bank_register.bank[2][69] ;
 wire \fifo_bank_register.bank[2][6] ;
 wire \fifo_bank_register.bank[2][70] ;
 wire \fifo_bank_register.bank[2][71] ;
 wire \fifo_bank_register.bank[2][72] ;
 wire \fifo_bank_register.bank[2][73] ;
 wire \fifo_bank_register.bank[2][74] ;
 wire \fifo_bank_register.bank[2][75] ;
 wire \fifo_bank_register.bank[2][76] ;
 wire \fifo_bank_register.bank[2][77] ;
 wire \fifo_bank_register.bank[2][78] ;
 wire \fifo_bank_register.bank[2][79] ;
 wire \fifo_bank_register.bank[2][7] ;
 wire \fifo_bank_register.bank[2][80] ;
 wire \fifo_bank_register.bank[2][81] ;
 wire \fifo_bank_register.bank[2][82] ;
 wire \fifo_bank_register.bank[2][83] ;
 wire \fifo_bank_register.bank[2][84] ;
 wire \fifo_bank_register.bank[2][85] ;
 wire \fifo_bank_register.bank[2][86] ;
 wire \fifo_bank_register.bank[2][87] ;
 wire \fifo_bank_register.bank[2][88] ;
 wire \fifo_bank_register.bank[2][89] ;
 wire \fifo_bank_register.bank[2][8] ;
 wire \fifo_bank_register.bank[2][90] ;
 wire \fifo_bank_register.bank[2][91] ;
 wire \fifo_bank_register.bank[2][92] ;
 wire \fifo_bank_register.bank[2][93] ;
 wire \fifo_bank_register.bank[2][94] ;
 wire \fifo_bank_register.bank[2][95] ;
 wire \fifo_bank_register.bank[2][96] ;
 wire \fifo_bank_register.bank[2][97] ;
 wire \fifo_bank_register.bank[2][98] ;
 wire \fifo_bank_register.bank[2][99] ;
 wire \fifo_bank_register.bank[2][9] ;
 wire \fifo_bank_register.bank[3][0] ;
 wire \fifo_bank_register.bank[3][100] ;
 wire \fifo_bank_register.bank[3][101] ;
 wire \fifo_bank_register.bank[3][102] ;
 wire \fifo_bank_register.bank[3][103] ;
 wire \fifo_bank_register.bank[3][104] ;
 wire \fifo_bank_register.bank[3][105] ;
 wire \fifo_bank_register.bank[3][106] ;
 wire \fifo_bank_register.bank[3][107] ;
 wire \fifo_bank_register.bank[3][108] ;
 wire \fifo_bank_register.bank[3][109] ;
 wire \fifo_bank_register.bank[3][10] ;
 wire \fifo_bank_register.bank[3][110] ;
 wire \fifo_bank_register.bank[3][111] ;
 wire \fifo_bank_register.bank[3][112] ;
 wire \fifo_bank_register.bank[3][113] ;
 wire \fifo_bank_register.bank[3][114] ;
 wire \fifo_bank_register.bank[3][115] ;
 wire \fifo_bank_register.bank[3][116] ;
 wire \fifo_bank_register.bank[3][117] ;
 wire \fifo_bank_register.bank[3][118] ;
 wire \fifo_bank_register.bank[3][119] ;
 wire \fifo_bank_register.bank[3][11] ;
 wire \fifo_bank_register.bank[3][120] ;
 wire \fifo_bank_register.bank[3][121] ;
 wire \fifo_bank_register.bank[3][122] ;
 wire \fifo_bank_register.bank[3][123] ;
 wire \fifo_bank_register.bank[3][124] ;
 wire \fifo_bank_register.bank[3][125] ;
 wire \fifo_bank_register.bank[3][126] ;
 wire \fifo_bank_register.bank[3][127] ;
 wire \fifo_bank_register.bank[3][12] ;
 wire \fifo_bank_register.bank[3][13] ;
 wire \fifo_bank_register.bank[3][14] ;
 wire \fifo_bank_register.bank[3][15] ;
 wire \fifo_bank_register.bank[3][16] ;
 wire \fifo_bank_register.bank[3][17] ;
 wire \fifo_bank_register.bank[3][18] ;
 wire \fifo_bank_register.bank[3][19] ;
 wire \fifo_bank_register.bank[3][1] ;
 wire \fifo_bank_register.bank[3][20] ;
 wire \fifo_bank_register.bank[3][21] ;
 wire \fifo_bank_register.bank[3][22] ;
 wire \fifo_bank_register.bank[3][23] ;
 wire \fifo_bank_register.bank[3][24] ;
 wire \fifo_bank_register.bank[3][25] ;
 wire \fifo_bank_register.bank[3][26] ;
 wire \fifo_bank_register.bank[3][27] ;
 wire \fifo_bank_register.bank[3][28] ;
 wire \fifo_bank_register.bank[3][29] ;
 wire \fifo_bank_register.bank[3][2] ;
 wire \fifo_bank_register.bank[3][30] ;
 wire \fifo_bank_register.bank[3][31] ;
 wire \fifo_bank_register.bank[3][32] ;
 wire \fifo_bank_register.bank[3][33] ;
 wire \fifo_bank_register.bank[3][34] ;
 wire \fifo_bank_register.bank[3][35] ;
 wire \fifo_bank_register.bank[3][36] ;
 wire \fifo_bank_register.bank[3][37] ;
 wire \fifo_bank_register.bank[3][38] ;
 wire \fifo_bank_register.bank[3][39] ;
 wire \fifo_bank_register.bank[3][3] ;
 wire \fifo_bank_register.bank[3][40] ;
 wire \fifo_bank_register.bank[3][41] ;
 wire \fifo_bank_register.bank[3][42] ;
 wire \fifo_bank_register.bank[3][43] ;
 wire \fifo_bank_register.bank[3][44] ;
 wire \fifo_bank_register.bank[3][45] ;
 wire \fifo_bank_register.bank[3][46] ;
 wire \fifo_bank_register.bank[3][47] ;
 wire \fifo_bank_register.bank[3][48] ;
 wire \fifo_bank_register.bank[3][49] ;
 wire \fifo_bank_register.bank[3][4] ;
 wire \fifo_bank_register.bank[3][50] ;
 wire \fifo_bank_register.bank[3][51] ;
 wire \fifo_bank_register.bank[3][52] ;
 wire \fifo_bank_register.bank[3][53] ;
 wire \fifo_bank_register.bank[3][54] ;
 wire \fifo_bank_register.bank[3][55] ;
 wire \fifo_bank_register.bank[3][56] ;
 wire \fifo_bank_register.bank[3][57] ;
 wire \fifo_bank_register.bank[3][58] ;
 wire \fifo_bank_register.bank[3][59] ;
 wire \fifo_bank_register.bank[3][5] ;
 wire \fifo_bank_register.bank[3][60] ;
 wire \fifo_bank_register.bank[3][61] ;
 wire \fifo_bank_register.bank[3][62] ;
 wire \fifo_bank_register.bank[3][63] ;
 wire \fifo_bank_register.bank[3][64] ;
 wire \fifo_bank_register.bank[3][65] ;
 wire \fifo_bank_register.bank[3][66] ;
 wire \fifo_bank_register.bank[3][67] ;
 wire \fifo_bank_register.bank[3][68] ;
 wire \fifo_bank_register.bank[3][69] ;
 wire \fifo_bank_register.bank[3][6] ;
 wire \fifo_bank_register.bank[3][70] ;
 wire \fifo_bank_register.bank[3][71] ;
 wire \fifo_bank_register.bank[3][72] ;
 wire \fifo_bank_register.bank[3][73] ;
 wire \fifo_bank_register.bank[3][74] ;
 wire \fifo_bank_register.bank[3][75] ;
 wire \fifo_bank_register.bank[3][76] ;
 wire \fifo_bank_register.bank[3][77] ;
 wire \fifo_bank_register.bank[3][78] ;
 wire \fifo_bank_register.bank[3][79] ;
 wire \fifo_bank_register.bank[3][7] ;
 wire \fifo_bank_register.bank[3][80] ;
 wire \fifo_bank_register.bank[3][81] ;
 wire \fifo_bank_register.bank[3][82] ;
 wire \fifo_bank_register.bank[3][83] ;
 wire \fifo_bank_register.bank[3][84] ;
 wire \fifo_bank_register.bank[3][85] ;
 wire \fifo_bank_register.bank[3][86] ;
 wire \fifo_bank_register.bank[3][87] ;
 wire \fifo_bank_register.bank[3][88] ;
 wire \fifo_bank_register.bank[3][89] ;
 wire \fifo_bank_register.bank[3][8] ;
 wire \fifo_bank_register.bank[3][90] ;
 wire \fifo_bank_register.bank[3][91] ;
 wire \fifo_bank_register.bank[3][92] ;
 wire \fifo_bank_register.bank[3][93] ;
 wire \fifo_bank_register.bank[3][94] ;
 wire \fifo_bank_register.bank[3][95] ;
 wire \fifo_bank_register.bank[3][96] ;
 wire \fifo_bank_register.bank[3][97] ;
 wire \fifo_bank_register.bank[3][98] ;
 wire \fifo_bank_register.bank[3][99] ;
 wire \fifo_bank_register.bank[3][9] ;
 wire \fifo_bank_register.bank[4][0] ;
 wire \fifo_bank_register.bank[4][100] ;
 wire \fifo_bank_register.bank[4][101] ;
 wire \fifo_bank_register.bank[4][102] ;
 wire \fifo_bank_register.bank[4][103] ;
 wire \fifo_bank_register.bank[4][104] ;
 wire \fifo_bank_register.bank[4][105] ;
 wire \fifo_bank_register.bank[4][106] ;
 wire \fifo_bank_register.bank[4][107] ;
 wire \fifo_bank_register.bank[4][108] ;
 wire \fifo_bank_register.bank[4][109] ;
 wire \fifo_bank_register.bank[4][10] ;
 wire \fifo_bank_register.bank[4][110] ;
 wire \fifo_bank_register.bank[4][111] ;
 wire \fifo_bank_register.bank[4][112] ;
 wire \fifo_bank_register.bank[4][113] ;
 wire \fifo_bank_register.bank[4][114] ;
 wire \fifo_bank_register.bank[4][115] ;
 wire \fifo_bank_register.bank[4][116] ;
 wire \fifo_bank_register.bank[4][117] ;
 wire \fifo_bank_register.bank[4][118] ;
 wire \fifo_bank_register.bank[4][119] ;
 wire \fifo_bank_register.bank[4][11] ;
 wire \fifo_bank_register.bank[4][120] ;
 wire \fifo_bank_register.bank[4][121] ;
 wire \fifo_bank_register.bank[4][122] ;
 wire \fifo_bank_register.bank[4][123] ;
 wire \fifo_bank_register.bank[4][124] ;
 wire \fifo_bank_register.bank[4][125] ;
 wire \fifo_bank_register.bank[4][126] ;
 wire \fifo_bank_register.bank[4][127] ;
 wire \fifo_bank_register.bank[4][12] ;
 wire \fifo_bank_register.bank[4][13] ;
 wire \fifo_bank_register.bank[4][14] ;
 wire \fifo_bank_register.bank[4][15] ;
 wire \fifo_bank_register.bank[4][16] ;
 wire \fifo_bank_register.bank[4][17] ;
 wire \fifo_bank_register.bank[4][18] ;
 wire \fifo_bank_register.bank[4][19] ;
 wire \fifo_bank_register.bank[4][1] ;
 wire \fifo_bank_register.bank[4][20] ;
 wire \fifo_bank_register.bank[4][21] ;
 wire \fifo_bank_register.bank[4][22] ;
 wire \fifo_bank_register.bank[4][23] ;
 wire \fifo_bank_register.bank[4][24] ;
 wire \fifo_bank_register.bank[4][25] ;
 wire \fifo_bank_register.bank[4][26] ;
 wire \fifo_bank_register.bank[4][27] ;
 wire \fifo_bank_register.bank[4][28] ;
 wire \fifo_bank_register.bank[4][29] ;
 wire \fifo_bank_register.bank[4][2] ;
 wire \fifo_bank_register.bank[4][30] ;
 wire \fifo_bank_register.bank[4][31] ;
 wire \fifo_bank_register.bank[4][32] ;
 wire \fifo_bank_register.bank[4][33] ;
 wire \fifo_bank_register.bank[4][34] ;
 wire \fifo_bank_register.bank[4][35] ;
 wire \fifo_bank_register.bank[4][36] ;
 wire \fifo_bank_register.bank[4][37] ;
 wire \fifo_bank_register.bank[4][38] ;
 wire \fifo_bank_register.bank[4][39] ;
 wire \fifo_bank_register.bank[4][3] ;
 wire \fifo_bank_register.bank[4][40] ;
 wire \fifo_bank_register.bank[4][41] ;
 wire \fifo_bank_register.bank[4][42] ;
 wire \fifo_bank_register.bank[4][43] ;
 wire \fifo_bank_register.bank[4][44] ;
 wire \fifo_bank_register.bank[4][45] ;
 wire \fifo_bank_register.bank[4][46] ;
 wire \fifo_bank_register.bank[4][47] ;
 wire \fifo_bank_register.bank[4][48] ;
 wire \fifo_bank_register.bank[4][49] ;
 wire \fifo_bank_register.bank[4][4] ;
 wire \fifo_bank_register.bank[4][50] ;
 wire \fifo_bank_register.bank[4][51] ;
 wire \fifo_bank_register.bank[4][52] ;
 wire \fifo_bank_register.bank[4][53] ;
 wire \fifo_bank_register.bank[4][54] ;
 wire \fifo_bank_register.bank[4][55] ;
 wire \fifo_bank_register.bank[4][56] ;
 wire \fifo_bank_register.bank[4][57] ;
 wire \fifo_bank_register.bank[4][58] ;
 wire \fifo_bank_register.bank[4][59] ;
 wire \fifo_bank_register.bank[4][5] ;
 wire \fifo_bank_register.bank[4][60] ;
 wire \fifo_bank_register.bank[4][61] ;
 wire \fifo_bank_register.bank[4][62] ;
 wire \fifo_bank_register.bank[4][63] ;
 wire \fifo_bank_register.bank[4][64] ;
 wire \fifo_bank_register.bank[4][65] ;
 wire \fifo_bank_register.bank[4][66] ;
 wire \fifo_bank_register.bank[4][67] ;
 wire \fifo_bank_register.bank[4][68] ;
 wire \fifo_bank_register.bank[4][69] ;
 wire \fifo_bank_register.bank[4][6] ;
 wire \fifo_bank_register.bank[4][70] ;
 wire \fifo_bank_register.bank[4][71] ;
 wire \fifo_bank_register.bank[4][72] ;
 wire \fifo_bank_register.bank[4][73] ;
 wire \fifo_bank_register.bank[4][74] ;
 wire \fifo_bank_register.bank[4][75] ;
 wire \fifo_bank_register.bank[4][76] ;
 wire \fifo_bank_register.bank[4][77] ;
 wire \fifo_bank_register.bank[4][78] ;
 wire \fifo_bank_register.bank[4][79] ;
 wire \fifo_bank_register.bank[4][7] ;
 wire \fifo_bank_register.bank[4][80] ;
 wire \fifo_bank_register.bank[4][81] ;
 wire \fifo_bank_register.bank[4][82] ;
 wire \fifo_bank_register.bank[4][83] ;
 wire \fifo_bank_register.bank[4][84] ;
 wire \fifo_bank_register.bank[4][85] ;
 wire \fifo_bank_register.bank[4][86] ;
 wire \fifo_bank_register.bank[4][87] ;
 wire \fifo_bank_register.bank[4][88] ;
 wire \fifo_bank_register.bank[4][89] ;
 wire \fifo_bank_register.bank[4][8] ;
 wire \fifo_bank_register.bank[4][90] ;
 wire \fifo_bank_register.bank[4][91] ;
 wire \fifo_bank_register.bank[4][92] ;
 wire \fifo_bank_register.bank[4][93] ;
 wire \fifo_bank_register.bank[4][94] ;
 wire \fifo_bank_register.bank[4][95] ;
 wire \fifo_bank_register.bank[4][96] ;
 wire \fifo_bank_register.bank[4][97] ;
 wire \fifo_bank_register.bank[4][98] ;
 wire \fifo_bank_register.bank[4][99] ;
 wire \fifo_bank_register.bank[4][9] ;
 wire \fifo_bank_register.bank[5][0] ;
 wire \fifo_bank_register.bank[5][100] ;
 wire \fifo_bank_register.bank[5][101] ;
 wire \fifo_bank_register.bank[5][102] ;
 wire \fifo_bank_register.bank[5][103] ;
 wire \fifo_bank_register.bank[5][104] ;
 wire \fifo_bank_register.bank[5][105] ;
 wire \fifo_bank_register.bank[5][106] ;
 wire \fifo_bank_register.bank[5][107] ;
 wire \fifo_bank_register.bank[5][108] ;
 wire \fifo_bank_register.bank[5][109] ;
 wire \fifo_bank_register.bank[5][10] ;
 wire \fifo_bank_register.bank[5][110] ;
 wire \fifo_bank_register.bank[5][111] ;
 wire \fifo_bank_register.bank[5][112] ;
 wire \fifo_bank_register.bank[5][113] ;
 wire \fifo_bank_register.bank[5][114] ;
 wire \fifo_bank_register.bank[5][115] ;
 wire \fifo_bank_register.bank[5][116] ;
 wire \fifo_bank_register.bank[5][117] ;
 wire \fifo_bank_register.bank[5][118] ;
 wire \fifo_bank_register.bank[5][119] ;
 wire \fifo_bank_register.bank[5][11] ;
 wire \fifo_bank_register.bank[5][120] ;
 wire \fifo_bank_register.bank[5][121] ;
 wire \fifo_bank_register.bank[5][122] ;
 wire \fifo_bank_register.bank[5][123] ;
 wire \fifo_bank_register.bank[5][124] ;
 wire \fifo_bank_register.bank[5][125] ;
 wire \fifo_bank_register.bank[5][126] ;
 wire \fifo_bank_register.bank[5][127] ;
 wire \fifo_bank_register.bank[5][12] ;
 wire \fifo_bank_register.bank[5][13] ;
 wire \fifo_bank_register.bank[5][14] ;
 wire \fifo_bank_register.bank[5][15] ;
 wire \fifo_bank_register.bank[5][16] ;
 wire \fifo_bank_register.bank[5][17] ;
 wire \fifo_bank_register.bank[5][18] ;
 wire \fifo_bank_register.bank[5][19] ;
 wire \fifo_bank_register.bank[5][1] ;
 wire \fifo_bank_register.bank[5][20] ;
 wire \fifo_bank_register.bank[5][21] ;
 wire \fifo_bank_register.bank[5][22] ;
 wire \fifo_bank_register.bank[5][23] ;
 wire \fifo_bank_register.bank[5][24] ;
 wire \fifo_bank_register.bank[5][25] ;
 wire \fifo_bank_register.bank[5][26] ;
 wire \fifo_bank_register.bank[5][27] ;
 wire \fifo_bank_register.bank[5][28] ;
 wire \fifo_bank_register.bank[5][29] ;
 wire \fifo_bank_register.bank[5][2] ;
 wire \fifo_bank_register.bank[5][30] ;
 wire \fifo_bank_register.bank[5][31] ;
 wire \fifo_bank_register.bank[5][32] ;
 wire \fifo_bank_register.bank[5][33] ;
 wire \fifo_bank_register.bank[5][34] ;
 wire \fifo_bank_register.bank[5][35] ;
 wire \fifo_bank_register.bank[5][36] ;
 wire \fifo_bank_register.bank[5][37] ;
 wire \fifo_bank_register.bank[5][38] ;
 wire \fifo_bank_register.bank[5][39] ;
 wire \fifo_bank_register.bank[5][3] ;
 wire \fifo_bank_register.bank[5][40] ;
 wire \fifo_bank_register.bank[5][41] ;
 wire \fifo_bank_register.bank[5][42] ;
 wire \fifo_bank_register.bank[5][43] ;
 wire \fifo_bank_register.bank[5][44] ;
 wire \fifo_bank_register.bank[5][45] ;
 wire \fifo_bank_register.bank[5][46] ;
 wire \fifo_bank_register.bank[5][47] ;
 wire \fifo_bank_register.bank[5][48] ;
 wire \fifo_bank_register.bank[5][49] ;
 wire \fifo_bank_register.bank[5][4] ;
 wire \fifo_bank_register.bank[5][50] ;
 wire \fifo_bank_register.bank[5][51] ;
 wire \fifo_bank_register.bank[5][52] ;
 wire \fifo_bank_register.bank[5][53] ;
 wire \fifo_bank_register.bank[5][54] ;
 wire \fifo_bank_register.bank[5][55] ;
 wire \fifo_bank_register.bank[5][56] ;
 wire \fifo_bank_register.bank[5][57] ;
 wire \fifo_bank_register.bank[5][58] ;
 wire \fifo_bank_register.bank[5][59] ;
 wire \fifo_bank_register.bank[5][5] ;
 wire \fifo_bank_register.bank[5][60] ;
 wire \fifo_bank_register.bank[5][61] ;
 wire \fifo_bank_register.bank[5][62] ;
 wire \fifo_bank_register.bank[5][63] ;
 wire \fifo_bank_register.bank[5][64] ;
 wire \fifo_bank_register.bank[5][65] ;
 wire \fifo_bank_register.bank[5][66] ;
 wire \fifo_bank_register.bank[5][67] ;
 wire \fifo_bank_register.bank[5][68] ;
 wire \fifo_bank_register.bank[5][69] ;
 wire \fifo_bank_register.bank[5][6] ;
 wire \fifo_bank_register.bank[5][70] ;
 wire \fifo_bank_register.bank[5][71] ;
 wire \fifo_bank_register.bank[5][72] ;
 wire \fifo_bank_register.bank[5][73] ;
 wire \fifo_bank_register.bank[5][74] ;
 wire \fifo_bank_register.bank[5][75] ;
 wire \fifo_bank_register.bank[5][76] ;
 wire \fifo_bank_register.bank[5][77] ;
 wire \fifo_bank_register.bank[5][78] ;
 wire \fifo_bank_register.bank[5][79] ;
 wire \fifo_bank_register.bank[5][7] ;
 wire \fifo_bank_register.bank[5][80] ;
 wire \fifo_bank_register.bank[5][81] ;
 wire \fifo_bank_register.bank[5][82] ;
 wire \fifo_bank_register.bank[5][83] ;
 wire \fifo_bank_register.bank[5][84] ;
 wire \fifo_bank_register.bank[5][85] ;
 wire \fifo_bank_register.bank[5][86] ;
 wire \fifo_bank_register.bank[5][87] ;
 wire \fifo_bank_register.bank[5][88] ;
 wire \fifo_bank_register.bank[5][89] ;
 wire \fifo_bank_register.bank[5][8] ;
 wire \fifo_bank_register.bank[5][90] ;
 wire \fifo_bank_register.bank[5][91] ;
 wire \fifo_bank_register.bank[5][92] ;
 wire \fifo_bank_register.bank[5][93] ;
 wire \fifo_bank_register.bank[5][94] ;
 wire \fifo_bank_register.bank[5][95] ;
 wire \fifo_bank_register.bank[5][96] ;
 wire \fifo_bank_register.bank[5][97] ;
 wire \fifo_bank_register.bank[5][98] ;
 wire \fifo_bank_register.bank[5][99] ;
 wire \fifo_bank_register.bank[5][9] ;
 wire \fifo_bank_register.bank[6][0] ;
 wire \fifo_bank_register.bank[6][100] ;
 wire \fifo_bank_register.bank[6][101] ;
 wire \fifo_bank_register.bank[6][102] ;
 wire \fifo_bank_register.bank[6][103] ;
 wire \fifo_bank_register.bank[6][104] ;
 wire \fifo_bank_register.bank[6][105] ;
 wire \fifo_bank_register.bank[6][106] ;
 wire \fifo_bank_register.bank[6][107] ;
 wire \fifo_bank_register.bank[6][108] ;
 wire \fifo_bank_register.bank[6][109] ;
 wire \fifo_bank_register.bank[6][10] ;
 wire \fifo_bank_register.bank[6][110] ;
 wire \fifo_bank_register.bank[6][111] ;
 wire \fifo_bank_register.bank[6][112] ;
 wire \fifo_bank_register.bank[6][113] ;
 wire \fifo_bank_register.bank[6][114] ;
 wire \fifo_bank_register.bank[6][115] ;
 wire \fifo_bank_register.bank[6][116] ;
 wire \fifo_bank_register.bank[6][117] ;
 wire \fifo_bank_register.bank[6][118] ;
 wire \fifo_bank_register.bank[6][119] ;
 wire \fifo_bank_register.bank[6][11] ;
 wire \fifo_bank_register.bank[6][120] ;
 wire \fifo_bank_register.bank[6][121] ;
 wire \fifo_bank_register.bank[6][122] ;
 wire \fifo_bank_register.bank[6][123] ;
 wire \fifo_bank_register.bank[6][124] ;
 wire \fifo_bank_register.bank[6][125] ;
 wire \fifo_bank_register.bank[6][126] ;
 wire \fifo_bank_register.bank[6][127] ;
 wire \fifo_bank_register.bank[6][12] ;
 wire \fifo_bank_register.bank[6][13] ;
 wire \fifo_bank_register.bank[6][14] ;
 wire \fifo_bank_register.bank[6][15] ;
 wire \fifo_bank_register.bank[6][16] ;
 wire \fifo_bank_register.bank[6][17] ;
 wire \fifo_bank_register.bank[6][18] ;
 wire \fifo_bank_register.bank[6][19] ;
 wire \fifo_bank_register.bank[6][1] ;
 wire \fifo_bank_register.bank[6][20] ;
 wire \fifo_bank_register.bank[6][21] ;
 wire \fifo_bank_register.bank[6][22] ;
 wire \fifo_bank_register.bank[6][23] ;
 wire \fifo_bank_register.bank[6][24] ;
 wire \fifo_bank_register.bank[6][25] ;
 wire \fifo_bank_register.bank[6][26] ;
 wire \fifo_bank_register.bank[6][27] ;
 wire \fifo_bank_register.bank[6][28] ;
 wire \fifo_bank_register.bank[6][29] ;
 wire \fifo_bank_register.bank[6][2] ;
 wire \fifo_bank_register.bank[6][30] ;
 wire \fifo_bank_register.bank[6][31] ;
 wire \fifo_bank_register.bank[6][32] ;
 wire \fifo_bank_register.bank[6][33] ;
 wire \fifo_bank_register.bank[6][34] ;
 wire \fifo_bank_register.bank[6][35] ;
 wire \fifo_bank_register.bank[6][36] ;
 wire \fifo_bank_register.bank[6][37] ;
 wire \fifo_bank_register.bank[6][38] ;
 wire \fifo_bank_register.bank[6][39] ;
 wire \fifo_bank_register.bank[6][3] ;
 wire \fifo_bank_register.bank[6][40] ;
 wire \fifo_bank_register.bank[6][41] ;
 wire \fifo_bank_register.bank[6][42] ;
 wire \fifo_bank_register.bank[6][43] ;
 wire \fifo_bank_register.bank[6][44] ;
 wire \fifo_bank_register.bank[6][45] ;
 wire \fifo_bank_register.bank[6][46] ;
 wire \fifo_bank_register.bank[6][47] ;
 wire \fifo_bank_register.bank[6][48] ;
 wire \fifo_bank_register.bank[6][49] ;
 wire \fifo_bank_register.bank[6][4] ;
 wire \fifo_bank_register.bank[6][50] ;
 wire \fifo_bank_register.bank[6][51] ;
 wire \fifo_bank_register.bank[6][52] ;
 wire \fifo_bank_register.bank[6][53] ;
 wire \fifo_bank_register.bank[6][54] ;
 wire \fifo_bank_register.bank[6][55] ;
 wire \fifo_bank_register.bank[6][56] ;
 wire \fifo_bank_register.bank[6][57] ;
 wire \fifo_bank_register.bank[6][58] ;
 wire \fifo_bank_register.bank[6][59] ;
 wire \fifo_bank_register.bank[6][5] ;
 wire \fifo_bank_register.bank[6][60] ;
 wire \fifo_bank_register.bank[6][61] ;
 wire \fifo_bank_register.bank[6][62] ;
 wire \fifo_bank_register.bank[6][63] ;
 wire \fifo_bank_register.bank[6][64] ;
 wire \fifo_bank_register.bank[6][65] ;
 wire \fifo_bank_register.bank[6][66] ;
 wire \fifo_bank_register.bank[6][67] ;
 wire \fifo_bank_register.bank[6][68] ;
 wire \fifo_bank_register.bank[6][69] ;
 wire \fifo_bank_register.bank[6][6] ;
 wire \fifo_bank_register.bank[6][70] ;
 wire \fifo_bank_register.bank[6][71] ;
 wire \fifo_bank_register.bank[6][72] ;
 wire \fifo_bank_register.bank[6][73] ;
 wire \fifo_bank_register.bank[6][74] ;
 wire \fifo_bank_register.bank[6][75] ;
 wire \fifo_bank_register.bank[6][76] ;
 wire \fifo_bank_register.bank[6][77] ;
 wire \fifo_bank_register.bank[6][78] ;
 wire \fifo_bank_register.bank[6][79] ;
 wire \fifo_bank_register.bank[6][7] ;
 wire \fifo_bank_register.bank[6][80] ;
 wire \fifo_bank_register.bank[6][81] ;
 wire \fifo_bank_register.bank[6][82] ;
 wire \fifo_bank_register.bank[6][83] ;
 wire \fifo_bank_register.bank[6][84] ;
 wire \fifo_bank_register.bank[6][85] ;
 wire \fifo_bank_register.bank[6][86] ;
 wire \fifo_bank_register.bank[6][87] ;
 wire \fifo_bank_register.bank[6][88] ;
 wire \fifo_bank_register.bank[6][89] ;
 wire \fifo_bank_register.bank[6][8] ;
 wire \fifo_bank_register.bank[6][90] ;
 wire \fifo_bank_register.bank[6][91] ;
 wire \fifo_bank_register.bank[6][92] ;
 wire \fifo_bank_register.bank[6][93] ;
 wire \fifo_bank_register.bank[6][94] ;
 wire \fifo_bank_register.bank[6][95] ;
 wire \fifo_bank_register.bank[6][96] ;
 wire \fifo_bank_register.bank[6][97] ;
 wire \fifo_bank_register.bank[6][98] ;
 wire \fifo_bank_register.bank[6][99] ;
 wire \fifo_bank_register.bank[6][9] ;
 wire \fifo_bank_register.bank[7][0] ;
 wire \fifo_bank_register.bank[7][100] ;
 wire \fifo_bank_register.bank[7][101] ;
 wire \fifo_bank_register.bank[7][102] ;
 wire \fifo_bank_register.bank[7][103] ;
 wire \fifo_bank_register.bank[7][104] ;
 wire \fifo_bank_register.bank[7][105] ;
 wire \fifo_bank_register.bank[7][106] ;
 wire \fifo_bank_register.bank[7][107] ;
 wire \fifo_bank_register.bank[7][108] ;
 wire \fifo_bank_register.bank[7][109] ;
 wire \fifo_bank_register.bank[7][10] ;
 wire \fifo_bank_register.bank[7][110] ;
 wire \fifo_bank_register.bank[7][111] ;
 wire \fifo_bank_register.bank[7][112] ;
 wire \fifo_bank_register.bank[7][113] ;
 wire \fifo_bank_register.bank[7][114] ;
 wire \fifo_bank_register.bank[7][115] ;
 wire \fifo_bank_register.bank[7][116] ;
 wire \fifo_bank_register.bank[7][117] ;
 wire \fifo_bank_register.bank[7][118] ;
 wire \fifo_bank_register.bank[7][119] ;
 wire \fifo_bank_register.bank[7][11] ;
 wire \fifo_bank_register.bank[7][120] ;
 wire \fifo_bank_register.bank[7][121] ;
 wire \fifo_bank_register.bank[7][122] ;
 wire \fifo_bank_register.bank[7][123] ;
 wire \fifo_bank_register.bank[7][124] ;
 wire \fifo_bank_register.bank[7][125] ;
 wire \fifo_bank_register.bank[7][126] ;
 wire \fifo_bank_register.bank[7][127] ;
 wire \fifo_bank_register.bank[7][12] ;
 wire \fifo_bank_register.bank[7][13] ;
 wire \fifo_bank_register.bank[7][14] ;
 wire \fifo_bank_register.bank[7][15] ;
 wire \fifo_bank_register.bank[7][16] ;
 wire \fifo_bank_register.bank[7][17] ;
 wire \fifo_bank_register.bank[7][18] ;
 wire \fifo_bank_register.bank[7][19] ;
 wire \fifo_bank_register.bank[7][1] ;
 wire \fifo_bank_register.bank[7][20] ;
 wire \fifo_bank_register.bank[7][21] ;
 wire \fifo_bank_register.bank[7][22] ;
 wire \fifo_bank_register.bank[7][23] ;
 wire \fifo_bank_register.bank[7][24] ;
 wire \fifo_bank_register.bank[7][25] ;
 wire \fifo_bank_register.bank[7][26] ;
 wire \fifo_bank_register.bank[7][27] ;
 wire \fifo_bank_register.bank[7][28] ;
 wire \fifo_bank_register.bank[7][29] ;
 wire \fifo_bank_register.bank[7][2] ;
 wire \fifo_bank_register.bank[7][30] ;
 wire \fifo_bank_register.bank[7][31] ;
 wire \fifo_bank_register.bank[7][32] ;
 wire \fifo_bank_register.bank[7][33] ;
 wire \fifo_bank_register.bank[7][34] ;
 wire \fifo_bank_register.bank[7][35] ;
 wire \fifo_bank_register.bank[7][36] ;
 wire \fifo_bank_register.bank[7][37] ;
 wire \fifo_bank_register.bank[7][38] ;
 wire \fifo_bank_register.bank[7][39] ;
 wire \fifo_bank_register.bank[7][3] ;
 wire \fifo_bank_register.bank[7][40] ;
 wire \fifo_bank_register.bank[7][41] ;
 wire \fifo_bank_register.bank[7][42] ;
 wire \fifo_bank_register.bank[7][43] ;
 wire \fifo_bank_register.bank[7][44] ;
 wire \fifo_bank_register.bank[7][45] ;
 wire \fifo_bank_register.bank[7][46] ;
 wire \fifo_bank_register.bank[7][47] ;
 wire \fifo_bank_register.bank[7][48] ;
 wire \fifo_bank_register.bank[7][49] ;
 wire \fifo_bank_register.bank[7][4] ;
 wire \fifo_bank_register.bank[7][50] ;
 wire \fifo_bank_register.bank[7][51] ;
 wire \fifo_bank_register.bank[7][52] ;
 wire \fifo_bank_register.bank[7][53] ;
 wire \fifo_bank_register.bank[7][54] ;
 wire \fifo_bank_register.bank[7][55] ;
 wire \fifo_bank_register.bank[7][56] ;
 wire \fifo_bank_register.bank[7][57] ;
 wire \fifo_bank_register.bank[7][58] ;
 wire \fifo_bank_register.bank[7][59] ;
 wire \fifo_bank_register.bank[7][5] ;
 wire \fifo_bank_register.bank[7][60] ;
 wire \fifo_bank_register.bank[7][61] ;
 wire \fifo_bank_register.bank[7][62] ;
 wire \fifo_bank_register.bank[7][63] ;
 wire \fifo_bank_register.bank[7][64] ;
 wire \fifo_bank_register.bank[7][65] ;
 wire \fifo_bank_register.bank[7][66] ;
 wire \fifo_bank_register.bank[7][67] ;
 wire \fifo_bank_register.bank[7][68] ;
 wire \fifo_bank_register.bank[7][69] ;
 wire \fifo_bank_register.bank[7][6] ;
 wire \fifo_bank_register.bank[7][70] ;
 wire \fifo_bank_register.bank[7][71] ;
 wire \fifo_bank_register.bank[7][72] ;
 wire \fifo_bank_register.bank[7][73] ;
 wire \fifo_bank_register.bank[7][74] ;
 wire \fifo_bank_register.bank[7][75] ;
 wire \fifo_bank_register.bank[7][76] ;
 wire \fifo_bank_register.bank[7][77] ;
 wire \fifo_bank_register.bank[7][78] ;
 wire \fifo_bank_register.bank[7][79] ;
 wire \fifo_bank_register.bank[7][7] ;
 wire \fifo_bank_register.bank[7][80] ;
 wire \fifo_bank_register.bank[7][81] ;
 wire \fifo_bank_register.bank[7][82] ;
 wire \fifo_bank_register.bank[7][83] ;
 wire \fifo_bank_register.bank[7][84] ;
 wire \fifo_bank_register.bank[7][85] ;
 wire \fifo_bank_register.bank[7][86] ;
 wire \fifo_bank_register.bank[7][87] ;
 wire \fifo_bank_register.bank[7][88] ;
 wire \fifo_bank_register.bank[7][89] ;
 wire \fifo_bank_register.bank[7][8] ;
 wire \fifo_bank_register.bank[7][90] ;
 wire \fifo_bank_register.bank[7][91] ;
 wire \fifo_bank_register.bank[7][92] ;
 wire \fifo_bank_register.bank[7][93] ;
 wire \fifo_bank_register.bank[7][94] ;
 wire \fifo_bank_register.bank[7][95] ;
 wire \fifo_bank_register.bank[7][96] ;
 wire \fifo_bank_register.bank[7][97] ;
 wire \fifo_bank_register.bank[7][98] ;
 wire \fifo_bank_register.bank[7][99] ;
 wire \fifo_bank_register.bank[7][9] ;
 wire \fifo_bank_register.bank[8][0] ;
 wire \fifo_bank_register.bank[8][100] ;
 wire \fifo_bank_register.bank[8][101] ;
 wire \fifo_bank_register.bank[8][102] ;
 wire \fifo_bank_register.bank[8][103] ;
 wire \fifo_bank_register.bank[8][104] ;
 wire \fifo_bank_register.bank[8][105] ;
 wire \fifo_bank_register.bank[8][106] ;
 wire \fifo_bank_register.bank[8][107] ;
 wire \fifo_bank_register.bank[8][108] ;
 wire \fifo_bank_register.bank[8][109] ;
 wire \fifo_bank_register.bank[8][10] ;
 wire \fifo_bank_register.bank[8][110] ;
 wire \fifo_bank_register.bank[8][111] ;
 wire \fifo_bank_register.bank[8][112] ;
 wire \fifo_bank_register.bank[8][113] ;
 wire \fifo_bank_register.bank[8][114] ;
 wire \fifo_bank_register.bank[8][115] ;
 wire \fifo_bank_register.bank[8][116] ;
 wire \fifo_bank_register.bank[8][117] ;
 wire \fifo_bank_register.bank[8][118] ;
 wire \fifo_bank_register.bank[8][119] ;
 wire \fifo_bank_register.bank[8][11] ;
 wire \fifo_bank_register.bank[8][120] ;
 wire \fifo_bank_register.bank[8][121] ;
 wire \fifo_bank_register.bank[8][122] ;
 wire \fifo_bank_register.bank[8][123] ;
 wire \fifo_bank_register.bank[8][124] ;
 wire \fifo_bank_register.bank[8][125] ;
 wire \fifo_bank_register.bank[8][126] ;
 wire \fifo_bank_register.bank[8][127] ;
 wire \fifo_bank_register.bank[8][12] ;
 wire \fifo_bank_register.bank[8][13] ;
 wire \fifo_bank_register.bank[8][14] ;
 wire \fifo_bank_register.bank[8][15] ;
 wire \fifo_bank_register.bank[8][16] ;
 wire \fifo_bank_register.bank[8][17] ;
 wire \fifo_bank_register.bank[8][18] ;
 wire \fifo_bank_register.bank[8][19] ;
 wire \fifo_bank_register.bank[8][1] ;
 wire \fifo_bank_register.bank[8][20] ;
 wire \fifo_bank_register.bank[8][21] ;
 wire \fifo_bank_register.bank[8][22] ;
 wire \fifo_bank_register.bank[8][23] ;
 wire \fifo_bank_register.bank[8][24] ;
 wire \fifo_bank_register.bank[8][25] ;
 wire \fifo_bank_register.bank[8][26] ;
 wire \fifo_bank_register.bank[8][27] ;
 wire \fifo_bank_register.bank[8][28] ;
 wire \fifo_bank_register.bank[8][29] ;
 wire \fifo_bank_register.bank[8][2] ;
 wire \fifo_bank_register.bank[8][30] ;
 wire \fifo_bank_register.bank[8][31] ;
 wire \fifo_bank_register.bank[8][32] ;
 wire \fifo_bank_register.bank[8][33] ;
 wire \fifo_bank_register.bank[8][34] ;
 wire \fifo_bank_register.bank[8][35] ;
 wire \fifo_bank_register.bank[8][36] ;
 wire \fifo_bank_register.bank[8][37] ;
 wire \fifo_bank_register.bank[8][38] ;
 wire \fifo_bank_register.bank[8][39] ;
 wire \fifo_bank_register.bank[8][3] ;
 wire \fifo_bank_register.bank[8][40] ;
 wire \fifo_bank_register.bank[8][41] ;
 wire \fifo_bank_register.bank[8][42] ;
 wire \fifo_bank_register.bank[8][43] ;
 wire \fifo_bank_register.bank[8][44] ;
 wire \fifo_bank_register.bank[8][45] ;
 wire \fifo_bank_register.bank[8][46] ;
 wire \fifo_bank_register.bank[8][47] ;
 wire \fifo_bank_register.bank[8][48] ;
 wire \fifo_bank_register.bank[8][49] ;
 wire \fifo_bank_register.bank[8][4] ;
 wire \fifo_bank_register.bank[8][50] ;
 wire \fifo_bank_register.bank[8][51] ;
 wire \fifo_bank_register.bank[8][52] ;
 wire \fifo_bank_register.bank[8][53] ;
 wire \fifo_bank_register.bank[8][54] ;
 wire \fifo_bank_register.bank[8][55] ;
 wire \fifo_bank_register.bank[8][56] ;
 wire \fifo_bank_register.bank[8][57] ;
 wire \fifo_bank_register.bank[8][58] ;
 wire \fifo_bank_register.bank[8][59] ;
 wire \fifo_bank_register.bank[8][5] ;
 wire \fifo_bank_register.bank[8][60] ;
 wire \fifo_bank_register.bank[8][61] ;
 wire \fifo_bank_register.bank[8][62] ;
 wire \fifo_bank_register.bank[8][63] ;
 wire \fifo_bank_register.bank[8][64] ;
 wire \fifo_bank_register.bank[8][65] ;
 wire \fifo_bank_register.bank[8][66] ;
 wire \fifo_bank_register.bank[8][67] ;
 wire \fifo_bank_register.bank[8][68] ;
 wire \fifo_bank_register.bank[8][69] ;
 wire \fifo_bank_register.bank[8][6] ;
 wire \fifo_bank_register.bank[8][70] ;
 wire \fifo_bank_register.bank[8][71] ;
 wire \fifo_bank_register.bank[8][72] ;
 wire \fifo_bank_register.bank[8][73] ;
 wire \fifo_bank_register.bank[8][74] ;
 wire \fifo_bank_register.bank[8][75] ;
 wire \fifo_bank_register.bank[8][76] ;
 wire \fifo_bank_register.bank[8][77] ;
 wire \fifo_bank_register.bank[8][78] ;
 wire \fifo_bank_register.bank[8][79] ;
 wire \fifo_bank_register.bank[8][7] ;
 wire \fifo_bank_register.bank[8][80] ;
 wire \fifo_bank_register.bank[8][81] ;
 wire \fifo_bank_register.bank[8][82] ;
 wire \fifo_bank_register.bank[8][83] ;
 wire \fifo_bank_register.bank[8][84] ;
 wire \fifo_bank_register.bank[8][85] ;
 wire \fifo_bank_register.bank[8][86] ;
 wire \fifo_bank_register.bank[8][87] ;
 wire \fifo_bank_register.bank[8][88] ;
 wire \fifo_bank_register.bank[8][89] ;
 wire \fifo_bank_register.bank[8][8] ;
 wire \fifo_bank_register.bank[8][90] ;
 wire \fifo_bank_register.bank[8][91] ;
 wire \fifo_bank_register.bank[8][92] ;
 wire \fifo_bank_register.bank[8][93] ;
 wire \fifo_bank_register.bank[8][94] ;
 wire \fifo_bank_register.bank[8][95] ;
 wire \fifo_bank_register.bank[8][96] ;
 wire \fifo_bank_register.bank[8][97] ;
 wire \fifo_bank_register.bank[8][98] ;
 wire \fifo_bank_register.bank[8][99] ;
 wire \fifo_bank_register.bank[8][9] ;
 wire \fifo_bank_register.bank[9][0] ;
 wire \fifo_bank_register.bank[9][100] ;
 wire \fifo_bank_register.bank[9][101] ;
 wire \fifo_bank_register.bank[9][102] ;
 wire \fifo_bank_register.bank[9][103] ;
 wire \fifo_bank_register.bank[9][104] ;
 wire \fifo_bank_register.bank[9][105] ;
 wire \fifo_bank_register.bank[9][106] ;
 wire \fifo_bank_register.bank[9][107] ;
 wire \fifo_bank_register.bank[9][108] ;
 wire \fifo_bank_register.bank[9][109] ;
 wire \fifo_bank_register.bank[9][10] ;
 wire \fifo_bank_register.bank[9][110] ;
 wire \fifo_bank_register.bank[9][111] ;
 wire \fifo_bank_register.bank[9][112] ;
 wire \fifo_bank_register.bank[9][113] ;
 wire \fifo_bank_register.bank[9][114] ;
 wire \fifo_bank_register.bank[9][115] ;
 wire \fifo_bank_register.bank[9][116] ;
 wire \fifo_bank_register.bank[9][117] ;
 wire \fifo_bank_register.bank[9][118] ;
 wire \fifo_bank_register.bank[9][119] ;
 wire \fifo_bank_register.bank[9][11] ;
 wire \fifo_bank_register.bank[9][120] ;
 wire \fifo_bank_register.bank[9][121] ;
 wire \fifo_bank_register.bank[9][122] ;
 wire \fifo_bank_register.bank[9][123] ;
 wire \fifo_bank_register.bank[9][124] ;
 wire \fifo_bank_register.bank[9][125] ;
 wire \fifo_bank_register.bank[9][126] ;
 wire \fifo_bank_register.bank[9][127] ;
 wire \fifo_bank_register.bank[9][12] ;
 wire \fifo_bank_register.bank[9][13] ;
 wire \fifo_bank_register.bank[9][14] ;
 wire \fifo_bank_register.bank[9][15] ;
 wire \fifo_bank_register.bank[9][16] ;
 wire \fifo_bank_register.bank[9][17] ;
 wire \fifo_bank_register.bank[9][18] ;
 wire \fifo_bank_register.bank[9][19] ;
 wire \fifo_bank_register.bank[9][1] ;
 wire \fifo_bank_register.bank[9][20] ;
 wire \fifo_bank_register.bank[9][21] ;
 wire \fifo_bank_register.bank[9][22] ;
 wire \fifo_bank_register.bank[9][23] ;
 wire \fifo_bank_register.bank[9][24] ;
 wire \fifo_bank_register.bank[9][25] ;
 wire \fifo_bank_register.bank[9][26] ;
 wire \fifo_bank_register.bank[9][27] ;
 wire \fifo_bank_register.bank[9][28] ;
 wire \fifo_bank_register.bank[9][29] ;
 wire \fifo_bank_register.bank[9][2] ;
 wire \fifo_bank_register.bank[9][30] ;
 wire \fifo_bank_register.bank[9][31] ;
 wire \fifo_bank_register.bank[9][32] ;
 wire \fifo_bank_register.bank[9][33] ;
 wire \fifo_bank_register.bank[9][34] ;
 wire \fifo_bank_register.bank[9][35] ;
 wire \fifo_bank_register.bank[9][36] ;
 wire \fifo_bank_register.bank[9][37] ;
 wire \fifo_bank_register.bank[9][38] ;
 wire \fifo_bank_register.bank[9][39] ;
 wire \fifo_bank_register.bank[9][3] ;
 wire \fifo_bank_register.bank[9][40] ;
 wire \fifo_bank_register.bank[9][41] ;
 wire \fifo_bank_register.bank[9][42] ;
 wire \fifo_bank_register.bank[9][43] ;
 wire \fifo_bank_register.bank[9][44] ;
 wire \fifo_bank_register.bank[9][45] ;
 wire \fifo_bank_register.bank[9][46] ;
 wire \fifo_bank_register.bank[9][47] ;
 wire \fifo_bank_register.bank[9][48] ;
 wire \fifo_bank_register.bank[9][49] ;
 wire \fifo_bank_register.bank[9][4] ;
 wire \fifo_bank_register.bank[9][50] ;
 wire \fifo_bank_register.bank[9][51] ;
 wire \fifo_bank_register.bank[9][52] ;
 wire \fifo_bank_register.bank[9][53] ;
 wire \fifo_bank_register.bank[9][54] ;
 wire \fifo_bank_register.bank[9][55] ;
 wire \fifo_bank_register.bank[9][56] ;
 wire \fifo_bank_register.bank[9][57] ;
 wire \fifo_bank_register.bank[9][58] ;
 wire \fifo_bank_register.bank[9][59] ;
 wire \fifo_bank_register.bank[9][5] ;
 wire \fifo_bank_register.bank[9][60] ;
 wire \fifo_bank_register.bank[9][61] ;
 wire \fifo_bank_register.bank[9][62] ;
 wire \fifo_bank_register.bank[9][63] ;
 wire \fifo_bank_register.bank[9][64] ;
 wire \fifo_bank_register.bank[9][65] ;
 wire \fifo_bank_register.bank[9][66] ;
 wire \fifo_bank_register.bank[9][67] ;
 wire \fifo_bank_register.bank[9][68] ;
 wire \fifo_bank_register.bank[9][69] ;
 wire \fifo_bank_register.bank[9][6] ;
 wire \fifo_bank_register.bank[9][70] ;
 wire \fifo_bank_register.bank[9][71] ;
 wire \fifo_bank_register.bank[9][72] ;
 wire \fifo_bank_register.bank[9][73] ;
 wire \fifo_bank_register.bank[9][74] ;
 wire \fifo_bank_register.bank[9][75] ;
 wire \fifo_bank_register.bank[9][76] ;
 wire \fifo_bank_register.bank[9][77] ;
 wire \fifo_bank_register.bank[9][78] ;
 wire \fifo_bank_register.bank[9][79] ;
 wire \fifo_bank_register.bank[9][7] ;
 wire \fifo_bank_register.bank[9][80] ;
 wire \fifo_bank_register.bank[9][81] ;
 wire \fifo_bank_register.bank[9][82] ;
 wire \fifo_bank_register.bank[9][83] ;
 wire \fifo_bank_register.bank[9][84] ;
 wire \fifo_bank_register.bank[9][85] ;
 wire \fifo_bank_register.bank[9][86] ;
 wire \fifo_bank_register.bank[9][87] ;
 wire \fifo_bank_register.bank[9][88] ;
 wire \fifo_bank_register.bank[9][89] ;
 wire \fifo_bank_register.bank[9][8] ;
 wire \fifo_bank_register.bank[9][90] ;
 wire \fifo_bank_register.bank[9][91] ;
 wire \fifo_bank_register.bank[9][92] ;
 wire \fifo_bank_register.bank[9][93] ;
 wire \fifo_bank_register.bank[9][94] ;
 wire \fifo_bank_register.bank[9][95] ;
 wire \fifo_bank_register.bank[9][96] ;
 wire \fifo_bank_register.bank[9][97] ;
 wire \fifo_bank_register.bank[9][98] ;
 wire \fifo_bank_register.bank[9][99] ;
 wire \fifo_bank_register.bank[9][9] ;
 wire \fifo_bank_register.clk ;
 wire \fifo_bank_register.data_out[0] ;
 wire \fifo_bank_register.data_out[100] ;
 wire \fifo_bank_register.data_out[101] ;
 wire \fifo_bank_register.data_out[102] ;
 wire \fifo_bank_register.data_out[103] ;
 wire \fifo_bank_register.data_out[104] ;
 wire \fifo_bank_register.data_out[105] ;
 wire \fifo_bank_register.data_out[106] ;
 wire \fifo_bank_register.data_out[107] ;
 wire \fifo_bank_register.data_out[108] ;
 wire \fifo_bank_register.data_out[109] ;
 wire \fifo_bank_register.data_out[10] ;
 wire \fifo_bank_register.data_out[110] ;
 wire \fifo_bank_register.data_out[111] ;
 wire \fifo_bank_register.data_out[112] ;
 wire \fifo_bank_register.data_out[113] ;
 wire \fifo_bank_register.data_out[114] ;
 wire \fifo_bank_register.data_out[115] ;
 wire \fifo_bank_register.data_out[116] ;
 wire \fifo_bank_register.data_out[117] ;
 wire \fifo_bank_register.data_out[118] ;
 wire \fifo_bank_register.data_out[119] ;
 wire \fifo_bank_register.data_out[11] ;
 wire \fifo_bank_register.data_out[120] ;
 wire \fifo_bank_register.data_out[121] ;
 wire \fifo_bank_register.data_out[122] ;
 wire \fifo_bank_register.data_out[123] ;
 wire \fifo_bank_register.data_out[124] ;
 wire \fifo_bank_register.data_out[125] ;
 wire \fifo_bank_register.data_out[126] ;
 wire \fifo_bank_register.data_out[127] ;
 wire \fifo_bank_register.data_out[12] ;
 wire \fifo_bank_register.data_out[13] ;
 wire \fifo_bank_register.data_out[14] ;
 wire \fifo_bank_register.data_out[15] ;
 wire \fifo_bank_register.data_out[16] ;
 wire \fifo_bank_register.data_out[17] ;
 wire \fifo_bank_register.data_out[18] ;
 wire \fifo_bank_register.data_out[19] ;
 wire \fifo_bank_register.data_out[1] ;
 wire \fifo_bank_register.data_out[20] ;
 wire \fifo_bank_register.data_out[21] ;
 wire \fifo_bank_register.data_out[22] ;
 wire \fifo_bank_register.data_out[23] ;
 wire \fifo_bank_register.data_out[24] ;
 wire \fifo_bank_register.data_out[25] ;
 wire \fifo_bank_register.data_out[26] ;
 wire \fifo_bank_register.data_out[27] ;
 wire \fifo_bank_register.data_out[28] ;
 wire \fifo_bank_register.data_out[29] ;
 wire \fifo_bank_register.data_out[2] ;
 wire \fifo_bank_register.data_out[30] ;
 wire \fifo_bank_register.data_out[31] ;
 wire \fifo_bank_register.data_out[32] ;
 wire \fifo_bank_register.data_out[33] ;
 wire \fifo_bank_register.data_out[34] ;
 wire \fifo_bank_register.data_out[35] ;
 wire \fifo_bank_register.data_out[36] ;
 wire \fifo_bank_register.data_out[37] ;
 wire \fifo_bank_register.data_out[38] ;
 wire \fifo_bank_register.data_out[39] ;
 wire \fifo_bank_register.data_out[3] ;
 wire \fifo_bank_register.data_out[40] ;
 wire \fifo_bank_register.data_out[41] ;
 wire \fifo_bank_register.data_out[42] ;
 wire \fifo_bank_register.data_out[43] ;
 wire \fifo_bank_register.data_out[44] ;
 wire \fifo_bank_register.data_out[45] ;
 wire \fifo_bank_register.data_out[46] ;
 wire \fifo_bank_register.data_out[47] ;
 wire \fifo_bank_register.data_out[48] ;
 wire \fifo_bank_register.data_out[49] ;
 wire \fifo_bank_register.data_out[4] ;
 wire \fifo_bank_register.data_out[50] ;
 wire \fifo_bank_register.data_out[51] ;
 wire \fifo_bank_register.data_out[52] ;
 wire \fifo_bank_register.data_out[53] ;
 wire \fifo_bank_register.data_out[54] ;
 wire \fifo_bank_register.data_out[55] ;
 wire \fifo_bank_register.data_out[56] ;
 wire \fifo_bank_register.data_out[57] ;
 wire \fifo_bank_register.data_out[58] ;
 wire \fifo_bank_register.data_out[59] ;
 wire \fifo_bank_register.data_out[5] ;
 wire \fifo_bank_register.data_out[60] ;
 wire \fifo_bank_register.data_out[61] ;
 wire \fifo_bank_register.data_out[62] ;
 wire \fifo_bank_register.data_out[63] ;
 wire \fifo_bank_register.data_out[64] ;
 wire \fifo_bank_register.data_out[65] ;
 wire \fifo_bank_register.data_out[66] ;
 wire \fifo_bank_register.data_out[67] ;
 wire \fifo_bank_register.data_out[68] ;
 wire \fifo_bank_register.data_out[69] ;
 wire \fifo_bank_register.data_out[6] ;
 wire \fifo_bank_register.data_out[70] ;
 wire \fifo_bank_register.data_out[71] ;
 wire \fifo_bank_register.data_out[72] ;
 wire \fifo_bank_register.data_out[73] ;
 wire \fifo_bank_register.data_out[74] ;
 wire \fifo_bank_register.data_out[75] ;
 wire \fifo_bank_register.data_out[76] ;
 wire \fifo_bank_register.data_out[77] ;
 wire \fifo_bank_register.data_out[78] ;
 wire \fifo_bank_register.data_out[79] ;
 wire \fifo_bank_register.data_out[7] ;
 wire \fifo_bank_register.data_out[80] ;
 wire \fifo_bank_register.data_out[81] ;
 wire \fifo_bank_register.data_out[82] ;
 wire \fifo_bank_register.data_out[83] ;
 wire \fifo_bank_register.data_out[84] ;
 wire \fifo_bank_register.data_out[85] ;
 wire \fifo_bank_register.data_out[86] ;
 wire \fifo_bank_register.data_out[87] ;
 wire \fifo_bank_register.data_out[88] ;
 wire \fifo_bank_register.data_out[89] ;
 wire \fifo_bank_register.data_out[8] ;
 wire \fifo_bank_register.data_out[90] ;
 wire \fifo_bank_register.data_out[91] ;
 wire \fifo_bank_register.data_out[92] ;
 wire \fifo_bank_register.data_out[93] ;
 wire \fifo_bank_register.data_out[94] ;
 wire \fifo_bank_register.data_out[95] ;
 wire \fifo_bank_register.data_out[96] ;
 wire \fifo_bank_register.data_out[97] ;
 wire \fifo_bank_register.data_out[98] ;
 wire \fifo_bank_register.data_out[99] ;
 wire \fifo_bank_register.data_out[9] ;
 wire \fifo_bank_register.read_ptr[0] ;
 wire \fifo_bank_register.read_ptr[1] ;
 wire \fifo_bank_register.read_ptr[2] ;
 wire \fifo_bank_register.read_ptr[3] ;
 wire \fifo_bank_register.write_ptr[0] ;
 wire \fifo_bank_register.write_ptr[1] ;
 wire \fifo_bank_register.write_ptr[2] ;
 wire \fifo_bank_register.write_ptr[3] ;
 wire first_round_reg;
 wire \ks1.col[0] ;
 wire \ks1.col[16] ;
 wire \ks1.col[17] ;
 wire \ks1.col[18] ;
 wire \ks1.col[19] ;
 wire \ks1.col[1] ;
 wire \ks1.col[20] ;
 wire \ks1.col[21] ;
 wire \ks1.col[22] ;
 wire \ks1.col[23] ;
 wire \ks1.col[24] ;
 wire \ks1.col[25] ;
 wire \ks1.col[26] ;
 wire \ks1.col[27] ;
 wire \ks1.col[28] ;
 wire \ks1.col[29] ;
 wire \ks1.col[2] ;
 wire \ks1.col[30] ;
 wire \ks1.col[31] ;
 wire \ks1.col[3] ;
 wire \ks1.col[4] ;
 wire \ks1.col[5] ;
 wire \ks1.col[6] ;
 wire \ks1.col[7] ;
 wire \ks1.key_reg[0] ;
 wire \ks1.key_reg[100] ;
 wire \ks1.key_reg[101] ;
 wire \ks1.key_reg[102] ;
 wire \ks1.key_reg[103] ;
 wire \ks1.key_reg[104] ;
 wire \ks1.key_reg[105] ;
 wire \ks1.key_reg[106] ;
 wire \ks1.key_reg[107] ;
 wire \ks1.key_reg[108] ;
 wire \ks1.key_reg[109] ;
 wire \ks1.key_reg[10] ;
 wire \ks1.key_reg[110] ;
 wire \ks1.key_reg[111] ;
 wire \ks1.key_reg[112] ;
 wire \ks1.key_reg[113] ;
 wire \ks1.key_reg[114] ;
 wire \ks1.key_reg[115] ;
 wire \ks1.key_reg[116] ;
 wire \ks1.key_reg[117] ;
 wire \ks1.key_reg[118] ;
 wire \ks1.key_reg[119] ;
 wire \ks1.key_reg[11] ;
 wire \ks1.key_reg[120] ;
 wire \ks1.key_reg[121] ;
 wire \ks1.key_reg[122] ;
 wire \ks1.key_reg[123] ;
 wire \ks1.key_reg[124] ;
 wire \ks1.key_reg[125] ;
 wire \ks1.key_reg[126] ;
 wire \ks1.key_reg[127] ;
 wire \ks1.key_reg[12] ;
 wire \ks1.key_reg[13] ;
 wire \ks1.key_reg[14] ;
 wire \ks1.key_reg[15] ;
 wire \ks1.key_reg[16] ;
 wire \ks1.key_reg[17] ;
 wire \ks1.key_reg[18] ;
 wire \ks1.key_reg[19] ;
 wire \ks1.key_reg[1] ;
 wire \ks1.key_reg[20] ;
 wire \ks1.key_reg[21] ;
 wire \ks1.key_reg[22] ;
 wire \ks1.key_reg[23] ;
 wire \ks1.key_reg[24] ;
 wire \ks1.key_reg[25] ;
 wire \ks1.key_reg[26] ;
 wire \ks1.key_reg[27] ;
 wire \ks1.key_reg[28] ;
 wire \ks1.key_reg[29] ;
 wire \ks1.key_reg[2] ;
 wire \ks1.key_reg[30] ;
 wire \ks1.key_reg[31] ;
 wire \ks1.key_reg[32] ;
 wire \ks1.key_reg[33] ;
 wire \ks1.key_reg[34] ;
 wire \ks1.key_reg[35] ;
 wire \ks1.key_reg[36] ;
 wire \ks1.key_reg[37] ;
 wire \ks1.key_reg[38] ;
 wire \ks1.key_reg[39] ;
 wire \ks1.key_reg[3] ;
 wire \ks1.key_reg[40] ;
 wire \ks1.key_reg[41] ;
 wire \ks1.key_reg[42] ;
 wire \ks1.key_reg[43] ;
 wire \ks1.key_reg[44] ;
 wire \ks1.key_reg[45] ;
 wire \ks1.key_reg[46] ;
 wire \ks1.key_reg[47] ;
 wire \ks1.key_reg[48] ;
 wire \ks1.key_reg[49] ;
 wire \ks1.key_reg[4] ;
 wire \ks1.key_reg[50] ;
 wire \ks1.key_reg[51] ;
 wire \ks1.key_reg[52] ;
 wire \ks1.key_reg[53] ;
 wire \ks1.key_reg[54] ;
 wire \ks1.key_reg[55] ;
 wire \ks1.key_reg[56] ;
 wire \ks1.key_reg[57] ;
 wire \ks1.key_reg[58] ;
 wire \ks1.key_reg[59] ;
 wire \ks1.key_reg[5] ;
 wire \ks1.key_reg[60] ;
 wire \ks1.key_reg[61] ;
 wire \ks1.key_reg[62] ;
 wire \ks1.key_reg[63] ;
 wire \ks1.key_reg[64] ;
 wire \ks1.key_reg[65] ;
 wire \ks1.key_reg[66] ;
 wire \ks1.key_reg[67] ;
 wire \ks1.key_reg[68] ;
 wire \ks1.key_reg[69] ;
 wire \ks1.key_reg[6] ;
 wire \ks1.key_reg[70] ;
 wire \ks1.key_reg[71] ;
 wire \ks1.key_reg[72] ;
 wire \ks1.key_reg[73] ;
 wire \ks1.key_reg[74] ;
 wire \ks1.key_reg[75] ;
 wire \ks1.key_reg[76] ;
 wire \ks1.key_reg[77] ;
 wire \ks1.key_reg[78] ;
 wire \ks1.key_reg[79] ;
 wire \ks1.key_reg[7] ;
 wire \ks1.key_reg[80] ;
 wire \ks1.key_reg[81] ;
 wire \ks1.key_reg[82] ;
 wire \ks1.key_reg[83] ;
 wire \ks1.key_reg[84] ;
 wire \ks1.key_reg[85] ;
 wire \ks1.key_reg[86] ;
 wire \ks1.key_reg[87] ;
 wire \ks1.key_reg[88] ;
 wire \ks1.key_reg[89] ;
 wire \ks1.key_reg[8] ;
 wire \ks1.key_reg[90] ;
 wire \ks1.key_reg[91] ;
 wire \ks1.key_reg[92] ;
 wire \ks1.key_reg[93] ;
 wire \ks1.key_reg[94] ;
 wire \ks1.key_reg[95] ;
 wire \ks1.key_reg[96] ;
 wire \ks1.key_reg[97] ;
 wire \ks1.key_reg[98] ;
 wire \ks1.key_reg[99] ;
 wire \ks1.key_reg[9] ;
 wire \ks1.next_ready_o ;
 wire \ks1.ready_o ;
 wire \ks1.state[0] ;
 wire \ks1.state[1] ;
 wire \ks1.state[2] ;
 wire \mix1.data_o[0] ;
 wire \mix1.data_o[100] ;
 wire \mix1.data_o[101] ;
 wire \mix1.data_o[102] ;
 wire \mix1.data_o[103] ;
 wire \mix1.data_o[104] ;
 wire \mix1.data_o[105] ;
 wire \mix1.data_o[106] ;
 wire \mix1.data_o[107] ;
 wire \mix1.data_o[108] ;
 wire \mix1.data_o[109] ;
 wire \mix1.data_o[10] ;
 wire \mix1.data_o[110] ;
 wire \mix1.data_o[111] ;
 wire \mix1.data_o[112] ;
 wire \mix1.data_o[113] ;
 wire \mix1.data_o[114] ;
 wire \mix1.data_o[115] ;
 wire \mix1.data_o[116] ;
 wire \mix1.data_o[117] ;
 wire \mix1.data_o[118] ;
 wire \mix1.data_o[119] ;
 wire \mix1.data_o[11] ;
 wire \mix1.data_o[120] ;
 wire \mix1.data_o[121] ;
 wire \mix1.data_o[122] ;
 wire \mix1.data_o[123] ;
 wire \mix1.data_o[124] ;
 wire \mix1.data_o[125] ;
 wire \mix1.data_o[126] ;
 wire \mix1.data_o[127] ;
 wire \mix1.data_o[12] ;
 wire \mix1.data_o[13] ;
 wire \mix1.data_o[14] ;
 wire \mix1.data_o[15] ;
 wire \mix1.data_o[16] ;
 wire \mix1.data_o[17] ;
 wire \mix1.data_o[18] ;
 wire \mix1.data_o[19] ;
 wire \mix1.data_o[1] ;
 wire \mix1.data_o[20] ;
 wire \mix1.data_o[21] ;
 wire \mix1.data_o[22] ;
 wire \mix1.data_o[23] ;
 wire \mix1.data_o[24] ;
 wire \mix1.data_o[25] ;
 wire \mix1.data_o[26] ;
 wire \mix1.data_o[27] ;
 wire \mix1.data_o[28] ;
 wire \mix1.data_o[29] ;
 wire \mix1.data_o[2] ;
 wire \mix1.data_o[30] ;
 wire \mix1.data_o[31] ;
 wire \mix1.data_o[32] ;
 wire \mix1.data_o[33] ;
 wire \mix1.data_o[34] ;
 wire \mix1.data_o[35] ;
 wire \mix1.data_o[36] ;
 wire \mix1.data_o[37] ;
 wire \mix1.data_o[38] ;
 wire \mix1.data_o[39] ;
 wire \mix1.data_o[3] ;
 wire \mix1.data_o[40] ;
 wire \mix1.data_o[41] ;
 wire \mix1.data_o[42] ;
 wire \mix1.data_o[43] ;
 wire \mix1.data_o[44] ;
 wire \mix1.data_o[45] ;
 wire \mix1.data_o[46] ;
 wire \mix1.data_o[47] ;
 wire \mix1.data_o[48] ;
 wire \mix1.data_o[49] ;
 wire \mix1.data_o[4] ;
 wire \mix1.data_o[50] ;
 wire \mix1.data_o[51] ;
 wire \mix1.data_o[52] ;
 wire \mix1.data_o[53] ;
 wire \mix1.data_o[54] ;
 wire \mix1.data_o[55] ;
 wire \mix1.data_o[56] ;
 wire \mix1.data_o[57] ;
 wire \mix1.data_o[58] ;
 wire \mix1.data_o[59] ;
 wire \mix1.data_o[5] ;
 wire \mix1.data_o[60] ;
 wire \mix1.data_o[61] ;
 wire \mix1.data_o[62] ;
 wire \mix1.data_o[63] ;
 wire \mix1.data_o[64] ;
 wire \mix1.data_o[65] ;
 wire \mix1.data_o[66] ;
 wire \mix1.data_o[67] ;
 wire \mix1.data_o[68] ;
 wire \mix1.data_o[69] ;
 wire \mix1.data_o[6] ;
 wire \mix1.data_o[70] ;
 wire \mix1.data_o[71] ;
 wire \mix1.data_o[72] ;
 wire \mix1.data_o[73] ;
 wire \mix1.data_o[74] ;
 wire \mix1.data_o[75] ;
 wire \mix1.data_o[76] ;
 wire \mix1.data_o[77] ;
 wire \mix1.data_o[78] ;
 wire \mix1.data_o[79] ;
 wire \mix1.data_o[7] ;
 wire \mix1.data_o[80] ;
 wire \mix1.data_o[81] ;
 wire \mix1.data_o[82] ;
 wire \mix1.data_o[83] ;
 wire \mix1.data_o[84] ;
 wire \mix1.data_o[85] ;
 wire \mix1.data_o[86] ;
 wire \mix1.data_o[87] ;
 wire \mix1.data_o[88] ;
 wire \mix1.data_o[89] ;
 wire \mix1.data_o[8] ;
 wire \mix1.data_o[90] ;
 wire \mix1.data_o[91] ;
 wire \mix1.data_o[92] ;
 wire \mix1.data_o[93] ;
 wire \mix1.data_o[94] ;
 wire \mix1.data_o[95] ;
 wire \mix1.data_o[96] ;
 wire \mix1.data_o[97] ;
 wire \mix1.data_o[98] ;
 wire \mix1.data_o[99] ;
 wire \mix1.data_o[9] ;
 wire \mix1.data_reg[100] ;
 wire \mix1.data_reg[101] ;
 wire \mix1.data_reg[102] ;
 wire \mix1.data_reg[103] ;
 wire \mix1.data_reg[104] ;
 wire \mix1.data_reg[105] ;
 wire \mix1.data_reg[106] ;
 wire \mix1.data_reg[107] ;
 wire \mix1.data_reg[108] ;
 wire \mix1.data_reg[109] ;
 wire \mix1.data_reg[110] ;
 wire \mix1.data_reg[111] ;
 wire \mix1.data_reg[112] ;
 wire \mix1.data_reg[113] ;
 wire \mix1.data_reg[114] ;
 wire \mix1.data_reg[115] ;
 wire \mix1.data_reg[116] ;
 wire \mix1.data_reg[117] ;
 wire \mix1.data_reg[118] ;
 wire \mix1.data_reg[119] ;
 wire \mix1.data_reg[120] ;
 wire \mix1.data_reg[121] ;
 wire \mix1.data_reg[122] ;
 wire \mix1.data_reg[123] ;
 wire \mix1.data_reg[124] ;
 wire \mix1.data_reg[125] ;
 wire \mix1.data_reg[126] ;
 wire \mix1.data_reg[127] ;
 wire \mix1.data_reg[32] ;
 wire \mix1.data_reg[33] ;
 wire \mix1.data_reg[34] ;
 wire \mix1.data_reg[35] ;
 wire \mix1.data_reg[36] ;
 wire \mix1.data_reg[37] ;
 wire \mix1.data_reg[38] ;
 wire \mix1.data_reg[39] ;
 wire \mix1.data_reg[40] ;
 wire \mix1.data_reg[41] ;
 wire \mix1.data_reg[42] ;
 wire \mix1.data_reg[43] ;
 wire \mix1.data_reg[44] ;
 wire \mix1.data_reg[45] ;
 wire \mix1.data_reg[46] ;
 wire \mix1.data_reg[47] ;
 wire \mix1.data_reg[48] ;
 wire \mix1.data_reg[49] ;
 wire \mix1.data_reg[50] ;
 wire \mix1.data_reg[51] ;
 wire \mix1.data_reg[52] ;
 wire \mix1.data_reg[53] ;
 wire \mix1.data_reg[54] ;
 wire \mix1.data_reg[55] ;
 wire \mix1.data_reg[56] ;
 wire \mix1.data_reg[57] ;
 wire \mix1.data_reg[58] ;
 wire \mix1.data_reg[59] ;
 wire \mix1.data_reg[60] ;
 wire \mix1.data_reg[61] ;
 wire \mix1.data_reg[62] ;
 wire \mix1.data_reg[63] ;
 wire \mix1.data_reg[64] ;
 wire \mix1.data_reg[65] ;
 wire \mix1.data_reg[66] ;
 wire \mix1.data_reg[67] ;
 wire \mix1.data_reg[68] ;
 wire \mix1.data_reg[69] ;
 wire \mix1.data_reg[70] ;
 wire \mix1.data_reg[71] ;
 wire \mix1.data_reg[72] ;
 wire \mix1.data_reg[73] ;
 wire \mix1.data_reg[74] ;
 wire \mix1.data_reg[75] ;
 wire \mix1.data_reg[76] ;
 wire \mix1.data_reg[77] ;
 wire \mix1.data_reg[78] ;
 wire \mix1.data_reg[79] ;
 wire \mix1.data_reg[80] ;
 wire \mix1.data_reg[81] ;
 wire \mix1.data_reg[82] ;
 wire \mix1.data_reg[83] ;
 wire \mix1.data_reg[84] ;
 wire \mix1.data_reg[85] ;
 wire \mix1.data_reg[86] ;
 wire \mix1.data_reg[87] ;
 wire \mix1.data_reg[88] ;
 wire \mix1.data_reg[89] ;
 wire \mix1.data_reg[90] ;
 wire \mix1.data_reg[91] ;
 wire \mix1.data_reg[92] ;
 wire \mix1.data_reg[93] ;
 wire \mix1.data_reg[94] ;
 wire \mix1.data_reg[95] ;
 wire \mix1.data_reg[96] ;
 wire \mix1.data_reg[97] ;
 wire \mix1.data_reg[98] ;
 wire \mix1.data_reg[99] ;
 wire \mix1.next_ready_o ;
 wire \mix1.ready_o ;
 wire \mix1.state[0] ;
 wire \mix1.state[1] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire next_addroundkey_ready_o;
 wire next_addroundkey_start_i;
 wire next_first_round_reg;
 wire next_state;
 wire \round[0] ;
 wire \round[1] ;
 wire \round[2] ;
 wire \round[3] ;
 wire \sbox1.ah[0] ;
 wire \sbox1.ah[1] ;
 wire \sbox1.ah[2] ;
 wire \sbox1.ah[3] ;
 wire \sbox1.ah_reg[0] ;
 wire \sbox1.ah_reg[1] ;
 wire \sbox1.ah_reg[2] ;
 wire \sbox1.ah_reg[3] ;
 wire \sbox1.alph[0] ;
 wire \sbox1.alph[1] ;
 wire \sbox1.alph[2] ;
 wire \sbox1.alph[3] ;
 wire \sbox1.intermediate_to_invert_var[0] ;
 wire \sbox1.intermediate_to_invert_var[1] ;
 wire \sbox1.intermediate_to_invert_var[2] ;
 wire \sbox1.intermediate_to_invert_var[3] ;
 wire \sbox1.inversion_to_invert_var[0] ;
 wire \sbox1.inversion_to_invert_var[1] ;
 wire \sbox1.inversion_to_invert_var[2] ;
 wire \sbox1.inversion_to_invert_var[3] ;
 wire \sbox1.next_alph[0] ;
 wire \sbox1.next_alph[1] ;
 wire \sbox1.next_alph[2] ;
 wire \sbox1.next_alph[3] ;
 wire state;
 wire \sub1.data_o[0] ;
 wire \sub1.data_o[100] ;
 wire \sub1.data_o[101] ;
 wire \sub1.data_o[102] ;
 wire \sub1.data_o[103] ;
 wire \sub1.data_o[104] ;
 wire \sub1.data_o[105] ;
 wire \sub1.data_o[106] ;
 wire \sub1.data_o[107] ;
 wire \sub1.data_o[108] ;
 wire \sub1.data_o[109] ;
 wire \sub1.data_o[10] ;
 wire \sub1.data_o[110] ;
 wire \sub1.data_o[111] ;
 wire \sub1.data_o[112] ;
 wire \sub1.data_o[113] ;
 wire \sub1.data_o[114] ;
 wire \sub1.data_o[115] ;
 wire \sub1.data_o[116] ;
 wire \sub1.data_o[117] ;
 wire \sub1.data_o[118] ;
 wire \sub1.data_o[119] ;
 wire \sub1.data_o[11] ;
 wire \sub1.data_o[120] ;
 wire \sub1.data_o[121] ;
 wire \sub1.data_o[122] ;
 wire \sub1.data_o[123] ;
 wire \sub1.data_o[124] ;
 wire \sub1.data_o[125] ;
 wire \sub1.data_o[126] ;
 wire \sub1.data_o[127] ;
 wire \sub1.data_o[12] ;
 wire \sub1.data_o[13] ;
 wire \sub1.data_o[14] ;
 wire \sub1.data_o[15] ;
 wire \sub1.data_o[16] ;
 wire \sub1.data_o[17] ;
 wire \sub1.data_o[18] ;
 wire \sub1.data_o[19] ;
 wire \sub1.data_o[1] ;
 wire \sub1.data_o[20] ;
 wire \sub1.data_o[21] ;
 wire \sub1.data_o[22] ;
 wire \sub1.data_o[23] ;
 wire \sub1.data_o[24] ;
 wire \sub1.data_o[25] ;
 wire \sub1.data_o[26] ;
 wire \sub1.data_o[27] ;
 wire \sub1.data_o[28] ;
 wire \sub1.data_o[29] ;
 wire \sub1.data_o[2] ;
 wire \sub1.data_o[30] ;
 wire \sub1.data_o[31] ;
 wire \sub1.data_o[32] ;
 wire \sub1.data_o[33] ;
 wire \sub1.data_o[34] ;
 wire \sub1.data_o[35] ;
 wire \sub1.data_o[36] ;
 wire \sub1.data_o[37] ;
 wire \sub1.data_o[38] ;
 wire \sub1.data_o[39] ;
 wire \sub1.data_o[3] ;
 wire \sub1.data_o[40] ;
 wire \sub1.data_o[41] ;
 wire \sub1.data_o[42] ;
 wire \sub1.data_o[43] ;
 wire \sub1.data_o[44] ;
 wire \sub1.data_o[45] ;
 wire \sub1.data_o[46] ;
 wire \sub1.data_o[47] ;
 wire \sub1.data_o[48] ;
 wire \sub1.data_o[49] ;
 wire \sub1.data_o[4] ;
 wire \sub1.data_o[50] ;
 wire \sub1.data_o[51] ;
 wire \sub1.data_o[52] ;
 wire \sub1.data_o[53] ;
 wire \sub1.data_o[54] ;
 wire \sub1.data_o[55] ;
 wire \sub1.data_o[56] ;
 wire \sub1.data_o[57] ;
 wire \sub1.data_o[58] ;
 wire \sub1.data_o[59] ;
 wire \sub1.data_o[5] ;
 wire \sub1.data_o[60] ;
 wire \sub1.data_o[61] ;
 wire \sub1.data_o[62] ;
 wire \sub1.data_o[63] ;
 wire \sub1.data_o[64] ;
 wire \sub1.data_o[65] ;
 wire \sub1.data_o[66] ;
 wire \sub1.data_o[67] ;
 wire \sub1.data_o[68] ;
 wire \sub1.data_o[69] ;
 wire \sub1.data_o[6] ;
 wire \sub1.data_o[70] ;
 wire \sub1.data_o[71] ;
 wire \sub1.data_o[72] ;
 wire \sub1.data_o[73] ;
 wire \sub1.data_o[74] ;
 wire \sub1.data_o[75] ;
 wire \sub1.data_o[76] ;
 wire \sub1.data_o[77] ;
 wire \sub1.data_o[78] ;
 wire \sub1.data_o[79] ;
 wire \sub1.data_o[7] ;
 wire \sub1.data_o[80] ;
 wire \sub1.data_o[81] ;
 wire \sub1.data_o[82] ;
 wire \sub1.data_o[83] ;
 wire \sub1.data_o[84] ;
 wire \sub1.data_o[85] ;
 wire \sub1.data_o[86] ;
 wire \sub1.data_o[87] ;
 wire \sub1.data_o[88] ;
 wire \sub1.data_o[89] ;
 wire \sub1.data_o[8] ;
 wire \sub1.data_o[90] ;
 wire \sub1.data_o[91] ;
 wire \sub1.data_o[92] ;
 wire \sub1.data_o[93] ;
 wire \sub1.data_o[94] ;
 wire \sub1.data_o[95] ;
 wire \sub1.data_o[96] ;
 wire \sub1.data_o[97] ;
 wire \sub1.data_o[98] ;
 wire \sub1.data_o[99] ;
 wire \sub1.data_o[9] ;
 wire \sub1.next_ready_o ;
 wire \sub1.ready_o ;
 wire \sub1.state[0] ;
 wire \sub1.state[1] ;
 wire \sub1.state[2] ;
 wire \sub1.state[3] ;
 wire \sub1.state[4] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_03926_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(\fifo_bank_register.data_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(\fifo_bank_register.data_out[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(\fifo_bank_register.data_out[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(\fifo_bank_register.data_out[87] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_04391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(\fifo_bank_register.data_out[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(\fifo_bank_register.data_out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(\mix1.data_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(\mix1.data_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(\mix1.data_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(\mix1.data_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(\mix1.data_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(\mix1.data_o[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(\mix1.data_o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(\mix1.data_o[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_04435_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(\mix1.data_o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(\mix1.data_o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(\mix1.data_o[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(\mix1.data_o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(\mix1.data_o[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(\mix1.data_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(\mix1.data_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(\mix1.data_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(\mix1.data_o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(\mix1.data_o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_04470_));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(\mix1.data_o[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(\sub1.data_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(\sub1.data_o[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(\sub1.data_o[47] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_04487_));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_04492_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_04562_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_04573_));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_04577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_04577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(_04468_));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(_04490_));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(_04748_));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(_05757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_04577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(_05977_));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(\addroundkey_data_o[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(\addroundkey_data_o[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(\addroundkey_data_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(\addroundkey_data_o[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(\addroundkey_data_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(\addroundkey_data_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(\addroundkey_data_o[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(\addroundkey_data_o[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(\addroundkey_data_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_04591_));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(\fifo_bank_register.data_out[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(\fifo_bank_register.data_out[116] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(\fifo_bank_register.data_out[116] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(\mix1.data_o[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(\mix1.data_o[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(\mix1.data_o[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(\sub1.data_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(\sub1.data_o[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(\sub1.data_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(\sub1.data_o[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(\sub1.data_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(\sub1.data_o[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(\sub1.data_o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(\sub1.data_o[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(\sub1.data_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(\sub1.data_o[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_04606_));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(_04566_));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(_06485_));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(_06705_));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(\addroundkey_data_o[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_05245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_05547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_05553_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_05553_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_05553_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_05614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_05614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_05614_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_06368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\addroundkey_data_o[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\addroundkey_data_o[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\addroundkey_data_o[113] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\addroundkey_data_o[119] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\addroundkey_data_o[121] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\addroundkey_data_o[121] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\addroundkey_data_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\addroundkey_data_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\addroundkey_data_o[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_02208_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\addroundkey_data_o[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\addroundkey_data_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\addroundkey_data_o[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\addroundkey_data_o[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\addroundkey_data_o[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\addroundkey_data_o[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\addroundkey_data_o[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\addroundkey_data_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\addroundkey_data_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\addroundkey_data_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\addroundkey_data_o[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(\addroundkey_data_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(\addroundkey_data_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\addroundkey_data_o[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\addroundkey_data_o[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\addroundkey_data_o[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\addroundkey_data_o[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\addroundkey_data_o[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\addroundkey_data_o[64] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\addroundkey_data_o[67] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_03143_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(\addroundkey_data_o[69] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(\addroundkey_data_o[71] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(\addroundkey_data_o[71] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(\addroundkey_data_o[71] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(\addroundkey_data_o[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(\addroundkey_data_o[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(\addroundkey_data_o[79] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(\addroundkey_data_o[79] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(\fifo_bank_register.data_out[114] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(\fifo_bank_register.data_out[115] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_03926_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1060 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_157_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_158_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_159_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_159_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_160_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_161_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_162_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_162_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_163_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_1382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_164_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_164_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_164_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_165_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_166_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_166_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_167_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_167_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_168_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_168_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_168_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_170_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_170_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_170_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_171_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_171_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_172_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_1378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_174_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_174_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_174_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_175_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_176_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_176_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_176_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_177_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_178_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_178_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_178_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_179_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_179_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_179_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_180_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_180_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_180_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_181_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_182_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_182_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_182_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_183_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_183_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_183_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_184_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_184_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_184_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_185_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_185_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_186_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_186_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_187_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_187_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_188_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_188_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_188_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_189_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_189_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_189_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_190_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_190_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_191_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_191_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_192_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_192_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_192_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_193_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_195_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_195_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_196_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_196_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_196_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_198_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_198_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_198_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_199_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_199_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_199_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_200_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_200_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_200_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_201_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_202_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_203_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_205_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_205_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_206_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_206_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_206_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_207_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_207_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_210_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_212_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_215_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_217_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_218_1378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_218_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_220_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_225_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_1378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_226_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_226_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_1380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_227_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_227_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_227_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_228_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_228_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_228_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_229_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_229_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_229_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_898 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_4 _08202_ (.A(\sub1.state[1] ),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_4 _08203_ (.A(\sub1.state[0] ),
    .X(_04363_));
 sky130_fd_sc_hd__buf_2 _08204_ (.A(\sub1.state[3] ),
    .X(_04364_));
 sky130_fd_sc_hd__clkbuf_4 _08205_ (.A(\sub1.state[2] ),
    .X(_04365_));
 sky130_fd_sc_hd__nor4_1 _08206_ (.A(_04362_),
    .B(_04363_),
    .C(_04364_),
    .D(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2_2 _08207_ (.A(\sub1.state[4] ),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__inv_2 _08208_ (.A(_04367_),
    .Y(_04368_));
 sky130_fd_sc_hd__clkbuf_8 _08209_ (.A(_04368_),
    .X(_04369_));
 sky130_fd_sc_hd__clkbuf_4 _08210_ (.A(_04369_),
    .X(\sub1.next_ready_o ));
 sky130_fd_sc_hd__nor2_1 _08211_ (.A(\ks1.state[1] ),
    .B(\ks1.state[0] ),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2_4 _08212_ (.A(\ks1.state[2] ),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__inv_2 _08213_ (.A(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__buf_4 _08214_ (.A(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__buf_4 _08215_ (.A(_04373_),
    .X(\ks1.next_ready_o ));
 sky130_fd_sc_hd__and2_1 _08216_ (.A(\mix1.state[0] ),
    .B(\mix1.state[1] ),
    .X(_04374_));
 sky130_fd_sc_hd__clkbuf_4 _08217_ (.A(_04374_),
    .X(_04375_));
 sky130_fd_sc_hd__buf_4 _08218_ (.A(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__buf_4 _08219_ (.A(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__buf_4 _08220_ (.A(_04377_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_4 _08221_ (.A(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__buf_4 _08222_ (.A(_04379_),
    .X(\mix1.next_ready_o ));
 sky130_fd_sc_hd__or4_1 _08223_ (.A(net22),
    .B(net21),
    .C(net25),
    .D(net24),
    .X(_04380_));
 sky130_fd_sc_hd__or4_1 _08224_ (.A(net27),
    .B(net26),
    .C(net29),
    .D(net28),
    .X(_04381_));
 sky130_fd_sc_hd__or4b_1 _08225_ (.A(net31),
    .B(_04381_),
    .C(net30),
    .D_N(net594),
    .X(_04382_));
 sky130_fd_sc_hd__or4_1 _08226_ (.A(net9),
    .B(net8),
    .C(net11),
    .D(net10),
    .X(_04383_));
 sky130_fd_sc_hd__or4_1 _08227_ (.A(net5),
    .B(net4),
    .C(net7),
    .D(net6),
    .X(_04384_));
 sky130_fd_sc_hd__or4_1 _08228_ (.A(net14),
    .B(net13),
    .C(net16),
    .D(net15),
    .X(_04385_));
 sky130_fd_sc_hd__or4_1 _08229_ (.A(net18),
    .B(net17),
    .C(net20),
    .D(net19),
    .X(_04386_));
 sky130_fd_sc_hd__or4_1 _08230_ (.A(_04383_),
    .B(_04384_),
    .C(_04385_),
    .D(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__or4_1 _08231_ (.A(net119),
    .B(net118),
    .C(net121),
    .D(net120),
    .X(_04388_));
 sky130_fd_sc_hd__or4_1 _08232_ (.A(net114),
    .B(net113),
    .C(net116),
    .D(net115),
    .X(_04389_));
 sky130_fd_sc_hd__or4_1 _08233_ (.A(net123),
    .B(net122),
    .C(net125),
    .D(net124),
    .X(_04390_));
 sky130_fd_sc_hd__or4_2 _08234_ (.A(net127),
    .B(net126),
    .C(net3),
    .D(net2),
    .X(_04391_));
 sky130_fd_sc_hd__or4_1 _08235_ (.A(_04388_),
    .B(_04389_),
    .C(_04390_),
    .D(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__or4_4 _08236_ (.A(_04380_),
    .B(_04382_),
    .C(_04387_),
    .D(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__or4_4 _08237_ (.A(net66),
    .B(net65),
    .C(net68),
    .D(net67),
    .X(_04394_));
 sky130_fd_sc_hd__or4_1 _08238_ (.A(net61),
    .B(net60),
    .C(net64),
    .D(net63),
    .X(_04395_));
 sky130_fd_sc_hd__or4_1 _08239_ (.A(net70),
    .B(net69),
    .C(net72),
    .D(net71),
    .X(_04396_));
 sky130_fd_sc_hd__or4_1 _08240_ (.A(net75),
    .B(net74),
    .C(net77),
    .D(net76),
    .X(_04397_));
 sky130_fd_sc_hd__or4_1 _08241_ (.A(_04394_),
    .B(_04395_),
    .C(_04396_),
    .D(_04397_),
    .X(_04398_));
 sky130_fd_sc_hd__or4_1 _08242_ (.A(net48),
    .B(net47),
    .C(net50),
    .D(net49),
    .X(_04399_));
 sky130_fd_sc_hd__or4_1 _08243_ (.A(net44),
    .B(net43),
    .C(net46),
    .D(net45),
    .X(_04400_));
 sky130_fd_sc_hd__or4_1 _08244_ (.A(net53),
    .B(net52),
    .C(net55),
    .D(net54),
    .X(_04401_));
 sky130_fd_sc_hd__or4_1 _08245_ (.A(net57),
    .B(net56),
    .C(net59),
    .D(net58),
    .X(_04402_));
 sky130_fd_sc_hd__or4_1 _08246_ (.A(_04399_),
    .B(_04400_),
    .C(_04401_),
    .D(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__or4_1 _08247_ (.A(net83),
    .B(net82),
    .C(net86),
    .D(net85),
    .X(_04404_));
 sky130_fd_sc_hd__or4_1 _08248_ (.A(net79),
    .B(net78),
    .C(net81),
    .D(net80),
    .X(_04405_));
 sky130_fd_sc_hd__or4_1 _08249_ (.A(net88),
    .B(net87),
    .C(net90),
    .D(net89),
    .X(_04406_));
 sky130_fd_sc_hd__or4_1 _08250_ (.A(net92),
    .B(net91),
    .C(net94),
    .D(net93),
    .X(_04407_));
 sky130_fd_sc_hd__or4_1 _08251_ (.A(_04404_),
    .B(_04405_),
    .C(_04406_),
    .D(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__or4_1 _08252_ (.A(net101),
    .B(net100),
    .C(net103),
    .D(net102),
    .X(_04409_));
 sky130_fd_sc_hd__or4_2 _08253_ (.A(net97),
    .B(net96),
    .C(net99),
    .D(net98),
    .X(_04410_));
 sky130_fd_sc_hd__or4_1 _08254_ (.A(net105),
    .B(net104),
    .C(net108),
    .D(net107),
    .X(_04411_));
 sky130_fd_sc_hd__or4_1 _08255_ (.A(net110),
    .B(net109),
    .C(net112),
    .D(net111),
    .X(_04412_));
 sky130_fd_sc_hd__or4_2 _08256_ (.A(_04409_),
    .B(_04410_),
    .C(_04411_),
    .D(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__or4_1 _08257_ (.A(_04398_),
    .B(_04403_),
    .C(_04408_),
    .D(_04413_),
    .X(_04414_));
 sky130_fd_sc_hd__or4_1 _08258_ (.A(net23),
    .B(net12),
    .C(net33),
    .D(net32),
    .X(_04415_));
 sky130_fd_sc_hd__or4_1 _08259_ (.A(net106),
    .B(net95),
    .C(net128),
    .D(net117),
    .X(_04416_));
 sky130_fd_sc_hd__or4_1 _08260_ (.A(net35),
    .B(net34),
    .C(net37),
    .D(net36),
    .X(_04417_));
 sky130_fd_sc_hd__or4_1 _08261_ (.A(net39),
    .B(net38),
    .C(net42),
    .D(net41),
    .X(_04418_));
 sky130_fd_sc_hd__or4_1 _08262_ (.A(_04415_),
    .B(_04416_),
    .C(_04417_),
    .D(_04418_),
    .X(_04419_));
 sky130_fd_sc_hd__or4bb_4 _08263_ (.A(net156),
    .B(net158),
    .C_N(net157),
    .D_N(net155),
    .X(_04420_));
 sky130_fd_sc_hd__or4b_1 _08264_ (.A(net151),
    .B(net154),
    .C(net153),
    .D_N(net150),
    .X(_04421_));
 sky130_fd_sc_hd__or4b_1 _08265_ (.A(net160),
    .B(net40),
    .C(net1),
    .D_N(net159),
    .X(_04422_));
 sky130_fd_sc_hd__or4_1 _08266_ (.A(net62),
    .B(net51),
    .C(net84),
    .D(net73),
    .X(_04423_));
 sky130_fd_sc_hd__or4_1 _08267_ (.A(_04420_),
    .B(_04421_),
    .C(_04422_),
    .D(_04423_),
    .X(_04424_));
 sky130_fd_sc_hd__and4b_1 _08268_ (.A_N(net139),
    .B(net140),
    .C(net138),
    .D(net137),
    .X(_04425_));
 sky130_fd_sc_hd__and4b_1 _08269_ (.A_N(net134),
    .B(net133),
    .C(net136),
    .D(net135),
    .X(_04426_));
 sky130_fd_sc_hd__nand2_1 _08270_ (.A(_04425_),
    .B(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__or4bb_1 _08271_ (.A(net143),
    .B(net144),
    .C_N(net145),
    .D_N(net142),
    .X(_04428_));
 sky130_fd_sc_hd__or4bb_1 _08272_ (.A(net147),
    .B(net146),
    .C_N(net149),
    .D_N(net148),
    .X(_04429_));
 sky130_fd_sc_hd__or4b_1 _08273_ (.A(net248),
    .B(net247),
    .C(net249),
    .D_N(net250),
    .X(_04430_));
 sky130_fd_sc_hd__or4bb_1 _08274_ (.A(net243),
    .B(net245),
    .C_N(net244),
    .D_N(net242),
    .X(_04431_));
 sky130_fd_sc_hd__or4bb_1 _08275_ (.A(net252),
    .B(net253),
    .C_N(net254),
    .D_N(net251),
    .X(_04432_));
 sky130_fd_sc_hd__or4bb_1 _08276_ (.A(net255),
    .B(net131),
    .C_N(net132),
    .D_N(net256),
    .X(_04433_));
 sky130_fd_sc_hd__or4_1 _08277_ (.A(_04430_),
    .B(_04431_),
    .C(_04432_),
    .D(_04433_),
    .X(_04434_));
 sky130_fd_sc_hd__or4_4 _08278_ (.A(_04427_),
    .B(_04428_),
    .C(_04429_),
    .D(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__or4_4 _08279_ (.A(_04414_),
    .B(_04419_),
    .C(_04424_),
    .D(_04435_),
    .X(_04436_));
 sky130_fd_sc_hd__and4b_1 _08280_ (.A_N(net202),
    .B(net213),
    .C(net191),
    .D(net180),
    .X(_04437_));
 sky130_fd_sc_hd__nand3b_1 _08281_ (.A_N(net130),
    .B(net169),
    .C(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__and4b_1 _08282_ (.A_N(net161),
    .B(net162),
    .C(net152),
    .D(net141),
    .X(_04439_));
 sky130_fd_sc_hd__and4b_1 _08283_ (.A_N(net235),
    .B(net224),
    .C(net257),
    .D(net246),
    .X(_04440_));
 sky130_fd_sc_hd__nand2_1 _08284_ (.A(_04439_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__or4bb_1 _08285_ (.A(net164),
    .B(net166),
    .C_N(net165),
    .D_N(net163),
    .X(_04442_));
 sky130_fd_sc_hd__or4bb_1 _08286_ (.A(net167),
    .B(net170),
    .C_N(net171),
    .D_N(net168),
    .X(_04443_));
 sky130_fd_sc_hd__or4_2 _08287_ (.A(_04438_),
    .B(_04441_),
    .C(_04442_),
    .D(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__nand4b_1 _08288_ (.A_N(net212),
    .B(net211),
    .C(net215),
    .D(net214),
    .Y(_04445_));
 sky130_fd_sc_hd__or4b_1 _08289_ (.A(net208),
    .B(net210),
    .C(net209),
    .D_N(net207),
    .X(_04446_));
 sky130_fd_sc_hd__nand4b_1 _08290_ (.A_N(net217),
    .B(net216),
    .C(net219),
    .D(net218),
    .Y(_04447_));
 sky130_fd_sc_hd__or4b_1 _08291_ (.A(net221),
    .B(net220),
    .C(net222),
    .D_N(net223),
    .X(_04448_));
 sky130_fd_sc_hd__or4_1 _08292_ (.A(_04445_),
    .B(_04446_),
    .C(_04447_),
    .D(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__or4_1 _08293_ (.A(net230),
    .B(net229),
    .C(net232),
    .D(net231),
    .X(_04450_));
 sky130_fd_sc_hd__or4bb_1 _08294_ (.A(net226),
    .B(net228),
    .C_N(net227),
    .D_N(net225),
    .X(_04451_));
 sky130_fd_sc_hd__or4bb_1 _08295_ (.A(net234),
    .B(net236),
    .C_N(net237),
    .D_N(net233),
    .X(_04452_));
 sky130_fd_sc_hd__and4b_1 _08296_ (.A_N(net240),
    .B(net241),
    .C(net239),
    .D(net238),
    .X(_04453_));
 sky130_fd_sc_hd__or4b_1 _08297_ (.A(_04450_),
    .B(_04451_),
    .C(_04452_),
    .D_N(_04453_),
    .X(_04454_));
 sky130_fd_sc_hd__nand4b_1 _08298_ (.A_N(net195),
    .B(net194),
    .C(net197),
    .D(net196),
    .Y(_04455_));
 sky130_fd_sc_hd__or4bb_1 _08299_ (.A(net190),
    .B(net192),
    .C_N(net193),
    .D_N(net189),
    .X(_04456_));
 sky130_fd_sc_hd__or4bb_1 _08300_ (.A(net199),
    .B(net201),
    .C_N(net200),
    .D_N(net198),
    .X(_04457_));
 sky130_fd_sc_hd__or4bb_1 _08301_ (.A(net203),
    .B(net205),
    .C_N(net206),
    .D_N(net204),
    .X(_04458_));
 sky130_fd_sc_hd__or4_1 _08302_ (.A(_04455_),
    .B(_04456_),
    .C(_04457_),
    .D(_04458_),
    .X(_04459_));
 sky130_fd_sc_hd__nand4b_1 _08303_ (.A_N(net177),
    .B(net176),
    .C(net179),
    .D(net178),
    .Y(_04460_));
 sky130_fd_sc_hd__or4b_1 _08304_ (.A(net173),
    .B(net175),
    .C(net174),
    .D_N(net172),
    .X(_04461_));
 sky130_fd_sc_hd__or4bb_1 _08305_ (.A(net182),
    .B(net184),
    .C_N(net183),
    .D_N(net181),
    .X(_04462_));
 sky130_fd_sc_hd__or4b_1 _08306_ (.A(net186),
    .B(net185),
    .C(net187),
    .D_N(net188),
    .X(_04463_));
 sky130_fd_sc_hd__or4_1 _08307_ (.A(_04460_),
    .B(_04461_),
    .C(_04462_),
    .D(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__or4_2 _08308_ (.A(_04449_),
    .B(_04454_),
    .C(_04459_),
    .D(_04464_),
    .X(_04465_));
 sky130_fd_sc_hd__nor4_4 _08309_ (.A(_04393_),
    .B(_04436_),
    .C(_04444_),
    .D(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__buf_8 _08310_ (.A(_04466_),
    .X(_04467_));
 sky130_fd_sc_hd__buf_12 _08311_ (.A(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__mux2_1 _08312_ (.A0(\addroundkey_data_o[0] ),
    .A1(\fifo_bank_register.data_out[0] ),
    .S(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__buf_1 _08313_ (.A(_04469_),
    .X(net260));
 sky130_fd_sc_hd__mux2_2 _08314_ (.A0(\addroundkey_data_o[1] ),
    .A1(\fifo_bank_register.data_out[1] ),
    .S(_04468_),
    .X(_04470_));
 sky130_fd_sc_hd__clkbuf_1 _08315_ (.A(_04470_),
    .X(net299));
 sky130_fd_sc_hd__mux2_2 _08316_ (.A0(\addroundkey_data_o[2] ),
    .A1(\fifo_bank_register.data_out[2] ),
    .S(_04468_),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_1 _08317_ (.A(_04471_),
    .X(net310));
 sky130_fd_sc_hd__mux2_1 _08318_ (.A0(\addroundkey_data_o[3] ),
    .A1(\fifo_bank_register.data_out[3] ),
    .S(_04468_),
    .X(_04472_));
 sky130_fd_sc_hd__clkbuf_2 _08319_ (.A(_04472_),
    .X(net321));
 sky130_fd_sc_hd__mux2_1 _08320_ (.A0(\addroundkey_data_o[4] ),
    .A1(\fifo_bank_register.data_out[4] ),
    .S(_04468_),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_1 _08321_ (.A(_04473_),
    .X(net332));
 sky130_fd_sc_hd__mux2_2 _08322_ (.A0(\addroundkey_data_o[5] ),
    .A1(\fifo_bank_register.data_out[5] ),
    .S(_04468_),
    .X(_04474_));
 sky130_fd_sc_hd__clkbuf_1 _08323_ (.A(_04474_),
    .X(net343));
 sky130_fd_sc_hd__mux2_1 _08324_ (.A0(\addroundkey_data_o[6] ),
    .A1(\fifo_bank_register.data_out[6] ),
    .S(_04468_),
    .X(_04475_));
 sky130_fd_sc_hd__buf_2 _08325_ (.A(_04475_),
    .X(net354));
 sky130_fd_sc_hd__mux2_1 _08326_ (.A0(\addroundkey_data_o[7] ),
    .A1(\fifo_bank_register.data_out[7] ),
    .S(_04468_),
    .X(_04476_));
 sky130_fd_sc_hd__buf_2 _08327_ (.A(_04476_),
    .X(net365));
 sky130_fd_sc_hd__mux2_1 _08328_ (.A0(\addroundkey_data_o[8] ),
    .A1(\fifo_bank_register.data_out[8] ),
    .S(_04468_),
    .X(_04477_));
 sky130_fd_sc_hd__buf_2 _08329_ (.A(_04477_),
    .X(net376));
 sky130_fd_sc_hd__buf_6 _08330_ (.A(_04466_),
    .X(_04478_));
 sky130_fd_sc_hd__clkbuf_16 _08331_ (.A(_04478_),
    .X(_04479_));
 sky130_fd_sc_hd__mux2_1 _08332_ (.A0(\addroundkey_data_o[9] ),
    .A1(\fifo_bank_register.data_out[9] ),
    .S(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__buf_1 _08333_ (.A(_04480_),
    .X(net387));
 sky130_fd_sc_hd__mux2_2 _08334_ (.A0(\addroundkey_data_o[10] ),
    .A1(\fifo_bank_register.data_out[10] ),
    .S(_04479_),
    .X(_04481_));
 sky130_fd_sc_hd__clkbuf_1 _08335_ (.A(_04481_),
    .X(net271));
 sky130_fd_sc_hd__mux2_2 _08336_ (.A0(\addroundkey_data_o[11] ),
    .A1(\fifo_bank_register.data_out[11] ),
    .S(_04479_),
    .X(_04482_));
 sky130_fd_sc_hd__clkbuf_1 _08337_ (.A(_04482_),
    .X(net282));
 sky130_fd_sc_hd__mux2_4 _08338_ (.A0(\addroundkey_data_o[12] ),
    .A1(\fifo_bank_register.data_out[12] ),
    .S(_04479_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_1 _08339_ (.A(_04483_),
    .X(net291));
 sky130_fd_sc_hd__mux2_1 _08340_ (.A0(\addroundkey_data_o[13] ),
    .A1(\fifo_bank_register.data_out[13] ),
    .S(_04479_),
    .X(_04484_));
 sky130_fd_sc_hd__clkbuf_2 _08341_ (.A(_04484_),
    .X(net292));
 sky130_fd_sc_hd__mux2_2 _08342_ (.A0(\addroundkey_data_o[14] ),
    .A1(\fifo_bank_register.data_out[14] ),
    .S(_04479_),
    .X(_04485_));
 sky130_fd_sc_hd__clkbuf_1 _08343_ (.A(_04485_),
    .X(net293));
 sky130_fd_sc_hd__mux2_2 _08344_ (.A0(\addroundkey_data_o[15] ),
    .A1(\fifo_bank_register.data_out[15] ),
    .S(_04479_),
    .X(_04486_));
 sky130_fd_sc_hd__clkbuf_2 _08345_ (.A(_04486_),
    .X(net294));
 sky130_fd_sc_hd__mux2_4 _08346_ (.A0(\addroundkey_data_o[16] ),
    .A1(\fifo_bank_register.data_out[16] ),
    .S(_04479_),
    .X(_04487_));
 sky130_fd_sc_hd__clkbuf_1 _08347_ (.A(_04487_),
    .X(net295));
 sky130_fd_sc_hd__mux2_2 _08348_ (.A0(\addroundkey_data_o[17] ),
    .A1(\fifo_bank_register.data_out[17] ),
    .S(_04479_),
    .X(_04488_));
 sky130_fd_sc_hd__clkbuf_1 _08349_ (.A(_04488_),
    .X(net296));
 sky130_fd_sc_hd__mux2_1 _08350_ (.A0(\addroundkey_data_o[18] ),
    .A1(\fifo_bank_register.data_out[18] ),
    .S(_04479_),
    .X(_04489_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08351_ (.A(_04489_),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_16 _08352_ (.A(_04478_),
    .X(_04490_));
 sky130_fd_sc_hd__mux2_2 _08353_ (.A0(\addroundkey_data_o[19] ),
    .A1(\fifo_bank_register.data_out[19] ),
    .S(_04490_),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _08354_ (.A(_04491_),
    .X(net298));
 sky130_fd_sc_hd__mux2_4 _08355_ (.A0(\addroundkey_data_o[20] ),
    .A1(\fifo_bank_register.data_out[20] ),
    .S(_04490_),
    .X(_04492_));
 sky130_fd_sc_hd__clkbuf_1 _08356_ (.A(_04492_),
    .X(net300));
 sky130_fd_sc_hd__mux2_1 _08357_ (.A0(\addroundkey_data_o[21] ),
    .A1(\fifo_bank_register.data_out[21] ),
    .S(_04490_),
    .X(_04493_));
 sky130_fd_sc_hd__clkbuf_2 _08358_ (.A(_04493_),
    .X(net301));
 sky130_fd_sc_hd__mux2_1 _08359_ (.A0(\addroundkey_data_o[22] ),
    .A1(\fifo_bank_register.data_out[22] ),
    .S(_04490_),
    .X(_04494_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08360_ (.A(_04494_),
    .X(net302));
 sky130_fd_sc_hd__mux2_1 _08361_ (.A0(\addroundkey_data_o[23] ),
    .A1(\fifo_bank_register.data_out[23] ),
    .S(_04490_),
    .X(_04495_));
 sky130_fd_sc_hd__clkbuf_1 _08362_ (.A(_04495_),
    .X(net303));
 sky130_fd_sc_hd__mux2_1 _08363_ (.A0(\addroundkey_data_o[24] ),
    .A1(\fifo_bank_register.data_out[24] ),
    .S(_04490_),
    .X(_04496_));
 sky130_fd_sc_hd__clkbuf_1 _08364_ (.A(_04496_),
    .X(net304));
 sky130_fd_sc_hd__mux2_1 _08365_ (.A0(\addroundkey_data_o[25] ),
    .A1(\fifo_bank_register.data_out[25] ),
    .S(_04490_),
    .X(_04497_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08366_ (.A(_04497_),
    .X(net305));
 sky130_fd_sc_hd__mux2_2 _08367_ (.A0(\addroundkey_data_o[26] ),
    .A1(\fifo_bank_register.data_out[26] ),
    .S(_04490_),
    .X(_04498_));
 sky130_fd_sc_hd__clkbuf_1 _08368_ (.A(_04498_),
    .X(net306));
 sky130_fd_sc_hd__mux2_4 _08369_ (.A0(\addroundkey_data_o[27] ),
    .A1(\fifo_bank_register.data_out[27] ),
    .S(_04490_),
    .X(_04499_));
 sky130_fd_sc_hd__clkbuf_1 _08370_ (.A(_04499_),
    .X(net307));
 sky130_fd_sc_hd__mux2_1 _08371_ (.A0(\addroundkey_data_o[28] ),
    .A1(\fifo_bank_register.data_out[28] ),
    .S(_04490_),
    .X(_04500_));
 sky130_fd_sc_hd__clkbuf_2 _08372_ (.A(_04500_),
    .X(net308));
 sky130_fd_sc_hd__buf_8 _08373_ (.A(_04478_),
    .X(_04501_));
 sky130_fd_sc_hd__mux2_1 _08374_ (.A0(\addroundkey_data_o[29] ),
    .A1(\fifo_bank_register.data_out[29] ),
    .S(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__clkbuf_1 _08375_ (.A(_04502_),
    .X(net309));
 sky130_fd_sc_hd__mux2_2 _08376_ (.A0(\addroundkey_data_o[30] ),
    .A1(\fifo_bank_register.data_out[30] ),
    .S(_04501_),
    .X(_04503_));
 sky130_fd_sc_hd__clkbuf_1 _08377_ (.A(_04503_),
    .X(net311));
 sky130_fd_sc_hd__mux2_2 _08378_ (.A0(\addroundkey_data_o[31] ),
    .A1(\fifo_bank_register.data_out[31] ),
    .S(_04501_),
    .X(_04504_));
 sky130_fd_sc_hd__clkbuf_1 _08379_ (.A(_04504_),
    .X(net312));
 sky130_fd_sc_hd__mux2_1 _08380_ (.A0(\addroundkey_data_o[32] ),
    .A1(\fifo_bank_register.data_out[32] ),
    .S(_04501_),
    .X(_04505_));
 sky130_fd_sc_hd__clkbuf_2 _08381_ (.A(_04505_),
    .X(net313));
 sky130_fd_sc_hd__mux2_4 _08382_ (.A0(\addroundkey_data_o[33] ),
    .A1(\fifo_bank_register.data_out[33] ),
    .S(_04501_),
    .X(_04506_));
 sky130_fd_sc_hd__clkbuf_1 _08383_ (.A(_04506_),
    .X(net314));
 sky130_fd_sc_hd__mux2_1 _08384_ (.A0(\addroundkey_data_o[34] ),
    .A1(\fifo_bank_register.data_out[34] ),
    .S(_04501_),
    .X(_04507_));
 sky130_fd_sc_hd__clkbuf_2 _08385_ (.A(_04507_),
    .X(net315));
 sky130_fd_sc_hd__mux2_2 _08386_ (.A0(\addroundkey_data_o[35] ),
    .A1(\fifo_bank_register.data_out[35] ),
    .S(_04501_),
    .X(_04508_));
 sky130_fd_sc_hd__clkbuf_1 _08387_ (.A(_04508_),
    .X(net316));
 sky130_fd_sc_hd__mux2_2 _08388_ (.A0(\addroundkey_data_o[36] ),
    .A1(\fifo_bank_register.data_out[36] ),
    .S(_04501_),
    .X(_04509_));
 sky130_fd_sc_hd__clkbuf_1 _08389_ (.A(_04509_),
    .X(net317));
 sky130_fd_sc_hd__mux2_2 _08390_ (.A0(\addroundkey_data_o[37] ),
    .A1(\fifo_bank_register.data_out[37] ),
    .S(_04501_),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_2 _08391_ (.A(_04510_),
    .X(net318));
 sky130_fd_sc_hd__mux2_2 _08392_ (.A0(\addroundkey_data_o[38] ),
    .A1(\fifo_bank_register.data_out[38] ),
    .S(_04501_),
    .X(_04511_));
 sky130_fd_sc_hd__clkbuf_1 _08393_ (.A(_04511_),
    .X(net319));
 sky130_fd_sc_hd__buf_8 _08394_ (.A(_04478_),
    .X(_04512_));
 sky130_fd_sc_hd__mux2_1 _08395_ (.A0(\addroundkey_data_o[39] ),
    .A1(\fifo_bank_register.data_out[39] ),
    .S(_04512_),
    .X(_04513_));
 sky130_fd_sc_hd__clkbuf_1 _08396_ (.A(_04513_),
    .X(net320));
 sky130_fd_sc_hd__mux2_1 _08397_ (.A0(\addroundkey_data_o[40] ),
    .A1(\fifo_bank_register.data_out[40] ),
    .S(_04512_),
    .X(_04514_));
 sky130_fd_sc_hd__clkbuf_2 _08398_ (.A(_04514_),
    .X(net322));
 sky130_fd_sc_hd__mux2_2 _08399_ (.A0(\addroundkey_data_o[41] ),
    .A1(\fifo_bank_register.data_out[41] ),
    .S(_04512_),
    .X(_04515_));
 sky130_fd_sc_hd__clkbuf_1 _08400_ (.A(_04515_),
    .X(net323));
 sky130_fd_sc_hd__mux2_2 _08401_ (.A0(\addroundkey_data_o[42] ),
    .A1(\fifo_bank_register.data_out[42] ),
    .S(_04512_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_1 _08402_ (.A(_04516_),
    .X(net324));
 sky130_fd_sc_hd__mux2_4 _08403_ (.A0(\addroundkey_data_o[43] ),
    .A1(\fifo_bank_register.data_out[43] ),
    .S(_04512_),
    .X(_04517_));
 sky130_fd_sc_hd__clkbuf_1 _08404_ (.A(_04517_),
    .X(net325));
 sky130_fd_sc_hd__mux2_2 _08405_ (.A0(\addroundkey_data_o[44] ),
    .A1(\fifo_bank_register.data_out[44] ),
    .S(_04512_),
    .X(_04518_));
 sky130_fd_sc_hd__clkbuf_1 _08406_ (.A(_04518_),
    .X(net326));
 sky130_fd_sc_hd__mux2_2 _08407_ (.A0(\addroundkey_data_o[45] ),
    .A1(\fifo_bank_register.data_out[45] ),
    .S(_04512_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _08408_ (.A(_04519_),
    .X(net327));
 sky130_fd_sc_hd__mux2_2 _08409_ (.A0(\addroundkey_data_o[46] ),
    .A1(\fifo_bank_register.data_out[46] ),
    .S(_04512_),
    .X(_04520_));
 sky130_fd_sc_hd__clkbuf_1 _08410_ (.A(_04520_),
    .X(net328));
 sky130_fd_sc_hd__mux2_4 _08411_ (.A0(\addroundkey_data_o[47] ),
    .A1(\fifo_bank_register.data_out[47] ),
    .S(_04512_),
    .X(_04521_));
 sky130_fd_sc_hd__clkbuf_1 _08412_ (.A(_04521_),
    .X(net329));
 sky130_fd_sc_hd__mux2_1 _08413_ (.A0(\addroundkey_data_o[48] ),
    .A1(\fifo_bank_register.data_out[48] ),
    .S(_04512_),
    .X(_04522_));
 sky130_fd_sc_hd__clkbuf_1 _08414_ (.A(_04522_),
    .X(net330));
 sky130_fd_sc_hd__buf_12 _08415_ (.A(_04478_),
    .X(_04523_));
 sky130_fd_sc_hd__mux2_1 _08416_ (.A0(\addroundkey_data_o[49] ),
    .A1(\fifo_bank_register.data_out[49] ),
    .S(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__buf_1 _08417_ (.A(_04524_),
    .X(net331));
 sky130_fd_sc_hd__mux2_1 _08418_ (.A0(\addroundkey_data_o[50] ),
    .A1(\fifo_bank_register.data_out[50] ),
    .S(_04523_),
    .X(_04525_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08419_ (.A(_04525_),
    .X(net333));
 sky130_fd_sc_hd__mux2_1 _08420_ (.A0(\addroundkey_data_o[51] ),
    .A1(\fifo_bank_register.data_out[51] ),
    .S(_04523_),
    .X(_04526_));
 sky130_fd_sc_hd__buf_1 _08421_ (.A(_04526_),
    .X(net334));
 sky130_fd_sc_hd__mux2_2 _08422_ (.A0(\addroundkey_data_o[52] ),
    .A1(\fifo_bank_register.data_out[52] ),
    .S(_04523_),
    .X(_04527_));
 sky130_fd_sc_hd__clkbuf_1 _08423_ (.A(_04527_),
    .X(net335));
 sky130_fd_sc_hd__mux2_1 _08424_ (.A0(\addroundkey_data_o[53] ),
    .A1(\fifo_bank_register.data_out[53] ),
    .S(_04523_),
    .X(_04528_));
 sky130_fd_sc_hd__buf_1 _08425_ (.A(_04528_),
    .X(net336));
 sky130_fd_sc_hd__mux2_4 _08426_ (.A0(\addroundkey_data_o[54] ),
    .A1(\fifo_bank_register.data_out[54] ),
    .S(_04523_),
    .X(_04529_));
 sky130_fd_sc_hd__clkbuf_1 _08427_ (.A(_04529_),
    .X(net337));
 sky130_fd_sc_hd__mux2_1 _08428_ (.A0(\addroundkey_data_o[55] ),
    .A1(\fifo_bank_register.data_out[55] ),
    .S(_04523_),
    .X(_04530_));
 sky130_fd_sc_hd__buf_1 _08429_ (.A(_04530_),
    .X(net338));
 sky130_fd_sc_hd__mux2_1 _08430_ (.A0(\addroundkey_data_o[56] ),
    .A1(\fifo_bank_register.data_out[56] ),
    .S(_04523_),
    .X(_04531_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08431_ (.A(_04531_),
    .X(net339));
 sky130_fd_sc_hd__mux2_2 _08432_ (.A0(\addroundkey_data_o[57] ),
    .A1(\fifo_bank_register.data_out[57] ),
    .S(_04523_),
    .X(_04532_));
 sky130_fd_sc_hd__clkbuf_1 _08433_ (.A(_04532_),
    .X(net340));
 sky130_fd_sc_hd__mux2_2 _08434_ (.A0(\addroundkey_data_o[58] ),
    .A1(\fifo_bank_register.data_out[58] ),
    .S(_04523_),
    .X(_04533_));
 sky130_fd_sc_hd__buf_1 _08435_ (.A(_04533_),
    .X(net341));
 sky130_fd_sc_hd__buf_8 _08436_ (.A(_04478_),
    .X(_04534_));
 sky130_fd_sc_hd__mux2_2 _08437_ (.A0(\addroundkey_data_o[59] ),
    .A1(\fifo_bank_register.data_out[59] ),
    .S(_04534_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_2 _08438_ (.A(_04535_),
    .X(net342));
 sky130_fd_sc_hd__mux2_1 _08439_ (.A0(\addroundkey_data_o[60] ),
    .A1(\fifo_bank_register.data_out[60] ),
    .S(_04534_),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_1 _08440_ (.A(_04536_),
    .X(net344));
 sky130_fd_sc_hd__mux2_1 _08441_ (.A0(\addroundkey_data_o[61] ),
    .A1(\fifo_bank_register.data_out[61] ),
    .S(_04534_),
    .X(_04537_));
 sky130_fd_sc_hd__clkbuf_1 _08442_ (.A(_04537_),
    .X(net345));
 sky130_fd_sc_hd__mux2_1 _08443_ (.A0(\addroundkey_data_o[62] ),
    .A1(\fifo_bank_register.data_out[62] ),
    .S(_04534_),
    .X(_04538_));
 sky130_fd_sc_hd__clkbuf_1 _08444_ (.A(_04538_),
    .X(net346));
 sky130_fd_sc_hd__mux2_1 _08445_ (.A0(\addroundkey_data_o[63] ),
    .A1(\fifo_bank_register.data_out[63] ),
    .S(_04534_),
    .X(_04539_));
 sky130_fd_sc_hd__clkbuf_1 _08446_ (.A(_04539_),
    .X(net347));
 sky130_fd_sc_hd__mux2_2 _08447_ (.A0(\addroundkey_data_o[64] ),
    .A1(\fifo_bank_register.data_out[64] ),
    .S(_04534_),
    .X(_04540_));
 sky130_fd_sc_hd__buf_1 _08448_ (.A(_04540_),
    .X(net348));
 sky130_fd_sc_hd__mux2_4 _08449_ (.A0(\addroundkey_data_o[65] ),
    .A1(\fifo_bank_register.data_out[65] ),
    .S(_04534_),
    .X(_04541_));
 sky130_fd_sc_hd__clkbuf_2 _08450_ (.A(_04541_),
    .X(net349));
 sky130_fd_sc_hd__mux2_1 _08451_ (.A0(\addroundkey_data_o[66] ),
    .A1(\fifo_bank_register.data_out[66] ),
    .S(_04534_),
    .X(_04542_));
 sky130_fd_sc_hd__clkbuf_1 _08452_ (.A(_04542_),
    .X(net350));
 sky130_fd_sc_hd__mux2_1 _08453_ (.A0(\addroundkey_data_o[67] ),
    .A1(\fifo_bank_register.data_out[67] ),
    .S(_04534_),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_1 _08454_ (.A(_04543_),
    .X(net351));
 sky130_fd_sc_hd__mux2_1 _08455_ (.A0(\addroundkey_data_o[68] ),
    .A1(\fifo_bank_register.data_out[68] ),
    .S(_04534_),
    .X(_04544_));
 sky130_fd_sc_hd__clkbuf_1 _08456_ (.A(_04544_),
    .X(net352));
 sky130_fd_sc_hd__buf_8 _08457_ (.A(_04478_),
    .X(_04545_));
 sky130_fd_sc_hd__mux2_1 _08458_ (.A0(\addroundkey_data_o[69] ),
    .A1(\fifo_bank_register.data_out[69] ),
    .S(_04545_),
    .X(_04546_));
 sky130_fd_sc_hd__buf_2 _08459_ (.A(_04546_),
    .X(net353));
 sky130_fd_sc_hd__mux2_1 _08460_ (.A0(\addroundkey_data_o[70] ),
    .A1(\fifo_bank_register.data_out[70] ),
    .S(_04545_),
    .X(_04547_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08461_ (.A(_04547_),
    .X(net355));
 sky130_fd_sc_hd__mux2_1 _08462_ (.A0(\addroundkey_data_o[71] ),
    .A1(\fifo_bank_register.data_out[71] ),
    .S(_04545_),
    .X(_04548_));
 sky130_fd_sc_hd__clkbuf_2 _08463_ (.A(_04548_),
    .X(net356));
 sky130_fd_sc_hd__mux2_1 _08464_ (.A0(\addroundkey_data_o[72] ),
    .A1(\fifo_bank_register.data_out[72] ),
    .S(_04545_),
    .X(_04549_));
 sky130_fd_sc_hd__buf_1 _08465_ (.A(_04549_),
    .X(net357));
 sky130_fd_sc_hd__mux2_2 _08466_ (.A0(\addroundkey_data_o[73] ),
    .A1(\fifo_bank_register.data_out[73] ),
    .S(_04545_),
    .X(_04550_));
 sky130_fd_sc_hd__buf_1 _08467_ (.A(_04550_),
    .X(net358));
 sky130_fd_sc_hd__mux2_2 _08468_ (.A0(\addroundkey_data_o[74] ),
    .A1(\fifo_bank_register.data_out[74] ),
    .S(_04545_),
    .X(_04551_));
 sky130_fd_sc_hd__clkbuf_1 _08469_ (.A(_04551_),
    .X(net359));
 sky130_fd_sc_hd__mux2_2 _08470_ (.A0(\addroundkey_data_o[75] ),
    .A1(\fifo_bank_register.data_out[75] ),
    .S(_04545_),
    .X(_04552_));
 sky130_fd_sc_hd__clkbuf_1 _08471_ (.A(_04552_),
    .X(net360));
 sky130_fd_sc_hd__mux2_1 _08472_ (.A0(\addroundkey_data_o[76] ),
    .A1(\fifo_bank_register.data_out[76] ),
    .S(_04545_),
    .X(_04553_));
 sky130_fd_sc_hd__clkbuf_2 _08473_ (.A(_04553_),
    .X(net361));
 sky130_fd_sc_hd__mux2_1 _08474_ (.A0(\addroundkey_data_o[77] ),
    .A1(\fifo_bank_register.data_out[77] ),
    .S(_04545_),
    .X(_04554_));
 sky130_fd_sc_hd__buf_1 _08475_ (.A(_04554_),
    .X(net362));
 sky130_fd_sc_hd__mux2_1 _08476_ (.A0(\addroundkey_data_o[78] ),
    .A1(\fifo_bank_register.data_out[78] ),
    .S(_04545_),
    .X(_04555_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08477_ (.A(_04555_),
    .X(net363));
 sky130_fd_sc_hd__buf_8 _08478_ (.A(_04478_),
    .X(_04556_));
 sky130_fd_sc_hd__mux2_1 _08479_ (.A0(\addroundkey_data_o[79] ),
    .A1(\fifo_bank_register.data_out[79] ),
    .S(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__clkbuf_2 _08480_ (.A(_04557_),
    .X(net364));
 sky130_fd_sc_hd__mux2_2 _08481_ (.A0(\addroundkey_data_o[80] ),
    .A1(\fifo_bank_register.data_out[80] ),
    .S(_04556_),
    .X(_04558_));
 sky130_fd_sc_hd__clkbuf_1 _08482_ (.A(_04558_),
    .X(net366));
 sky130_fd_sc_hd__mux2_2 _08483_ (.A0(\addroundkey_data_o[81] ),
    .A1(\fifo_bank_register.data_out[81] ),
    .S(_04556_),
    .X(_04559_));
 sky130_fd_sc_hd__clkbuf_1 _08484_ (.A(_04559_),
    .X(net367));
 sky130_fd_sc_hd__mux2_1 _08485_ (.A0(\addroundkey_data_o[82] ),
    .A1(\fifo_bank_register.data_out[82] ),
    .S(_04556_),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_1 _08486_ (.A(_04560_),
    .X(net368));
 sky130_fd_sc_hd__mux2_1 _08487_ (.A0(\addroundkey_data_o[83] ),
    .A1(\fifo_bank_register.data_out[83] ),
    .S(_04556_),
    .X(_04561_));
 sky130_fd_sc_hd__clkbuf_1 _08488_ (.A(_04561_),
    .X(net369));
 sky130_fd_sc_hd__mux2_4 _08489_ (.A0(\addroundkey_data_o[84] ),
    .A1(\fifo_bank_register.data_out[84] ),
    .S(_04556_),
    .X(_04562_));
 sky130_fd_sc_hd__clkbuf_1 _08490_ (.A(_04562_),
    .X(net370));
 sky130_fd_sc_hd__mux2_1 _08491_ (.A0(\addroundkey_data_o[85] ),
    .A1(\fifo_bank_register.data_out[85] ),
    .S(_04556_),
    .X(_04563_));
 sky130_fd_sc_hd__clkbuf_1 _08492_ (.A(_04563_),
    .X(net371));
 sky130_fd_sc_hd__mux2_2 _08493_ (.A0(\addroundkey_data_o[86] ),
    .A1(\fifo_bank_register.data_out[86] ),
    .S(_04556_),
    .X(_04564_));
 sky130_fd_sc_hd__clkbuf_1 _08494_ (.A(_04564_),
    .X(net372));
 sky130_fd_sc_hd__mux2_2 _08495_ (.A0(\addroundkey_data_o[87] ),
    .A1(\fifo_bank_register.data_out[87] ),
    .S(_04556_),
    .X(_04565_));
 sky130_fd_sc_hd__buf_1 _08496_ (.A(_04565_),
    .X(net373));
 sky130_fd_sc_hd__mux2_2 _08497_ (.A0(\addroundkey_data_o[88] ),
    .A1(\fifo_bank_register.data_out[88] ),
    .S(_04556_),
    .X(_04566_));
 sky130_fd_sc_hd__clkbuf_1 _08498_ (.A(_04566_),
    .X(net374));
 sky130_fd_sc_hd__buf_6 _08499_ (.A(_04478_),
    .X(_04567_));
 sky130_fd_sc_hd__mux2_2 _08500_ (.A0(\addroundkey_data_o[89] ),
    .A1(\fifo_bank_register.data_out[89] ),
    .S(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__clkbuf_2 _08501_ (.A(_04568_),
    .X(net375));
 sky130_fd_sc_hd__mux2_1 _08502_ (.A0(\addroundkey_data_o[90] ),
    .A1(\fifo_bank_register.data_out[90] ),
    .S(_04567_),
    .X(_04569_));
 sky130_fd_sc_hd__clkbuf_1 _08503_ (.A(_04569_),
    .X(net377));
 sky130_fd_sc_hd__mux2_4 _08504_ (.A0(\addroundkey_data_o[91] ),
    .A1(\fifo_bank_register.data_out[91] ),
    .S(_04567_),
    .X(_04570_));
 sky130_fd_sc_hd__clkbuf_1 _08505_ (.A(_04570_),
    .X(net378));
 sky130_fd_sc_hd__mux2_8 _08506_ (.A0(\addroundkey_data_o[92] ),
    .A1(\fifo_bank_register.data_out[92] ),
    .S(_04567_),
    .X(_04571_));
 sky130_fd_sc_hd__clkbuf_1 _08507_ (.A(_04571_),
    .X(net379));
 sky130_fd_sc_hd__mux2_4 _08508_ (.A0(\addroundkey_data_o[93] ),
    .A1(\fifo_bank_register.data_out[93] ),
    .S(_04567_),
    .X(_04572_));
 sky130_fd_sc_hd__clkbuf_1 _08509_ (.A(_04572_),
    .X(net380));
 sky130_fd_sc_hd__mux2_4 _08510_ (.A0(\addroundkey_data_o[94] ),
    .A1(\fifo_bank_register.data_out[94] ),
    .S(_04567_),
    .X(_04573_));
 sky130_fd_sc_hd__clkbuf_1 _08511_ (.A(_04573_),
    .X(net381));
 sky130_fd_sc_hd__mux2_1 _08512_ (.A0(\addroundkey_data_o[95] ),
    .A1(\fifo_bank_register.data_out[95] ),
    .S(_04567_),
    .X(_04574_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _08513_ (.A(_04574_),
    .X(net382));
 sky130_fd_sc_hd__mux2_2 _08514_ (.A0(\addroundkey_data_o[96] ),
    .A1(\fifo_bank_register.data_out[96] ),
    .S(_04567_),
    .X(_04575_));
 sky130_fd_sc_hd__clkbuf_1 _08515_ (.A(_04575_),
    .X(net383));
 sky130_fd_sc_hd__mux2_1 _08516_ (.A0(\addroundkey_data_o[97] ),
    .A1(\fifo_bank_register.data_out[97] ),
    .S(_04567_),
    .X(_04576_));
 sky130_fd_sc_hd__clkbuf_2 _08517_ (.A(_04576_),
    .X(net384));
 sky130_fd_sc_hd__mux2_4 _08518_ (.A0(\addroundkey_data_o[98] ),
    .A1(\fifo_bank_register.data_out[98] ),
    .S(_04567_),
    .X(_04577_));
 sky130_fd_sc_hd__buf_2 _08519_ (.A(_04577_),
    .X(net385));
 sky130_fd_sc_hd__buf_6 _08520_ (.A(_04478_),
    .X(_04578_));
 sky130_fd_sc_hd__mux2_2 _08521_ (.A0(\addroundkey_data_o[99] ),
    .A1(\fifo_bank_register.data_out[99] ),
    .S(_04578_),
    .X(_04579_));
 sky130_fd_sc_hd__clkbuf_1 _08522_ (.A(_04579_),
    .X(net386));
 sky130_fd_sc_hd__mux2_2 _08523_ (.A0(\addroundkey_data_o[100] ),
    .A1(\fifo_bank_register.data_out[100] ),
    .S(_04578_),
    .X(_04580_));
 sky130_fd_sc_hd__buf_1 _08524_ (.A(_04580_),
    .X(net261));
 sky130_fd_sc_hd__mux2_1 _08525_ (.A0(\addroundkey_data_o[101] ),
    .A1(\fifo_bank_register.data_out[101] ),
    .S(_04578_),
    .X(_04581_));
 sky130_fd_sc_hd__clkbuf_2 _08526_ (.A(_04581_),
    .X(net262));
 sky130_fd_sc_hd__mux2_2 _08527_ (.A0(\addroundkey_data_o[102] ),
    .A1(\fifo_bank_register.data_out[102] ),
    .S(_04578_),
    .X(_04582_));
 sky130_fd_sc_hd__clkbuf_1 _08528_ (.A(_04582_),
    .X(net263));
 sky130_fd_sc_hd__mux2_2 _08529_ (.A0(\addroundkey_data_o[103] ),
    .A1(\fifo_bank_register.data_out[103] ),
    .S(_04578_),
    .X(_04583_));
 sky130_fd_sc_hd__clkbuf_1 _08530_ (.A(_04583_),
    .X(net264));
 sky130_fd_sc_hd__mux2_1 _08531_ (.A0(\addroundkey_data_o[104] ),
    .A1(\fifo_bank_register.data_out[104] ),
    .S(_04578_),
    .X(_04584_));
 sky130_fd_sc_hd__clkbuf_4 _08532_ (.A(_04584_),
    .X(net265));
 sky130_fd_sc_hd__mux2_1 _08533_ (.A0(\addroundkey_data_o[105] ),
    .A1(\fifo_bank_register.data_out[105] ),
    .S(_04578_),
    .X(_04585_));
 sky130_fd_sc_hd__clkbuf_4 _08534_ (.A(_04585_),
    .X(net266));
 sky130_fd_sc_hd__mux2_1 _08535_ (.A0(\addroundkey_data_o[106] ),
    .A1(\fifo_bank_register.data_out[106] ),
    .S(_04578_),
    .X(_04586_));
 sky130_fd_sc_hd__clkbuf_1 _08536_ (.A(_04586_),
    .X(net267));
 sky130_fd_sc_hd__mux2_2 _08537_ (.A0(\addroundkey_data_o[107] ),
    .A1(\fifo_bank_register.data_out[107] ),
    .S(_04578_),
    .X(_04587_));
 sky130_fd_sc_hd__clkbuf_1 _08538_ (.A(_04587_),
    .X(net268));
 sky130_fd_sc_hd__mux2_2 _08539_ (.A0(\addroundkey_data_o[108] ),
    .A1(\fifo_bank_register.data_out[108] ),
    .S(_04578_),
    .X(_04588_));
 sky130_fd_sc_hd__clkbuf_1 _08540_ (.A(_04588_),
    .X(net269));
 sky130_fd_sc_hd__buf_8 _08541_ (.A(_04466_),
    .X(_04589_));
 sky130_fd_sc_hd__mux2_2 _08542_ (.A0(\addroundkey_data_o[109] ),
    .A1(\fifo_bank_register.data_out[109] ),
    .S(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__buf_1 _08543_ (.A(_04590_),
    .X(net270));
 sky130_fd_sc_hd__mux2_4 _08544_ (.A0(\addroundkey_data_o[110] ),
    .A1(\fifo_bank_register.data_out[110] ),
    .S(_04589_),
    .X(_04591_));
 sky130_fd_sc_hd__clkbuf_1 _08545_ (.A(_04591_),
    .X(net272));
 sky130_fd_sc_hd__mux2_1 _08546_ (.A0(\addroundkey_data_o[111] ),
    .A1(\fifo_bank_register.data_out[111] ),
    .S(_04589_),
    .X(_04592_));
 sky130_fd_sc_hd__clkbuf_2 _08547_ (.A(_04592_),
    .X(net273));
 sky130_fd_sc_hd__mux2_4 _08548_ (.A0(\addroundkey_data_o[112] ),
    .A1(\fifo_bank_register.data_out[112] ),
    .S(_04589_),
    .X(_04593_));
 sky130_fd_sc_hd__clkbuf_1 _08549_ (.A(_04593_),
    .X(net274));
 sky130_fd_sc_hd__mux2_2 _08550_ (.A0(\addroundkey_data_o[113] ),
    .A1(\fifo_bank_register.data_out[113] ),
    .S(_04589_),
    .X(_04594_));
 sky130_fd_sc_hd__clkbuf_1 _08551_ (.A(_04594_),
    .X(net275));
 sky130_fd_sc_hd__mux2_1 _08552_ (.A0(\addroundkey_data_o[114] ),
    .A1(\fifo_bank_register.data_out[114] ),
    .S(_04589_),
    .X(_04595_));
 sky130_fd_sc_hd__clkbuf_2 _08553_ (.A(_04595_),
    .X(net276));
 sky130_fd_sc_hd__mux2_4 _08554_ (.A0(\addroundkey_data_o[115] ),
    .A1(\fifo_bank_register.data_out[115] ),
    .S(_04589_),
    .X(_04596_));
 sky130_fd_sc_hd__clkbuf_1 _08555_ (.A(_04596_),
    .X(net277));
 sky130_fd_sc_hd__mux2_2 _08556_ (.A0(\addroundkey_data_o[116] ),
    .A1(\fifo_bank_register.data_out[116] ),
    .S(_04589_),
    .X(_04597_));
 sky130_fd_sc_hd__buf_1 _08557_ (.A(_04597_),
    .X(net278));
 sky130_fd_sc_hd__mux2_4 _08558_ (.A0(\addroundkey_data_o[117] ),
    .A1(\fifo_bank_register.data_out[117] ),
    .S(_04589_),
    .X(_04598_));
 sky130_fd_sc_hd__clkbuf_1 _08559_ (.A(_04598_),
    .X(net279));
 sky130_fd_sc_hd__mux2_1 _08560_ (.A0(\addroundkey_data_o[118] ),
    .A1(\fifo_bank_register.data_out[118] ),
    .S(_04589_),
    .X(_04599_));
 sky130_fd_sc_hd__buf_2 _08561_ (.A(_04599_),
    .X(net280));
 sky130_fd_sc_hd__mux2_2 _08562_ (.A0(\addroundkey_data_o[119] ),
    .A1(\fifo_bank_register.data_out[119] ),
    .S(_04467_),
    .X(_04600_));
 sky130_fd_sc_hd__buf_1 _08563_ (.A(_04600_),
    .X(net281));
 sky130_fd_sc_hd__mux2_4 _08564_ (.A0(\addroundkey_data_o[120] ),
    .A1(\fifo_bank_register.data_out[120] ),
    .S(_04467_),
    .X(_04601_));
 sky130_fd_sc_hd__clkbuf_1 _08565_ (.A(_04601_),
    .X(net283));
 sky130_fd_sc_hd__mux2_1 _08566_ (.A0(\addroundkey_data_o[121] ),
    .A1(\fifo_bank_register.data_out[121] ),
    .S(_04467_),
    .X(_04602_));
 sky130_fd_sc_hd__buf_1 _08567_ (.A(_04602_),
    .X(net284));
 sky130_fd_sc_hd__mux2_1 _08568_ (.A0(\addroundkey_data_o[122] ),
    .A1(\fifo_bank_register.data_out[122] ),
    .S(_04467_),
    .X(_04603_));
 sky130_fd_sc_hd__clkbuf_2 _08569_ (.A(_04603_),
    .X(net285));
 sky130_fd_sc_hd__mux2_1 _08570_ (.A0(\addroundkey_data_o[123] ),
    .A1(\fifo_bank_register.data_out[123] ),
    .S(_04467_),
    .X(_04604_));
 sky130_fd_sc_hd__buf_1 _08571_ (.A(_04604_),
    .X(net286));
 sky130_fd_sc_hd__mux2_2 _08572_ (.A0(\addroundkey_data_o[124] ),
    .A1(\fifo_bank_register.data_out[124] ),
    .S(_04467_),
    .X(_04605_));
 sky130_fd_sc_hd__clkbuf_2 _08573_ (.A(_04605_),
    .X(net287));
 sky130_fd_sc_hd__mux2_2 _08574_ (.A0(\addroundkey_data_o[125] ),
    .A1(\fifo_bank_register.data_out[125] ),
    .S(_04467_),
    .X(_04606_));
 sky130_fd_sc_hd__clkbuf_2 _08575_ (.A(_04606_),
    .X(net288));
 sky130_fd_sc_hd__mux2_2 _08576_ (.A0(\addroundkey_data_o[126] ),
    .A1(\fifo_bank_register.data_out[126] ),
    .S(_04467_),
    .X(_04607_));
 sky130_fd_sc_hd__clkbuf_1 _08577_ (.A(_04607_),
    .X(net289));
 sky130_fd_sc_hd__mux2_2 _08578_ (.A0(\addroundkey_data_o[127] ),
    .A1(\fifo_bank_register.data_out[127] ),
    .S(_04467_),
    .X(_04608_));
 sky130_fd_sc_hd__clkbuf_1 _08579_ (.A(_04608_),
    .X(net290));
 sky130_fd_sc_hd__buf_4 _08580_ (.A(state),
    .X(_04609_));
 sky130_fd_sc_hd__clkinv_4 _08581_ (.A(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__clkbuf_4 _08582_ (.A(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__and2_1 _08583_ (.A(_04611_),
    .B(net258),
    .X(_04612_));
 sky130_fd_sc_hd__clkbuf_1 _08584_ (.A(_04612_),
    .X(next_first_round_reg));
 sky130_fd_sc_hd__buf_2 _08585_ (.A(\round[0] ),
    .X(_04613_));
 sky130_fd_sc_hd__or3_2 _08586_ (.A(\round[1] ),
    .B(_04613_),
    .C(\round[2] ),
    .X(_04614_));
 sky130_fd_sc_hd__nor2_1 _08587_ (.A(\round[3] ),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__and4bb_2 _08588_ (.A_N(_04613_),
    .B_N(\round[2] ),
    .C(\round[3] ),
    .D(\round[1] ),
    .X(_04616_));
 sky130_fd_sc_hd__inv_4 _08589_ (.A(net129),
    .Y(_04617_));
 sky130_fd_sc_hd__mux2_4 _08590_ (.A0(_04615_),
    .A1(_04616_),
    .S(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__a21oi_2 _08591_ (.A1(addroundkey_ready_o),
    .A2(_04618_),
    .B1(_04611_),
    .Y(_04619_));
 sky130_fd_sc_hd__or2_1 _08592_ (.A(next_first_round_reg),
    .B(_04619_),
    .X(_04620_));
 sky130_fd_sc_hd__clkbuf_1 _08593_ (.A(_04620_),
    .X(next_state));
 sky130_fd_sc_hd__and4bb_1 _08594_ (.A_N(\round[1] ),
    .B_N(\round[2] ),
    .C(\round[3] ),
    .D(_04613_),
    .X(_04621_));
 sky130_fd_sc_hd__mux2_1 _08595_ (.A0(_04615_),
    .A1(_04621_),
    .S(_04617_),
    .X(_04622_));
 sky130_fd_sc_hd__inv_2 _08596_ (.A(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__clkbuf_8 _08597_ (.A(net129),
    .X(_04624_));
 sky130_fd_sc_hd__nand2_2 _08598_ (.A(_04624_),
    .B(\sub1.ready_o ),
    .Y(_04625_));
 sky130_fd_sc_hd__nand2_4 _08599_ (.A(_04617_),
    .B(\mix1.ready_o ),
    .Y(_04626_));
 sky130_fd_sc_hd__nand2_2 _08600_ (.A(_04625_),
    .B(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__or2_1 _08601_ (.A(first_round_reg),
    .B(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__and2_2 _08602_ (.A(\sub1.ready_o ),
    .B(_04622_),
    .X(_04629_));
 sky130_fd_sc_hd__a21o_1 _08603_ (.A1(_04623_),
    .A2(_04628_),
    .B1(_04629_),
    .X(_04630_));
 sky130_fd_sc_hd__a22o_1 _08604_ (.A1(_04611_),
    .A2(net671),
    .B1(_04619_),
    .B2(_04630_),
    .X(next_addroundkey_start_i));
 sky130_fd_sc_hd__or2_1 _08605_ (.A(net258),
    .B(_04468_),
    .X(_04631_));
 sky130_fd_sc_hd__clkbuf_2 _08606_ (.A(_04631_),
    .X(\fifo_bank_register.clk ));
 sky130_fd_sc_hd__xor2_1 _08607_ (.A(\round[1] ),
    .B(\addroundkey_round[1] ),
    .X(_04632_));
 sky130_fd_sc_hd__xor2_1 _08608_ (.A(\round[0] ),
    .B(\addroundkey_round[0] ),
    .X(_04633_));
 sky130_fd_sc_hd__xor2_1 _08609_ (.A(\round[3] ),
    .B(\addroundkey_round[3] ),
    .X(_04634_));
 sky130_fd_sc_hd__xor2_1 _08610_ (.A(\round[2] ),
    .B(\addroundkey_round[2] ),
    .X(_04635_));
 sky130_fd_sc_hd__or4_2 _08611_ (.A(_04632_),
    .B(_04633_),
    .C(_04634_),
    .D(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__nand2b_2 _08612_ (.A_N(addroundkey_start_i),
    .B(\ks1.ready_o ),
    .Y(_04637_));
 sky130_fd_sc_hd__nand2_2 _08613_ (.A(addroundkey_start_i),
    .B(_04615_),
    .Y(_04638_));
 sky130_fd_sc_hd__clkbuf_8 _08614_ (.A(_04638_),
    .X(_04639_));
 sky130_fd_sc_hd__o21ai_2 _08615_ (.A1(_04636_),
    .A2(_04637_),
    .B1(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__buf_4 _08616_ (.A(_04640_),
    .X(next_addroundkey_ready_o));
 sky130_fd_sc_hd__or2_2 _08617_ (.A(\round[3] ),
    .B(_04614_),
    .X(_04641_));
 sky130_fd_sc_hd__nand2_4 _08618_ (.A(addroundkey_start_i),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__or2b_1 _08619_ (.A(_04637_),
    .B_N(_04636_),
    .X(_04643_));
 sky130_fd_sc_hd__clkbuf_4 _08620_ (.A(_04643_),
    .X(_04644_));
 sky130_fd_sc_hd__a2111o_1 _08621_ (.A1(_04642_),
    .A2(_04644_),
    .B1(\ks1.state[1] ),
    .C1(\ks1.state[0] ),
    .D1(\ks1.state[2] ),
    .X(_04645_));
 sky130_fd_sc_hd__or2_1 _08622_ (.A(\ks1.state[2] ),
    .B(_04370_),
    .X(_04646_));
 sky130_fd_sc_hd__and3_1 _08623_ (.A(_04371_),
    .B(_04645_),
    .C(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__buf_4 _08624_ (.A(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__nand2_4 _08625_ (.A(_04624_),
    .B(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__or2_4 _08626_ (.A(_04617_),
    .B(_04616_),
    .X(_04650_));
 sky130_fd_sc_hd__a22oi_2 _08627_ (.A1(net129),
    .A2(\mix1.ready_o ),
    .B1(_04650_),
    .B2(addroundkey_ready_o),
    .Y(_04651_));
 sky130_fd_sc_hd__a21oi_4 _08628_ (.A1(state),
    .A2(_04618_),
    .B1(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__and3b_4 _08629_ (.A_N(\sub1.state[4] ),
    .B(_04366_),
    .C(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__nor2_1 _08630_ (.A(_04617_),
    .B(_04616_),
    .Y(_04654_));
 sky130_fd_sc_hd__clkbuf_4 _08631_ (.A(_04654_),
    .X(_04655_));
 sky130_fd_sc_hd__buf_4 _08632_ (.A(_04655_),
    .X(_04656_));
 sky130_fd_sc_hd__buf_4 _08633_ (.A(_04656_),
    .X(_04657_));
 sky130_fd_sc_hd__buf_4 _08634_ (.A(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__mux2_1 _08635_ (.A0(\addroundkey_data_o[124] ),
    .A1(\mix1.data_o[124] ),
    .S(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__and4b_1 _08636_ (.A_N(\sub1.state[1] ),
    .B(_04363_),
    .C(\sub1.state[3] ),
    .D(\sub1.state[2] ),
    .X(_04660_));
 sky130_fd_sc_hd__clkbuf_4 _08637_ (.A(_04660_),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_4 _08638_ (.A(_04654_),
    .X(_04662_));
 sky130_fd_sc_hd__buf_4 _08639_ (.A(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__mux2_1 _08640_ (.A0(\addroundkey_data_o[20] ),
    .A1(\mix1.data_o[20] ),
    .S(_04663_),
    .X(_04664_));
 sky130_fd_sc_hd__buf_4 _08641_ (.A(_04655_),
    .X(_04665_));
 sky130_fd_sc_hd__buf_4 _08642_ (.A(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__mux2_1 _08643_ (.A0(\addroundkey_data_o[76] ),
    .A1(\mix1.data_o[76] ),
    .S(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__and4bb_4 _08644_ (.A_N(_04363_),
    .B_N(_04364_),
    .C(_04365_),
    .D(_04362_),
    .X(_04668_));
 sky130_fd_sc_hd__a22o_1 _08645_ (.A1(_04661_),
    .A2(_04664_),
    .B1(_04667_),
    .B2(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__and4bb_4 _08646_ (.A_N(\sub1.state[1] ),
    .B_N(\sub1.state[2] ),
    .C(\sub1.state[3] ),
    .D(_04363_),
    .X(_04670_));
 sky130_fd_sc_hd__mux2_1 _08647_ (.A0(\addroundkey_data_o[52] ),
    .A1(\mix1.data_o[52] ),
    .S(_04663_),
    .X(_04671_));
 sky130_fd_sc_hd__mux2_1 _08648_ (.A0(\addroundkey_data_o[28] ),
    .A1(\mix1.data_o[28] ),
    .S(_04666_),
    .X(_04672_));
 sky130_fd_sc_hd__inv_2 _08649_ (.A(\sub1.state[0] ),
    .Y(_04673_));
 sky130_fd_sc_hd__and4b_1 _08650_ (.A_N(\sub1.state[1] ),
    .B(_04673_),
    .C(\sub1.state[3] ),
    .D(\sub1.state[2] ),
    .X(_04674_));
 sky130_fd_sc_hd__clkbuf_4 _08651_ (.A(_04674_),
    .X(_04675_));
 sky130_fd_sc_hd__a22o_1 _08652_ (.A1(_04670_),
    .A2(_04671_),
    .B1(_04672_),
    .B2(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__and4bb_4 _08653_ (.A_N(_04362_),
    .B_N(_04364_),
    .C(_04365_),
    .D(_04363_),
    .X(_04677_));
 sky130_fd_sc_hd__mux2_1 _08654_ (.A0(\addroundkey_data_o[84] ),
    .A1(\mix1.data_o[84] ),
    .S(_04663_),
    .X(_04678_));
 sky130_fd_sc_hd__mux2_1 _08655_ (.A0(\addroundkey_data_o[116] ),
    .A1(\mix1.data_o[116] ),
    .S(_04666_),
    .X(_04679_));
 sky130_fd_sc_hd__or2_1 _08656_ (.A(\sub1.state[1] ),
    .B(_04673_),
    .X(_04680_));
 sky130_fd_sc_hd__or2_2 _08657_ (.A(\sub1.state[3] ),
    .B(\sub1.state[2] ),
    .X(_04681_));
 sky130_fd_sc_hd__nor2_2 _08658_ (.A(_04680_),
    .B(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__a22o_1 _08659_ (.A1(_04677_),
    .A2(_04678_),
    .B1(_04679_),
    .B2(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__nor4b_4 _08660_ (.A(_04362_),
    .B(_04363_),
    .C(_04365_),
    .D_N(_04364_),
    .Y(_04684_));
 sky130_fd_sc_hd__mux2_1 _08661_ (.A0(\addroundkey_data_o[60] ),
    .A1(\mix1.data_o[60] ),
    .S(_04663_),
    .X(_04685_));
 sky130_fd_sc_hd__mux2_1 _08662_ (.A0(\addroundkey_data_o[4] ),
    .A1(\mix1.data_o[4] ),
    .S(_04666_),
    .X(_04686_));
 sky130_fd_sc_hd__and2_1 _08663_ (.A(\sub1.state[1] ),
    .B(\sub1.state[0] ),
    .X(_04687_));
 sky130_fd_sc_hd__and3_1 _08664_ (.A(_04364_),
    .B(_04365_),
    .C(_04687_),
    .X(_04688_));
 sky130_fd_sc_hd__clkbuf_4 _08665_ (.A(_04688_),
    .X(_04689_));
 sky130_fd_sc_hd__a22o_1 _08666_ (.A1(_04684_),
    .A2(_04685_),
    .B1(_04686_),
    .B2(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__or4_1 _08667_ (.A(_04669_),
    .B(_04676_),
    .C(_04683_),
    .D(_04690_),
    .X(_04691_));
 sky130_fd_sc_hd__and4bb_2 _08668_ (.A_N(_04363_),
    .B_N(\sub1.state[2] ),
    .C(\sub1.state[3] ),
    .D(_04362_),
    .X(_04692_));
 sky130_fd_sc_hd__clkbuf_4 _08669_ (.A(_04692_),
    .X(_04693_));
 sky130_fd_sc_hd__and3b_2 _08670_ (.A_N(\sub1.state[2] ),
    .B(_04687_),
    .C(_04364_),
    .X(_04694_));
 sky130_fd_sc_hd__clkbuf_4 _08671_ (.A(_04694_),
    .X(_04695_));
 sky130_fd_sc_hd__a22o_1 _08672_ (.A1(\mix1.data_o[44] ),
    .A2(_04693_),
    .B1(_04695_),
    .B2(\mix1.data_o[36] ),
    .X(_04696_));
 sky130_fd_sc_hd__a22o_1 _08673_ (.A1(\addroundkey_data_o[44] ),
    .A2(_04693_),
    .B1(_04695_),
    .B2(\addroundkey_data_o[36] ),
    .X(_04697_));
 sky130_fd_sc_hd__clkbuf_4 _08674_ (.A(_04650_),
    .X(_04698_));
 sky130_fd_sc_hd__mux2_1 _08675_ (.A0(_04696_),
    .A1(_04697_),
    .S(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__nand2_2 _08676_ (.A(_04362_),
    .B(_04363_),
    .Y(_04700_));
 sky130_fd_sc_hd__nor2_4 _08677_ (.A(_04700_),
    .B(_04681_),
    .Y(_04701_));
 sky130_fd_sc_hd__buf_4 _08678_ (.A(_04656_),
    .X(_04702_));
 sky130_fd_sc_hd__or2_1 _08679_ (.A(\addroundkey_data_o[100] ),
    .B(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__o211a_1 _08680_ (.A1(\mix1.data_o[100] ),
    .A2(_04698_),
    .B1(_04701_),
    .C1(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__nand2_1 _08681_ (.A(_04362_),
    .B(_04673_),
    .Y(_04705_));
 sky130_fd_sc_hd__nor2_4 _08682_ (.A(_04705_),
    .B(_04681_),
    .Y(_04706_));
 sky130_fd_sc_hd__mux2_1 _08683_ (.A0(\addroundkey_data_o[108] ),
    .A1(\mix1.data_o[108] ),
    .S(_04663_),
    .X(_04707_));
 sky130_fd_sc_hd__mux2_1 _08684_ (.A0(\addroundkey_data_o[12] ),
    .A1(\mix1.data_o[12] ),
    .S(_04666_),
    .X(_04708_));
 sky130_fd_sc_hd__and4_1 _08685_ (.A(_04362_),
    .B(_04673_),
    .C(_04364_),
    .D(_04365_),
    .X(_04709_));
 sky130_fd_sc_hd__buf_2 _08686_ (.A(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__a22o_1 _08687_ (.A1(_04706_),
    .A2(_04707_),
    .B1(_04708_),
    .B2(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__and3b_1 _08688_ (.A_N(\sub1.state[3] ),
    .B(\sub1.state[2] ),
    .C(_04687_),
    .X(_04712_));
 sky130_fd_sc_hd__clkbuf_4 _08689_ (.A(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__mux2_1 _08690_ (.A0(\addroundkey_data_o[68] ),
    .A1(\mix1.data_o[68] ),
    .S(_04663_),
    .X(_04714_));
 sky130_fd_sc_hd__mux2_1 _08691_ (.A0(\addroundkey_data_o[92] ),
    .A1(\mix1.data_o[92] ),
    .S(_04666_),
    .X(_04715_));
 sky130_fd_sc_hd__nor4b_4 _08692_ (.A(_04362_),
    .B(_04363_),
    .C(_04364_),
    .D_N(_04365_),
    .Y(_04716_));
 sky130_fd_sc_hd__a22o_1 _08693_ (.A1(_04713_),
    .A2(_04714_),
    .B1(_04715_),
    .B2(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__or4_1 _08694_ (.A(_04699_),
    .B(_04704_),
    .C(_04711_),
    .D(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__a211o_1 _08695_ (.A1(_04653_),
    .A2(_04659_),
    .B1(_04691_),
    .C1(_04718_),
    .X(_04719_));
 sky130_fd_sc_hd__inv_2 _08696_ (.A(\ks1.state[2] ),
    .Y(_04720_));
 sky130_fd_sc_hd__nand3_2 _08697_ (.A(\ks1.state[1] ),
    .B(\ks1.state[0] ),
    .C(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nor3_1 _08698_ (.A(\addroundkey_round[1] ),
    .B(\addroundkey_round[2] ),
    .C(\addroundkey_round[3] ),
    .Y(_04722_));
 sky130_fd_sc_hd__and2_1 _08699_ (.A(addroundkey_start_i),
    .B(_04641_),
    .X(_04723_));
 sky130_fd_sc_hd__a21oi_1 _08700_ (.A1(_04644_),
    .A2(_04722_),
    .B1(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__clkbuf_4 _08701_ (.A(_04724_),
    .X(_04725_));
 sky130_fd_sc_hd__clkbuf_4 _08702_ (.A(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__nand2_1 _08703_ (.A(\ks1.ready_o ),
    .B(_04636_),
    .Y(_04727_));
 sky130_fd_sc_hd__and2_1 _08704_ (.A(_04722_),
    .B(_04727_),
    .X(_04728_));
 sky130_fd_sc_hd__clkbuf_4 _08705_ (.A(_04728_),
    .X(_04729_));
 sky130_fd_sc_hd__buf_2 _08706_ (.A(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__o21a_4 _08707_ (.A1(_04641_),
    .A2(_04722_),
    .B1(addroundkey_start_i),
    .X(_04731_));
 sky130_fd_sc_hd__buf_2 _08708_ (.A(_04731_),
    .X(_04732_));
 sky130_fd_sc_hd__o31a_1 _08709_ (.A1(\ks1.key_reg[4] ),
    .A2(_04730_),
    .A3(_04732_),
    .B1(net202),
    .X(_04733_));
 sky130_fd_sc_hd__a21oi_1 _08710_ (.A1(\ks1.key_reg[4] ),
    .A2(_04726_),
    .B1(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__buf_4 _08711_ (.A(_04724_),
    .X(_04735_));
 sky130_fd_sc_hd__mux2_1 _08712_ (.A0(net161),
    .A1(\ks1.key_reg[12] ),
    .S(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__nor2_1 _08713_ (.A(\ks1.state[0] ),
    .B(\ks1.state[2] ),
    .Y(_04737_));
 sky130_fd_sc_hd__and2_1 _08714_ (.A(\ks1.state[1] ),
    .B(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__a2bb2o_1 _08715_ (.A1_N(_04721_),
    .A2_N(_04734_),
    .B1(_04736_),
    .B2(_04738_),
    .X(_04739_));
 sky130_fd_sc_hd__or3b_1 _08716_ (.A(\ks1.state[1] ),
    .B(\ks1.state[2] ),
    .C_N(\ks1.state[0] ),
    .X(_04740_));
 sky130_fd_sc_hd__buf_2 _08717_ (.A(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__buf_4 _08718_ (.A(_04735_),
    .X(_04742_));
 sky130_fd_sc_hd__o31a_1 _08719_ (.A1(\ks1.key_reg[20] ),
    .A2(_04730_),
    .A3(_04732_),
    .B1(net170),
    .X(_04743_));
 sky130_fd_sc_hd__a21oi_1 _08720_ (.A1(\ks1.key_reg[20] ),
    .A2(_04742_),
    .B1(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__clkbuf_4 _08721_ (.A(_04729_),
    .X(_04745_));
 sky130_fd_sc_hd__buf_2 _08722_ (.A(_04731_),
    .X(_04746_));
 sky130_fd_sc_hd__or3_1 _08723_ (.A(\ks1.key_reg[28] ),
    .B(_04745_),
    .C(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__a22o_1 _08724_ (.A1(\ks1.key_reg[28] ),
    .A2(_04735_),
    .B1(_04747_),
    .B2(net178),
    .X(_04748_));
 sky130_fd_sc_hd__inv_2 _08725_ (.A(_04644_),
    .Y(_04749_));
 sky130_fd_sc_hd__o211a_1 _08726_ (.A1(_04723_),
    .A2(_04749_),
    .B1(_04720_),
    .C1(_04370_),
    .X(_04750_));
 sky130_fd_sc_hd__a2bb2o_1 _08727_ (.A1_N(_04741_),
    .A2_N(_04744_),
    .B1(_04748_),
    .B2(_04750_),
    .X(_04751_));
 sky130_fd_sc_hd__a211o_2 _08728_ (.A1(_04648_),
    .A2(_04719_),
    .B1(_04739_),
    .C1(_04751_),
    .X(_04752_));
 sky130_fd_sc_hd__o31a_1 _08729_ (.A1(\ks1.key_reg[17] ),
    .A2(_04730_),
    .A3(_04732_),
    .B1(net166),
    .X(_04753_));
 sky130_fd_sc_hd__a21oi_1 _08730_ (.A1(\ks1.key_reg[17] ),
    .A2(_04742_),
    .B1(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__nand2_2 _08731_ (.A(\ks1.state[1] ),
    .B(_04737_),
    .Y(_04755_));
 sky130_fd_sc_hd__o31a_1 _08732_ (.A1(\ks1.key_reg[9] ),
    .A2(_04730_),
    .A3(_04732_),
    .B1(net257),
    .X(_04756_));
 sky130_fd_sc_hd__a21oi_2 _08733_ (.A1(\ks1.key_reg[9] ),
    .A2(_04742_),
    .B1(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__o31a_1 _08734_ (.A1(\ks1.key_reg[1] ),
    .A2(_04730_),
    .A3(_04732_),
    .B1(net169),
    .X(_04758_));
 sky130_fd_sc_hd__a21oi_1 _08735_ (.A1(\ks1.key_reg[1] ),
    .A2(_04726_),
    .B1(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__o31a_1 _08736_ (.A1(\ks1.key_reg[25] ),
    .A2(_04730_),
    .A3(_04732_),
    .B1(net175),
    .X(_04760_));
 sky130_fd_sc_hd__a21oi_2 _08737_ (.A1(\ks1.key_reg[25] ),
    .A2(_04726_),
    .B1(_04760_),
    .Y(_04761_));
 sky130_fd_sc_hd__or2_1 _08738_ (.A(\mix1.data_o[121] ),
    .B(_04698_),
    .X(_04762_));
 sky130_fd_sc_hd__o211a_1 _08739_ (.A1(\addroundkey_data_o[121] ),
    .A2(_04658_),
    .B1(_04762_),
    .C1(_04653_),
    .X(_04763_));
 sky130_fd_sc_hd__mux2_1 _08740_ (.A0(\addroundkey_data_o[65] ),
    .A1(\mix1.data_o[65] ),
    .S(_04655_),
    .X(_04764_));
 sky130_fd_sc_hd__mux2_1 _08741_ (.A0(\addroundkey_data_o[73] ),
    .A1(\mix1.data_o[73] ),
    .S(_04655_),
    .X(_04765_));
 sky130_fd_sc_hd__a22o_1 _08742_ (.A1(_04713_),
    .A2(_04764_),
    .B1(_04668_),
    .B2(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__mux2_1 _08743_ (.A0(\addroundkey_data_o[113] ),
    .A1(\mix1.data_o[113] ),
    .S(_04655_),
    .X(_04767_));
 sky130_fd_sc_hd__mux2_1 _08744_ (.A0(\addroundkey_data_o[97] ),
    .A1(\mix1.data_o[97] ),
    .S(_04655_),
    .X(_04768_));
 sky130_fd_sc_hd__a22o_1 _08745_ (.A1(_04682_),
    .A2(_04767_),
    .B1(_04701_),
    .B2(_04768_),
    .X(_04769_));
 sky130_fd_sc_hd__mux2_1 _08746_ (.A0(\addroundkey_data_o[81] ),
    .A1(\mix1.data_o[81] ),
    .S(_04654_),
    .X(_04770_));
 sky130_fd_sc_hd__mux2_1 _08747_ (.A0(\addroundkey_data_o[105] ),
    .A1(\mix1.data_o[105] ),
    .S(_04655_),
    .X(_04771_));
 sky130_fd_sc_hd__a22o_1 _08748_ (.A1(_04677_),
    .A2(_04770_),
    .B1(_04706_),
    .B2(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__mux2_1 _08749_ (.A0(\addroundkey_data_o[17] ),
    .A1(\mix1.data_o[17] ),
    .S(_04655_),
    .X(_04773_));
 sky130_fd_sc_hd__a22o_1 _08750_ (.A1(\mix1.data_o[25] ),
    .A2(_04675_),
    .B1(_04670_),
    .B2(\mix1.data_o[49] ),
    .X(_04774_));
 sky130_fd_sc_hd__a22o_1 _08751_ (.A1(_04661_),
    .A2(_04773_),
    .B1(_04774_),
    .B2(_04656_),
    .X(_04775_));
 sky130_fd_sc_hd__or4_1 _08752_ (.A(_04766_),
    .B(_04769_),
    .C(_04772_),
    .D(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__buf_4 _08753_ (.A(_04693_),
    .X(_04777_));
 sky130_fd_sc_hd__buf_4 _08754_ (.A(_04662_),
    .X(_04778_));
 sky130_fd_sc_hd__mux2_1 _08755_ (.A0(\addroundkey_data_o[41] ),
    .A1(\mix1.data_o[41] ),
    .S(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__mux2_1 _08756_ (.A0(\addroundkey_data_o[1] ),
    .A1(\mix1.data_o[1] ),
    .S(_04662_),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_1 _08757_ (.A0(\addroundkey_data_o[89] ),
    .A1(\mix1.data_o[89] ),
    .S(_04662_),
    .X(_04781_));
 sky130_fd_sc_hd__a22o_1 _08758_ (.A1(_04689_),
    .A2(_04780_),
    .B1(_04716_),
    .B2(_04781_),
    .X(_04782_));
 sky130_fd_sc_hd__a21o_1 _08759_ (.A1(_04777_),
    .A2(_04779_),
    .B1(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__clkbuf_4 _08760_ (.A(_04695_),
    .X(_04784_));
 sky130_fd_sc_hd__mux2_1 _08761_ (.A0(\addroundkey_data_o[33] ),
    .A1(\mix1.data_o[33] ),
    .S(_04656_),
    .X(_04785_));
 sky130_fd_sc_hd__a22o_1 _08762_ (.A1(\addroundkey_data_o[25] ),
    .A2(_04675_),
    .B1(_04670_),
    .B2(\addroundkey_data_o[49] ),
    .X(_04786_));
 sky130_fd_sc_hd__a22o_1 _08763_ (.A1(_04784_),
    .A2(_04785_),
    .B1(_04786_),
    .B2(_04698_),
    .X(_04787_));
 sky130_fd_sc_hd__mux2_1 _08764_ (.A0(\addroundkey_data_o[9] ),
    .A1(\mix1.data_o[9] ),
    .S(_04656_),
    .X(_04788_));
 sky130_fd_sc_hd__mux2_1 _08765_ (.A0(\addroundkey_data_o[57] ),
    .A1(\mix1.data_o[57] ),
    .S(_04778_),
    .X(_04789_));
 sky130_fd_sc_hd__a22o_1 _08766_ (.A1(_04710_),
    .A2(_04788_),
    .B1(_04684_),
    .B2(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__or4_2 _08767_ (.A(_04776_),
    .B(_04783_),
    .C(_04787_),
    .D(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__o21ai_2 _08768_ (.A1(_04763_),
    .A2(_04791_),
    .B1(_04648_),
    .Y(_04792_));
 sky130_fd_sc_hd__o221a_1 _08769_ (.A1(_04721_),
    .A2(_04759_),
    .B1(_04761_),
    .B2(_04645_),
    .C1(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__o221a_2 _08770_ (.A1(_04741_),
    .A2(_04754_),
    .B1(_04755_),
    .B2(_04757_),
    .C1(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__o31a_1 _08771_ (.A1(\ks1.key_reg[19] ),
    .A2(_04730_),
    .A3(_04732_),
    .B1(net168),
    .X(_04795_));
 sky130_fd_sc_hd__a21oi_1 _08772_ (.A1(\ks1.key_reg[19] ),
    .A2(_04742_),
    .B1(_04795_),
    .Y(_04796_));
 sky130_fd_sc_hd__or3_1 _08773_ (.A(\ks1.key_reg[11] ),
    .B(_04745_),
    .C(_04746_),
    .X(_04797_));
 sky130_fd_sc_hd__a22o_1 _08774_ (.A1(\ks1.key_reg[11] ),
    .A2(_04735_),
    .B1(_04797_),
    .B2(net152),
    .X(_04798_));
 sky130_fd_sc_hd__o31a_1 _08775_ (.A1(\ks1.key_reg[3] ),
    .A2(_04730_),
    .A3(_04732_),
    .B1(net191),
    .X(_04799_));
 sky130_fd_sc_hd__a21oi_1 _08776_ (.A1(\ks1.key_reg[3] ),
    .A2(_04726_),
    .B1(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__o2bb2a_1 _08777_ (.A1_N(_04798_),
    .A2_N(_04738_),
    .B1(_04721_),
    .B2(_04800_),
    .X(_04801_));
 sky130_fd_sc_hd__mux2_1 _08778_ (.A0(\addroundkey_data_o[123] ),
    .A1(\mix1.data_o[123] ),
    .S(_04657_),
    .X(_04802_));
 sky130_fd_sc_hd__clkbuf_8 _08779_ (.A(_04655_),
    .X(_04803_));
 sky130_fd_sc_hd__mux2_1 _08780_ (.A0(\addroundkey_data_o[75] ),
    .A1(\mix1.data_o[75] ),
    .S(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__buf_4 _08781_ (.A(_04655_),
    .X(_04805_));
 sky130_fd_sc_hd__mux2_1 _08782_ (.A0(\addroundkey_data_o[91] ),
    .A1(\mix1.data_o[91] ),
    .S(_04805_),
    .X(_04806_));
 sky130_fd_sc_hd__a22o_1 _08783_ (.A1(_04668_),
    .A2(_04804_),
    .B1(_04806_),
    .B2(_04716_),
    .X(_04807_));
 sky130_fd_sc_hd__mux2_1 _08784_ (.A0(\addroundkey_data_o[107] ),
    .A1(\mix1.data_o[107] ),
    .S(_04803_),
    .X(_04808_));
 sky130_fd_sc_hd__mux2_1 _08785_ (.A0(\addroundkey_data_o[27] ),
    .A1(\mix1.data_o[27] ),
    .S(_04805_),
    .X(_04809_));
 sky130_fd_sc_hd__a22o_1 _08786_ (.A1(_04706_),
    .A2(_04808_),
    .B1(_04809_),
    .B2(_04675_),
    .X(_04810_));
 sky130_fd_sc_hd__mux2_1 _08787_ (.A0(\addroundkey_data_o[11] ),
    .A1(\mix1.data_o[11] ),
    .S(_04665_),
    .X(_04811_));
 sky130_fd_sc_hd__mux2_1 _08788_ (.A0(\addroundkey_data_o[59] ),
    .A1(\mix1.data_o[59] ),
    .S(_04805_),
    .X(_04812_));
 sky130_fd_sc_hd__a22o_1 _08789_ (.A1(_04710_),
    .A2(_04811_),
    .B1(_04812_),
    .B2(_04684_),
    .X(_04813_));
 sky130_fd_sc_hd__mux2_1 _08790_ (.A0(\addroundkey_data_o[51] ),
    .A1(\mix1.data_o[51] ),
    .S(_04803_),
    .X(_04814_));
 sky130_fd_sc_hd__mux2_1 _08791_ (.A0(\addroundkey_data_o[67] ),
    .A1(\mix1.data_o[67] ),
    .S(_04805_),
    .X(_04815_));
 sky130_fd_sc_hd__a22o_1 _08792_ (.A1(_04670_),
    .A2(_04814_),
    .B1(_04815_),
    .B2(_04713_),
    .X(_04816_));
 sky130_fd_sc_hd__or4_1 _08793_ (.A(_04807_),
    .B(_04810_),
    .C(_04813_),
    .D(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__a22o_1 _08794_ (.A1(\addroundkey_data_o[83] ),
    .A2(_04677_),
    .B1(_04661_),
    .B2(\addroundkey_data_o[19] ),
    .X(_04818_));
 sky130_fd_sc_hd__a22o_1 _08795_ (.A1(\mix1.data_o[83] ),
    .A2(_04677_),
    .B1(_04661_),
    .B2(\mix1.data_o[19] ),
    .X(_04819_));
 sky130_fd_sc_hd__mux2_1 _08796_ (.A0(_04818_),
    .A1(_04819_),
    .S(_04702_),
    .X(_04820_));
 sky130_fd_sc_hd__or2_1 _08797_ (.A(\addroundkey_data_o[43] ),
    .B(_04663_),
    .X(_04821_));
 sky130_fd_sc_hd__o211a_1 _08798_ (.A1(\mix1.data_o[43] ),
    .A2(_04698_),
    .B1(_04693_),
    .C1(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__mux2_1 _08799_ (.A0(\addroundkey_data_o[99] ),
    .A1(\mix1.data_o[99] ),
    .S(_04803_),
    .X(_04823_));
 sky130_fd_sc_hd__mux2_1 _08800_ (.A0(\addroundkey_data_o[115] ),
    .A1(\mix1.data_o[115] ),
    .S(_04656_),
    .X(_04824_));
 sky130_fd_sc_hd__a22o_1 _08801_ (.A1(_04701_),
    .A2(_04823_),
    .B1(_04824_),
    .B2(_04682_),
    .X(_04825_));
 sky130_fd_sc_hd__mux2_1 _08802_ (.A0(\addroundkey_data_o[35] ),
    .A1(\mix1.data_o[35] ),
    .S(_04805_),
    .X(_04826_));
 sky130_fd_sc_hd__mux2_1 _08803_ (.A0(\addroundkey_data_o[3] ),
    .A1(\mix1.data_o[3] ),
    .S(_04656_),
    .X(_04827_));
 sky130_fd_sc_hd__a22o_1 _08804_ (.A1(_04695_),
    .A2(_04826_),
    .B1(_04827_),
    .B2(_04689_),
    .X(_04828_));
 sky130_fd_sc_hd__or4_1 _08805_ (.A(_04820_),
    .B(_04822_),
    .C(_04825_),
    .D(_04828_),
    .X(_04829_));
 sky130_fd_sc_hd__a211o_2 _08806_ (.A1(_04653_),
    .A2(_04802_),
    .B1(_04817_),
    .C1(_04829_),
    .X(_04830_));
 sky130_fd_sc_hd__mux2_1 _08807_ (.A0(net177),
    .A1(\ks1.key_reg[27] ),
    .S(_04726_),
    .X(_04831_));
 sky130_fd_sc_hd__a22oi_1 _08808_ (.A1(_04648_),
    .A2(_04830_),
    .B1(_04831_),
    .B2(_04750_),
    .Y(_04832_));
 sky130_fd_sc_hd__o211a_1 _08809_ (.A1(_04741_),
    .A2(_04796_),
    .B1(_04801_),
    .C1(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__mux2_1 _08810_ (.A0(\addroundkey_data_o[126] ),
    .A1(\mix1.data_o[126] ),
    .S(_04657_),
    .X(_04834_));
 sky130_fd_sc_hd__mux2_1 _08811_ (.A0(\addroundkey_data_o[22] ),
    .A1(\mix1.data_o[22] ),
    .S(_04662_),
    .X(_04835_));
 sky130_fd_sc_hd__mux2_1 _08812_ (.A0(\addroundkey_data_o[78] ),
    .A1(\mix1.data_o[78] ),
    .S(_04803_),
    .X(_04836_));
 sky130_fd_sc_hd__a22o_1 _08813_ (.A1(_04661_),
    .A2(_04835_),
    .B1(_04836_),
    .B2(_04668_),
    .X(_04837_));
 sky130_fd_sc_hd__mux2_1 _08814_ (.A0(\addroundkey_data_o[54] ),
    .A1(\mix1.data_o[54] ),
    .S(_04662_),
    .X(_04838_));
 sky130_fd_sc_hd__mux2_1 _08815_ (.A0(\addroundkey_data_o[30] ),
    .A1(\mix1.data_o[30] ),
    .S(_04665_),
    .X(_04839_));
 sky130_fd_sc_hd__a22o_1 _08816_ (.A1(_04670_),
    .A2(_04838_),
    .B1(_04839_),
    .B2(_04675_),
    .X(_04840_));
 sky130_fd_sc_hd__mux2_1 _08817_ (.A0(\addroundkey_data_o[86] ),
    .A1(\mix1.data_o[86] ),
    .S(_04662_),
    .X(_04841_));
 sky130_fd_sc_hd__mux2_1 _08818_ (.A0(\addroundkey_data_o[118] ),
    .A1(\mix1.data_o[118] ),
    .S(_04665_),
    .X(_04842_));
 sky130_fd_sc_hd__a22o_1 _08819_ (.A1(_04677_),
    .A2(_04841_),
    .B1(_04842_),
    .B2(_04682_),
    .X(_04843_));
 sky130_fd_sc_hd__mux2_1 _08820_ (.A0(\addroundkey_data_o[62] ),
    .A1(\mix1.data_o[62] ),
    .S(_04662_),
    .X(_04844_));
 sky130_fd_sc_hd__mux2_1 _08821_ (.A0(\addroundkey_data_o[6] ),
    .A1(\mix1.data_o[6] ),
    .S(_04803_),
    .X(_04845_));
 sky130_fd_sc_hd__a22o_1 _08822_ (.A1(_04684_),
    .A2(_04844_),
    .B1(_04845_),
    .B2(_04689_),
    .X(_04846_));
 sky130_fd_sc_hd__or4_1 _08823_ (.A(_04837_),
    .B(_04840_),
    .C(_04843_),
    .D(_04846_),
    .X(_04847_));
 sky130_fd_sc_hd__a22o_1 _08824_ (.A1(\mix1.data_o[46] ),
    .A2(_04692_),
    .B1(_04694_),
    .B2(\mix1.data_o[38] ),
    .X(_04848_));
 sky130_fd_sc_hd__a22o_1 _08825_ (.A1(\addroundkey_data_o[46] ),
    .A2(_04692_),
    .B1(_04694_),
    .B2(\addroundkey_data_o[38] ),
    .X(_04849_));
 sky130_fd_sc_hd__mux2_1 _08826_ (.A0(_04848_),
    .A1(_04849_),
    .S(_04650_),
    .X(_04850_));
 sky130_fd_sc_hd__or2_1 _08827_ (.A(\addroundkey_data_o[102] ),
    .B(_04778_),
    .X(_04851_));
 sky130_fd_sc_hd__o211a_1 _08828_ (.A1(\mix1.data_o[102] ),
    .A2(_04650_),
    .B1(_04701_),
    .C1(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__mux2_1 _08829_ (.A0(\addroundkey_data_o[110] ),
    .A1(\mix1.data_o[110] ),
    .S(_04665_),
    .X(_04853_));
 sky130_fd_sc_hd__mux2_1 _08830_ (.A0(\addroundkey_data_o[14] ),
    .A1(\mix1.data_o[14] ),
    .S(_04803_),
    .X(_04854_));
 sky130_fd_sc_hd__a22o_1 _08831_ (.A1(_04706_),
    .A2(_04853_),
    .B1(_04854_),
    .B2(_04710_),
    .X(_04855_));
 sky130_fd_sc_hd__mux2_1 _08832_ (.A0(\addroundkey_data_o[70] ),
    .A1(\mix1.data_o[70] ),
    .S(_04665_),
    .X(_04856_));
 sky130_fd_sc_hd__mux2_1 _08833_ (.A0(\addroundkey_data_o[94] ),
    .A1(\mix1.data_o[94] ),
    .S(_04805_),
    .X(_04857_));
 sky130_fd_sc_hd__a22o_1 _08834_ (.A1(_04713_),
    .A2(_04856_),
    .B1(_04857_),
    .B2(_04716_),
    .X(_04858_));
 sky130_fd_sc_hd__or4_2 _08835_ (.A(_04850_),
    .B(_04852_),
    .C(_04855_),
    .D(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__a211o_1 _08836_ (.A1(_04653_),
    .A2(_04834_),
    .B1(_04847_),
    .C1(_04859_),
    .X(_04860_));
 sky130_fd_sc_hd__o31a_1 _08837_ (.A1(\ks1.key_reg[14] ),
    .A2(_04729_),
    .A3(_04731_),
    .B1(net163),
    .X(_04861_));
 sky130_fd_sc_hd__a21oi_1 _08838_ (.A1(\ks1.key_reg[14] ),
    .A2(_04725_),
    .B1(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__inv_2 _08839_ (.A(_04721_),
    .Y(_04863_));
 sky130_fd_sc_hd__or3_1 _08840_ (.A(\ks1.key_reg[6] ),
    .B(_04729_),
    .C(_04731_),
    .X(_04864_));
 sky130_fd_sc_hd__a22o_1 _08841_ (.A1(\ks1.key_reg[6] ),
    .A2(_04725_),
    .B1(_04864_),
    .B2(net224),
    .X(_04865_));
 sky130_fd_sc_hd__a2bb2o_1 _08842_ (.A1_N(_04862_),
    .A2_N(_04755_),
    .B1(_04863_),
    .B2(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__o31a_1 _08843_ (.A1(\ks1.key_reg[22] ),
    .A2(_04729_),
    .A3(_04731_),
    .B1(net172),
    .X(_04867_));
 sky130_fd_sc_hd__a21oi_1 _08844_ (.A1(\ks1.key_reg[22] ),
    .A2(_04725_),
    .B1(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__mux2_1 _08845_ (.A0(net181),
    .A1(\ks1.key_reg[30] ),
    .S(_04725_),
    .X(_04869_));
 sky130_fd_sc_hd__a2bb2o_1 _08846_ (.A1_N(_04741_),
    .A2_N(_04868_),
    .B1(_04869_),
    .B2(_04750_),
    .X(_04870_));
 sky130_fd_sc_hd__a211o_1 _08847_ (.A1(_04648_),
    .A2(_04860_),
    .B1(_04866_),
    .C1(_04870_),
    .X(_04871_));
 sky130_fd_sc_hd__inv_2 _08848_ (.A(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__xnor2_1 _08849_ (.A(_04833_),
    .B(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__and2_2 _08850_ (.A(_04624_),
    .B(_04648_),
    .X(_04874_));
 sky130_fd_sc_hd__o21a_1 _08851_ (.A1(_04794_),
    .A2(_04873_),
    .B1(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__nand2_1 _08852_ (.A(_04794_),
    .B(_04873_),
    .Y(_04876_));
 sky130_fd_sc_hd__a22o_4 _08853_ (.A1(_04649_),
    .A2(_04752_),
    .B1(_04875_),
    .B2(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__mux2_1 _08854_ (.A0(\addroundkey_data_o[120] ),
    .A1(\mix1.data_o[120] ),
    .S(_04658_),
    .X(_04878_));
 sky130_fd_sc_hd__buf_4 _08855_ (.A(_04661_),
    .X(_04879_));
 sky130_fd_sc_hd__buf_4 _08856_ (.A(_04805_),
    .X(_04880_));
 sky130_fd_sc_hd__mux2_1 _08857_ (.A0(\addroundkey_data_o[16] ),
    .A1(\mix1.data_o[16] ),
    .S(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__mux2_1 _08858_ (.A0(\addroundkey_data_o[72] ),
    .A1(\mix1.data_o[72] ),
    .S(_04702_),
    .X(_04882_));
 sky130_fd_sc_hd__a22o_1 _08859_ (.A1(_04879_),
    .A2(_04881_),
    .B1(_04882_),
    .B2(_04668_),
    .X(_04883_));
 sky130_fd_sc_hd__buf_4 _08860_ (.A(_04670_),
    .X(_04884_));
 sky130_fd_sc_hd__mux2_1 _08861_ (.A0(\addroundkey_data_o[48] ),
    .A1(\mix1.data_o[48] ),
    .S(_04666_),
    .X(_04885_));
 sky130_fd_sc_hd__mux2_1 _08862_ (.A0(\addroundkey_data_o[24] ),
    .A1(\mix1.data_o[24] ),
    .S(_04880_),
    .X(_04886_));
 sky130_fd_sc_hd__a22o_1 _08863_ (.A1(_04884_),
    .A2(_04885_),
    .B1(_04886_),
    .B2(_04675_),
    .X(_04887_));
 sky130_fd_sc_hd__buf_4 _08864_ (.A(_04677_),
    .X(_04888_));
 sky130_fd_sc_hd__mux2_1 _08865_ (.A0(\addroundkey_data_o[80] ),
    .A1(\mix1.data_o[80] ),
    .S(_04666_),
    .X(_04889_));
 sky130_fd_sc_hd__mux2_1 _08866_ (.A0(\addroundkey_data_o[112] ),
    .A1(\mix1.data_o[112] ),
    .S(_04880_),
    .X(_04890_));
 sky130_fd_sc_hd__clkbuf_8 _08867_ (.A(_04682_),
    .X(_04891_));
 sky130_fd_sc_hd__a22o_1 _08868_ (.A1(_04888_),
    .A2(_04889_),
    .B1(_04890_),
    .B2(_04891_),
    .X(_04892_));
 sky130_fd_sc_hd__mux2_1 _08869_ (.A0(\addroundkey_data_o[56] ),
    .A1(\mix1.data_o[56] ),
    .S(_04880_),
    .X(_04893_));
 sky130_fd_sc_hd__mux2_1 _08870_ (.A0(\addroundkey_data_o[0] ),
    .A1(\mix1.data_o[0] ),
    .S(_04702_),
    .X(_04894_));
 sky130_fd_sc_hd__a22o_1 _08871_ (.A1(_04684_),
    .A2(_04893_),
    .B1(_04894_),
    .B2(_04689_),
    .X(_04895_));
 sky130_fd_sc_hd__or4_1 _08872_ (.A(_04883_),
    .B(_04887_),
    .C(_04892_),
    .D(_04895_),
    .X(_04896_));
 sky130_fd_sc_hd__a22o_1 _08873_ (.A1(\mix1.data_o[40] ),
    .A2(_04693_),
    .B1(_04695_),
    .B2(\mix1.data_o[32] ),
    .X(_04897_));
 sky130_fd_sc_hd__a22o_1 _08874_ (.A1(\addroundkey_data_o[40] ),
    .A2(_04693_),
    .B1(_04695_),
    .B2(\addroundkey_data_o[32] ),
    .X(_04898_));
 sky130_fd_sc_hd__mux2_1 _08875_ (.A0(_04897_),
    .A1(_04898_),
    .S(_04698_),
    .X(_04899_));
 sky130_fd_sc_hd__clkbuf_4 _08876_ (.A(_04698_),
    .X(_04900_));
 sky130_fd_sc_hd__or2_1 _08877_ (.A(\addroundkey_data_o[96] ),
    .B(_04657_),
    .X(_04901_));
 sky130_fd_sc_hd__o211a_1 _08878_ (.A1(\mix1.data_o[96] ),
    .A2(_04900_),
    .B1(_04701_),
    .C1(_04901_),
    .X(_04902_));
 sky130_fd_sc_hd__mux2_1 _08879_ (.A0(\addroundkey_data_o[104] ),
    .A1(\mix1.data_o[104] ),
    .S(_04880_),
    .X(_04903_));
 sky130_fd_sc_hd__mux2_1 _08880_ (.A0(\addroundkey_data_o[8] ),
    .A1(\mix1.data_o[8] ),
    .S(_04702_),
    .X(_04904_));
 sky130_fd_sc_hd__a22o_1 _08881_ (.A1(_04706_),
    .A2(_04903_),
    .B1(_04904_),
    .B2(_04710_),
    .X(_04905_));
 sky130_fd_sc_hd__mux2_1 _08882_ (.A0(\addroundkey_data_o[64] ),
    .A1(\mix1.data_o[64] ),
    .S(_04880_),
    .X(_04906_));
 sky130_fd_sc_hd__mux2_1 _08883_ (.A0(\addroundkey_data_o[88] ),
    .A1(\mix1.data_o[88] ),
    .S(_04702_),
    .X(_04907_));
 sky130_fd_sc_hd__a22o_1 _08884_ (.A1(_04713_),
    .A2(_04906_),
    .B1(_04907_),
    .B2(_04716_),
    .X(_04908_));
 sky130_fd_sc_hd__or4_1 _08885_ (.A(_04899_),
    .B(_04902_),
    .C(_04905_),
    .D(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__a211o_2 _08886_ (.A1(_04653_),
    .A2(_04878_),
    .B1(_04896_),
    .C1(_04909_),
    .X(_04910_));
 sky130_fd_sc_hd__buf_4 _08887_ (.A(_04738_),
    .X(_04911_));
 sky130_fd_sc_hd__or3_1 _08888_ (.A(\ks1.key_reg[8] ),
    .B(_04745_),
    .C(_04746_),
    .X(_04912_));
 sky130_fd_sc_hd__a22o_1 _08889_ (.A1(\ks1.key_reg[8] ),
    .A2(_04726_),
    .B1(_04912_),
    .B2(net246),
    .X(_04913_));
 sky130_fd_sc_hd__or3_1 _08890_ (.A(\ks1.key_reg[16] ),
    .B(_04745_),
    .C(_04746_),
    .X(_04914_));
 sky130_fd_sc_hd__a22o_1 _08891_ (.A1(\ks1.key_reg[16] ),
    .A2(_04726_),
    .B1(_04914_),
    .B2(net165),
    .X(_04915_));
 sky130_fd_sc_hd__inv_4 _08892_ (.A(_04741_),
    .Y(_04916_));
 sky130_fd_sc_hd__o31a_1 _08893_ (.A1(\ks1.key_reg[24] ),
    .A2(_04729_),
    .A3(_04731_),
    .B1(net174),
    .X(_04917_));
 sky130_fd_sc_hd__a21oi_1 _08894_ (.A1(\ks1.key_reg[24] ),
    .A2(_04735_),
    .B1(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__or3_1 _08895_ (.A(\ks1.key_reg[0] ),
    .B(_04729_),
    .C(_04731_),
    .X(_04919_));
 sky130_fd_sc_hd__a22o_1 _08896_ (.A1(\ks1.key_reg[0] ),
    .A2(_04725_),
    .B1(_04919_),
    .B2(net130),
    .X(_04920_));
 sky130_fd_sc_hd__a2bb2o_1 _08897_ (.A1_N(_04645_),
    .A2_N(_04918_),
    .B1(_04863_),
    .B2(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__a221o_2 _08898_ (.A1(_04911_),
    .A2(_04913_),
    .B1(_04915_),
    .B2(_04916_),
    .C1(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__a21oi_2 _08899_ (.A1(_04648_),
    .A2(_04910_),
    .B1(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__mux2_1 _08900_ (.A0(\addroundkey_data_o[125] ),
    .A1(\mix1.data_o[125] ),
    .S(_04658_),
    .X(_04924_));
 sky130_fd_sc_hd__mux2_1 _08901_ (.A0(\addroundkey_data_o[21] ),
    .A1(\mix1.data_o[21] ),
    .S(_04880_),
    .X(_04925_));
 sky130_fd_sc_hd__mux2_1 _08902_ (.A0(\addroundkey_data_o[77] ),
    .A1(\mix1.data_o[77] ),
    .S(_04657_),
    .X(_04926_));
 sky130_fd_sc_hd__buf_4 _08903_ (.A(_04668_),
    .X(_04927_));
 sky130_fd_sc_hd__a22o_1 _08904_ (.A1(_04879_),
    .A2(_04925_),
    .B1(_04926_),
    .B2(_04927_),
    .X(_04928_));
 sky130_fd_sc_hd__mux2_1 _08905_ (.A0(\addroundkey_data_o[53] ),
    .A1(\mix1.data_o[53] ),
    .S(_04880_),
    .X(_04929_));
 sky130_fd_sc_hd__mux2_1 _08906_ (.A0(\addroundkey_data_o[29] ),
    .A1(\mix1.data_o[29] ),
    .S(_04702_),
    .X(_04930_));
 sky130_fd_sc_hd__a22o_1 _08907_ (.A1(_04884_),
    .A2(_04929_),
    .B1(_04930_),
    .B2(_04675_),
    .X(_04931_));
 sky130_fd_sc_hd__mux2_1 _08908_ (.A0(\addroundkey_data_o[85] ),
    .A1(\mix1.data_o[85] ),
    .S(_04880_),
    .X(_04932_));
 sky130_fd_sc_hd__mux2_1 _08909_ (.A0(\addroundkey_data_o[117] ),
    .A1(\mix1.data_o[117] ),
    .S(_04702_),
    .X(_04933_));
 sky130_fd_sc_hd__a22o_1 _08910_ (.A1(_04888_),
    .A2(_04932_),
    .B1(_04933_),
    .B2(_04891_),
    .X(_04934_));
 sky130_fd_sc_hd__clkbuf_4 _08911_ (.A(_04684_),
    .X(_04935_));
 sky130_fd_sc_hd__mux2_1 _08912_ (.A0(\addroundkey_data_o[61] ),
    .A1(\mix1.data_o[61] ),
    .S(_04880_),
    .X(_04936_));
 sky130_fd_sc_hd__mux2_1 _08913_ (.A0(\addroundkey_data_o[5] ),
    .A1(\mix1.data_o[5] ),
    .S(_04657_),
    .X(_04937_));
 sky130_fd_sc_hd__a22o_1 _08914_ (.A1(_04935_),
    .A2(_04936_),
    .B1(_04937_),
    .B2(_04689_),
    .X(_04938_));
 sky130_fd_sc_hd__or4_1 _08915_ (.A(_04928_),
    .B(_04931_),
    .C(_04934_),
    .D(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__a22o_1 _08916_ (.A1(\mix1.data_o[45] ),
    .A2(_04693_),
    .B1(_04695_),
    .B2(\mix1.data_o[37] ),
    .X(_04940_));
 sky130_fd_sc_hd__a22o_1 _08917_ (.A1(\addroundkey_data_o[45] ),
    .A2(_04693_),
    .B1(_04695_),
    .B2(\addroundkey_data_o[37] ),
    .X(_04941_));
 sky130_fd_sc_hd__mux2_1 _08918_ (.A0(_04940_),
    .A1(_04941_),
    .S(_04900_),
    .X(_04942_));
 sky130_fd_sc_hd__clkbuf_4 _08919_ (.A(_04701_),
    .X(_04943_));
 sky130_fd_sc_hd__or2_1 _08920_ (.A(\addroundkey_data_o[101] ),
    .B(_04657_),
    .X(_04944_));
 sky130_fd_sc_hd__o211a_1 _08921_ (.A1(\mix1.data_o[101] ),
    .A2(_04900_),
    .B1(_04943_),
    .C1(_04944_),
    .X(_04945_));
 sky130_fd_sc_hd__clkbuf_4 _08922_ (.A(_04706_),
    .X(_04946_));
 sky130_fd_sc_hd__mux2_1 _08923_ (.A0(\addroundkey_data_o[109] ),
    .A1(\mix1.data_o[109] ),
    .S(_04702_),
    .X(_04947_));
 sky130_fd_sc_hd__mux2_1 _08924_ (.A0(\addroundkey_data_o[13] ),
    .A1(\mix1.data_o[13] ),
    .S(_04657_),
    .X(_04948_));
 sky130_fd_sc_hd__clkbuf_4 _08925_ (.A(_04710_),
    .X(_04949_));
 sky130_fd_sc_hd__a22o_1 _08926_ (.A1(_04946_),
    .A2(_04947_),
    .B1(_04948_),
    .B2(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__mux2_1 _08927_ (.A0(\addroundkey_data_o[69] ),
    .A1(\mix1.data_o[69] ),
    .S(_04702_),
    .X(_04951_));
 sky130_fd_sc_hd__mux2_1 _08928_ (.A0(\addroundkey_data_o[93] ),
    .A1(\mix1.data_o[93] ),
    .S(_04657_),
    .X(_04952_));
 sky130_fd_sc_hd__a22o_1 _08929_ (.A1(_04713_),
    .A2(_04951_),
    .B1(_04952_),
    .B2(_04716_),
    .X(_04953_));
 sky130_fd_sc_hd__or4_1 _08930_ (.A(_04942_),
    .B(_04945_),
    .C(_04950_),
    .D(_04953_),
    .X(_04954_));
 sky130_fd_sc_hd__a211o_2 _08931_ (.A1(_04653_),
    .A2(_04924_),
    .B1(_04939_),
    .C1(_04954_),
    .X(_04955_));
 sky130_fd_sc_hd__or3_1 _08932_ (.A(\ks1.key_reg[21] ),
    .B(_04730_),
    .C(_04732_),
    .X(_04956_));
 sky130_fd_sc_hd__a22o_1 _08933_ (.A1(\ks1.key_reg[21] ),
    .A2(_04726_),
    .B1(_04956_),
    .B2(net171),
    .X(_04957_));
 sky130_fd_sc_hd__or3_1 _08934_ (.A(\ks1.key_reg[13] ),
    .B(_04730_),
    .C(_04732_),
    .X(_04958_));
 sky130_fd_sc_hd__a22o_1 _08935_ (.A1(\ks1.key_reg[13] ),
    .A2(_04726_),
    .B1(_04958_),
    .B2(net162),
    .X(_04959_));
 sky130_fd_sc_hd__o31a_1 _08936_ (.A1(\ks1.key_reg[5] ),
    .A2(_04745_),
    .A3(_04746_),
    .B1(net213),
    .X(_04960_));
 sky130_fd_sc_hd__a21oi_2 _08937_ (.A1(\ks1.key_reg[5] ),
    .A2(_04735_),
    .B1(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__or3_1 _08938_ (.A(\ks1.key_reg[29] ),
    .B(_04729_),
    .C(_04731_),
    .X(_04962_));
 sky130_fd_sc_hd__a22o_1 _08939_ (.A1(\ks1.key_reg[29] ),
    .A2(_04725_),
    .B1(_04962_),
    .B2(net179),
    .X(_04963_));
 sky130_fd_sc_hd__a2bb2o_1 _08940_ (.A1_N(_04721_),
    .A2_N(_04961_),
    .B1(_04963_),
    .B2(_04750_),
    .X(_04964_));
 sky130_fd_sc_hd__a221o_2 _08941_ (.A1(_04916_),
    .A2(_04957_),
    .B1(_04959_),
    .B2(_04911_),
    .C1(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__a21oi_2 _08942_ (.A1(_04648_),
    .A2(_04955_),
    .B1(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__xnor2_2 _08943_ (.A(_04923_),
    .B(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__nor2_1 _08944_ (.A(_04833_),
    .B(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__a21o_1 _08945_ (.A1(_04833_),
    .A2(_04967_),
    .B1(_04649_),
    .X(_04969_));
 sky130_fd_sc_hd__o22a_2 _08946_ (.A1(_04874_),
    .A2(_04872_),
    .B1(_04968_),
    .B2(_04969_),
    .X(_04970_));
 sky130_fd_sc_hd__xor2_4 _08947_ (.A(_04877_),
    .B(_04970_),
    .X(_04971_));
 sky130_fd_sc_hd__mux2_1 _08948_ (.A0(\addroundkey_data_o[127] ),
    .A1(\mix1.data_o[127] ),
    .S(_04658_),
    .X(_04972_));
 sky130_fd_sc_hd__mux2_1 _08949_ (.A0(\addroundkey_data_o[23] ),
    .A1(\mix1.data_o[23] ),
    .S(_04656_),
    .X(_04973_));
 sky130_fd_sc_hd__mux2_1 _08950_ (.A0(\addroundkey_data_o[79] ),
    .A1(\mix1.data_o[79] ),
    .S(_04778_),
    .X(_04974_));
 sky130_fd_sc_hd__a22o_1 _08951_ (.A1(_04661_),
    .A2(_04973_),
    .B1(_04974_),
    .B2(_04668_),
    .X(_04975_));
 sky130_fd_sc_hd__mux2_1 _08952_ (.A0(\addroundkey_data_o[55] ),
    .A1(\mix1.data_o[55] ),
    .S(_04656_),
    .X(_04976_));
 sky130_fd_sc_hd__mux2_1 _08953_ (.A0(\addroundkey_data_o[31] ),
    .A1(\mix1.data_o[31] ),
    .S(_04778_),
    .X(_04977_));
 sky130_fd_sc_hd__a22o_1 _08954_ (.A1(_04670_),
    .A2(_04976_),
    .B1(_04977_),
    .B2(_04675_),
    .X(_04978_));
 sky130_fd_sc_hd__mux2_1 _08955_ (.A0(\addroundkey_data_o[87] ),
    .A1(\mix1.data_o[87] ),
    .S(_04656_),
    .X(_04979_));
 sky130_fd_sc_hd__mux2_1 _08956_ (.A0(\addroundkey_data_o[119] ),
    .A1(\mix1.data_o[119] ),
    .S(_04778_),
    .X(_04980_));
 sky130_fd_sc_hd__a22o_1 _08957_ (.A1(_04677_),
    .A2(_04979_),
    .B1(_04980_),
    .B2(_04682_),
    .X(_04981_));
 sky130_fd_sc_hd__mux2_1 _08958_ (.A0(\addroundkey_data_o[63] ),
    .A1(\mix1.data_o[63] ),
    .S(_04778_),
    .X(_04982_));
 sky130_fd_sc_hd__mux2_1 _08959_ (.A0(\addroundkey_data_o[7] ),
    .A1(\mix1.data_o[7] ),
    .S(_04663_),
    .X(_04983_));
 sky130_fd_sc_hd__a22o_1 _08960_ (.A1(_04684_),
    .A2(_04982_),
    .B1(_04983_),
    .B2(_04689_),
    .X(_04984_));
 sky130_fd_sc_hd__or4_1 _08961_ (.A(_04975_),
    .B(_04978_),
    .C(_04981_),
    .D(_04984_),
    .X(_04985_));
 sky130_fd_sc_hd__a22o_1 _08962_ (.A1(\mix1.data_o[47] ),
    .A2(_04693_),
    .B1(_04695_),
    .B2(\mix1.data_o[39] ),
    .X(_04986_));
 sky130_fd_sc_hd__a22o_1 _08963_ (.A1(\addroundkey_data_o[47] ),
    .A2(_04693_),
    .B1(_04695_),
    .B2(\addroundkey_data_o[39] ),
    .X(_04987_));
 sky130_fd_sc_hd__mux2_1 _08964_ (.A0(_04986_),
    .A1(_04987_),
    .S(_04698_),
    .X(_04988_));
 sky130_fd_sc_hd__or2_1 _08965_ (.A(\addroundkey_data_o[103] ),
    .B(_04666_),
    .X(_04989_));
 sky130_fd_sc_hd__o211a_1 _08966_ (.A1(\mix1.data_o[103] ),
    .A2(_04698_),
    .B1(_04701_),
    .C1(_04989_),
    .X(_04990_));
 sky130_fd_sc_hd__mux2_1 _08967_ (.A0(\addroundkey_data_o[111] ),
    .A1(\mix1.data_o[111] ),
    .S(_04778_),
    .X(_04991_));
 sky130_fd_sc_hd__mux2_1 _08968_ (.A0(\addroundkey_data_o[15] ),
    .A1(\mix1.data_o[15] ),
    .S(_04663_),
    .X(_04992_));
 sky130_fd_sc_hd__a22o_1 _08969_ (.A1(_04706_),
    .A2(_04991_),
    .B1(_04992_),
    .B2(_04710_),
    .X(_04993_));
 sky130_fd_sc_hd__mux2_1 _08970_ (.A0(\addroundkey_data_o[71] ),
    .A1(\mix1.data_o[71] ),
    .S(_04778_),
    .X(_04994_));
 sky130_fd_sc_hd__mux2_1 _08971_ (.A0(\addroundkey_data_o[95] ),
    .A1(\mix1.data_o[95] ),
    .S(_04663_),
    .X(_04995_));
 sky130_fd_sc_hd__a22o_1 _08972_ (.A1(_04713_),
    .A2(_04994_),
    .B1(_04995_),
    .B2(_04716_),
    .X(_04996_));
 sky130_fd_sc_hd__or4_2 _08973_ (.A(_04988_),
    .B(_04990_),
    .C(_04993_),
    .D(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__a211o_1 _08974_ (.A1(_04653_),
    .A2(_04972_),
    .B1(_04985_),
    .C1(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__o31a_1 _08975_ (.A1(\ks1.key_reg[23] ),
    .A2(_04745_),
    .A3(_04746_),
    .B1(net173),
    .X(_04999_));
 sky130_fd_sc_hd__a21oi_1 _08976_ (.A1(\ks1.key_reg[23] ),
    .A2(_04735_),
    .B1(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__or3_1 _08977_ (.A(\ks1.key_reg[31] ),
    .B(_04729_),
    .C(_04731_),
    .X(_05001_));
 sky130_fd_sc_hd__a22o_1 _08978_ (.A1(\ks1.key_reg[31] ),
    .A2(_04725_),
    .B1(_05001_),
    .B2(net182),
    .X(_05002_));
 sky130_fd_sc_hd__a2bb2o_1 _08979_ (.A1_N(_05000_),
    .A2_N(_04741_),
    .B1(_04750_),
    .B2(_05002_),
    .X(_05003_));
 sky130_fd_sc_hd__o31a_1 _08980_ (.A1(\ks1.key_reg[15] ),
    .A2(_04745_),
    .A3(_04746_),
    .B1(net164),
    .X(_05004_));
 sky130_fd_sc_hd__a21oi_1 _08981_ (.A1(\ks1.key_reg[15] ),
    .A2(_04726_),
    .B1(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__or3_1 _08982_ (.A(\ks1.key_reg[7] ),
    .B(_04729_),
    .C(_04731_),
    .X(_05006_));
 sky130_fd_sc_hd__a22o_1 _08983_ (.A1(\ks1.key_reg[7] ),
    .A2(_04725_),
    .B1(_05006_),
    .B2(net235),
    .X(_05007_));
 sky130_fd_sc_hd__clkbuf_8 _08984_ (.A(_04863_),
    .X(_00007_));
 sky130_fd_sc_hd__a2bb2o_1 _08985_ (.A1_N(_04755_),
    .A2_N(_05005_),
    .B1(_05007_),
    .B2(_00007_),
    .X(_05008_));
 sky130_fd_sc_hd__a211o_2 _08986_ (.A1(_04648_),
    .A2(_04998_),
    .B1(_05003_),
    .C1(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__xor2_1 _08987_ (.A(_04794_),
    .B(_04752_),
    .X(_05010_));
 sky130_fd_sc_hd__a21o_1 _08988_ (.A1(_04872_),
    .A2(_05010_),
    .B1(_04649_),
    .X(_05011_));
 sky130_fd_sc_hd__nor2_1 _08989_ (.A(_04872_),
    .B(_05010_),
    .Y(_05012_));
 sky130_fd_sc_hd__o2bb2a_4 _08990_ (.A1_N(_04649_),
    .A2_N(_05009_),
    .B1(_05011_),
    .B2(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__xnor2_1 _08991_ (.A(_04873_),
    .B(_04923_),
    .Y(_05014_));
 sky130_fd_sc_hd__mux2_4 _08992_ (.A0(_04794_),
    .A1(_05014_),
    .S(_04874_),
    .X(_05015_));
 sky130_fd_sc_hd__xor2_4 _08993_ (.A(_05013_),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__xnor2_4 _08994_ (.A(_04971_),
    .B(_05016_),
    .Y(\sbox1.ah[1] ));
 sky130_fd_sc_hd__mux2_1 _08995_ (.A0(\addroundkey_data_o[122] ),
    .A1(\mix1.data_o[122] ),
    .S(_04657_),
    .X(_05017_));
 sky130_fd_sc_hd__mux2_1 _08996_ (.A0(\addroundkey_data_o[18] ),
    .A1(\mix1.data_o[18] ),
    .S(_04665_),
    .X(_05018_));
 sky130_fd_sc_hd__mux2_1 _08997_ (.A0(\addroundkey_data_o[74] ),
    .A1(\mix1.data_o[74] ),
    .S(_04803_),
    .X(_05019_));
 sky130_fd_sc_hd__a22o_1 _08998_ (.A1(_04661_),
    .A2(_05018_),
    .B1(_05019_),
    .B2(_04668_),
    .X(_05020_));
 sky130_fd_sc_hd__mux2_1 _08999_ (.A0(\addroundkey_data_o[50] ),
    .A1(\mix1.data_o[50] ),
    .S(_04662_),
    .X(_05021_));
 sky130_fd_sc_hd__mux2_1 _09000_ (.A0(\addroundkey_data_o[26] ),
    .A1(\mix1.data_o[26] ),
    .S(_04803_),
    .X(_05022_));
 sky130_fd_sc_hd__a22o_1 _09001_ (.A1(_04670_),
    .A2(_05021_),
    .B1(_05022_),
    .B2(_04675_),
    .X(_05023_));
 sky130_fd_sc_hd__mux2_1 _09002_ (.A0(\addroundkey_data_o[82] ),
    .A1(\mix1.data_o[82] ),
    .S(_04662_),
    .X(_05024_));
 sky130_fd_sc_hd__mux2_1 _09003_ (.A0(\addroundkey_data_o[114] ),
    .A1(\mix1.data_o[114] ),
    .S(_04803_),
    .X(_05025_));
 sky130_fd_sc_hd__a22o_1 _09004_ (.A1(_04677_),
    .A2(_05024_),
    .B1(_05025_),
    .B2(_04682_),
    .X(_05026_));
 sky130_fd_sc_hd__mux2_1 _09005_ (.A0(\addroundkey_data_o[58] ),
    .A1(\mix1.data_o[58] ),
    .S(_04665_),
    .X(_05027_));
 sky130_fd_sc_hd__mux2_1 _09006_ (.A0(\addroundkey_data_o[2] ),
    .A1(\mix1.data_o[2] ),
    .S(_04805_),
    .X(_05028_));
 sky130_fd_sc_hd__a22o_1 _09007_ (.A1(_04684_),
    .A2(_05027_),
    .B1(_05028_),
    .B2(_04689_),
    .X(_05029_));
 sky130_fd_sc_hd__or4_1 _09008_ (.A(_05020_),
    .B(_05023_),
    .C(_05026_),
    .D(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__a22o_1 _09009_ (.A1(\mix1.data_o[42] ),
    .A2(_04692_),
    .B1(_04694_),
    .B2(\mix1.data_o[34] ),
    .X(_05031_));
 sky130_fd_sc_hd__a22o_1 _09010_ (.A1(\addroundkey_data_o[42] ),
    .A2(_04692_),
    .B1(_04694_),
    .B2(\addroundkey_data_o[34] ),
    .X(_05032_));
 sky130_fd_sc_hd__mux2_1 _09011_ (.A0(_05031_),
    .A1(_05032_),
    .S(_04650_),
    .X(_05033_));
 sky130_fd_sc_hd__or2_1 _09012_ (.A(\addroundkey_data_o[98] ),
    .B(_04778_),
    .X(_05034_));
 sky130_fd_sc_hd__o211a_1 _09013_ (.A1(\mix1.data_o[98] ),
    .A2(_04698_),
    .B1(_04701_),
    .C1(_05034_),
    .X(_05035_));
 sky130_fd_sc_hd__mux2_1 _09014_ (.A0(\addroundkey_data_o[106] ),
    .A1(\mix1.data_o[106] ),
    .S(_04665_),
    .X(_05036_));
 sky130_fd_sc_hd__mux2_1 _09015_ (.A0(\addroundkey_data_o[10] ),
    .A1(\mix1.data_o[10] ),
    .S(_04805_),
    .X(_05037_));
 sky130_fd_sc_hd__a22o_1 _09016_ (.A1(_04706_),
    .A2(_05036_),
    .B1(_05037_),
    .B2(_04710_),
    .X(_05038_));
 sky130_fd_sc_hd__mux2_1 _09017_ (.A0(\addroundkey_data_o[66] ),
    .A1(\mix1.data_o[66] ),
    .S(_04665_),
    .X(_05039_));
 sky130_fd_sc_hd__mux2_1 _09018_ (.A0(\addroundkey_data_o[90] ),
    .A1(\mix1.data_o[90] ),
    .S(_04805_),
    .X(_05040_));
 sky130_fd_sc_hd__a22o_1 _09019_ (.A1(_04713_),
    .A2(_05039_),
    .B1(_05040_),
    .B2(_04716_),
    .X(_05041_));
 sky130_fd_sc_hd__or4_1 _09020_ (.A(_05033_),
    .B(_05035_),
    .C(_05038_),
    .D(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__a211o_2 _09021_ (.A1(_04653_),
    .A2(_05017_),
    .B1(_05030_),
    .C1(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__nand2_1 _09022_ (.A(_04648_),
    .B(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__o31a_1 _09023_ (.A1(\ks1.key_reg[26] ),
    .A2(_04745_),
    .A3(_04746_),
    .B1(net176),
    .X(_05045_));
 sky130_fd_sc_hd__a21oi_2 _09024_ (.A1(\ks1.key_reg[26] ),
    .A2(_04735_),
    .B1(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__o31a_1 _09025_ (.A1(\ks1.key_reg[10] ),
    .A2(_04745_),
    .A3(_04746_),
    .B1(net141),
    .X(_05047_));
 sky130_fd_sc_hd__a21oi_1 _09026_ (.A1(\ks1.key_reg[10] ),
    .A2(_04735_),
    .B1(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__o22a_1 _09027_ (.A1(_04645_),
    .A2(_05046_),
    .B1(_05048_),
    .B2(_04755_),
    .X(_05049_));
 sky130_fd_sc_hd__mux2_1 _09028_ (.A0(net180),
    .A1(\ks1.key_reg[2] ),
    .S(_04725_),
    .X(_05050_));
 sky130_fd_sc_hd__o31a_1 _09029_ (.A1(\ks1.key_reg[18] ),
    .A2(_04745_),
    .A3(_04746_),
    .B1(net167),
    .X(_05051_));
 sky130_fd_sc_hd__a21oi_1 _09030_ (.A1(\ks1.key_reg[18] ),
    .A2(_04735_),
    .B1(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__o2bb2a_1 _09031_ (.A1_N(_04863_),
    .A2_N(_05050_),
    .B1(_05052_),
    .B2(_04741_),
    .X(_05053_));
 sky130_fd_sc_hd__and3_2 _09032_ (.A(_05044_),
    .B(_05049_),
    .C(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__xnor2_2 _09033_ (.A(_05009_),
    .B(_05054_),
    .Y(_05055_));
 sky130_fd_sc_hd__xnor2_1 _09034_ (.A(_04752_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__mux2_4 _09035_ (.A0(_04966_),
    .A1(_05056_),
    .S(_04874_),
    .X(_05057_));
 sky130_fd_sc_hd__xnor2_4 _09036_ (.A(_05013_),
    .B(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__inv_2 _09037_ (.A(_05058_),
    .Y(\sbox1.ah[3] ));
 sky130_fd_sc_hd__xor2_4 _09038_ (.A(_04971_),
    .B(_05057_),
    .X(\sbox1.ah[0] ));
 sky130_fd_sc_hd__xnor2_1 _09039_ (.A(_04967_),
    .B(_05054_),
    .Y(_05059_));
 sky130_fd_sc_hd__buf_4 _09040_ (.A(_04874_),
    .X(_05060_));
 sky130_fd_sc_hd__mux2_1 _09041_ (.A0(_04833_),
    .A1(_05059_),
    .S(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__nand2_1 _09042_ (.A(_05010_),
    .B(_05009_),
    .Y(_05062_));
 sky130_fd_sc_hd__or2_1 _09043_ (.A(_05010_),
    .B(_05009_),
    .X(_05063_));
 sky130_fd_sc_hd__nor2_1 _09044_ (.A(_05060_),
    .B(_05054_),
    .Y(_05064_));
 sky130_fd_sc_hd__a31o_4 _09045_ (.A1(_05060_),
    .A2(_05062_),
    .A3(_05063_),
    .B1(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__xnor2_1 _09046_ (.A(_05058_),
    .B(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__xnor2_2 _09047_ (.A(_05061_),
    .B(_05066_),
    .Y(\sbox1.ah[2] ));
 sky130_fd_sc_hd__xnor2_4 _09048_ (.A(_04877_),
    .B(_05065_),
    .Y(_05067_));
 sky130_fd_sc_hd__xor2_1 _09049_ (.A(_05058_),
    .B(_05067_),
    .X(\sbox1.next_alph[3] ));
 sky130_fd_sc_hd__or2_1 _09050_ (.A(_05016_),
    .B(\sbox1.ah[2] ),
    .X(_05068_));
 sky130_fd_sc_hd__nand2_1 _09051_ (.A(_05016_),
    .B(\sbox1.ah[2] ),
    .Y(_05069_));
 sky130_fd_sc_hd__and2_1 _09052_ (.A(_05068_),
    .B(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__clkbuf_1 _09053_ (.A(_05070_),
    .X(\sbox1.next_alph[2] ));
 sky130_fd_sc_hd__xnor2_4 _09054_ (.A(_05015_),
    .B(_05065_),
    .Y(_05071_));
 sky130_fd_sc_hd__xor2_1 _09055_ (.A(\sbox1.ah[1] ),
    .B(_05071_),
    .X(\sbox1.next_alph[1] ));
 sky130_fd_sc_hd__nor2_1 _09056_ (.A(_04966_),
    .B(_05055_),
    .Y(_05072_));
 sky130_fd_sc_hd__a21o_1 _09057_ (.A1(_04966_),
    .A2(_05055_),
    .B1(_04649_),
    .X(_05073_));
 sky130_fd_sc_hd__o22a_1 _09058_ (.A1(_05060_),
    .A2(_04923_),
    .B1(_05072_),
    .B2(_05073_),
    .X(_05074_));
 sky130_fd_sc_hd__inv_2 _09059_ (.A(_05074_),
    .Y(\sbox1.next_alph[0] ));
 sky130_fd_sc_hd__nand2_1 _09060_ (.A(\sbox1.ah[2] ),
    .B(_05071_),
    .Y(_05075_));
 sky130_fd_sc_hd__nor2_1 _09061_ (.A(_04971_),
    .B(_05016_),
    .Y(_05076_));
 sky130_fd_sc_hd__xnor2_1 _09062_ (.A(\sbox1.ah[0] ),
    .B(\sbox1.next_alph[0] ),
    .Y(_05077_));
 sky130_fd_sc_hd__mux2_1 _09063_ (.A0(_05058_),
    .A1(\sbox1.ah[0] ),
    .S(_05067_),
    .X(_05078_));
 sky130_fd_sc_hd__o21ba_1 _09064_ (.A1(_05058_),
    .A2(_05077_),
    .B1_N(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__a41o_1 _09065_ (.A1(\sbox1.ah[3] ),
    .A2(\sbox1.ah[0] ),
    .A3(_05067_),
    .A4(_05074_),
    .B1(_05079_),
    .X(_05080_));
 sky130_fd_sc_hd__xnor2_1 _09066_ (.A(_05076_),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__xnor2_1 _09067_ (.A(_05075_),
    .B(_05081_),
    .Y(\sbox1.intermediate_to_invert_var[3] ));
 sky130_fd_sc_hd__a22oi_1 _09068_ (.A1(_05016_),
    .A2(\sbox1.ah[0] ),
    .B1(_05071_),
    .B2(\sbox1.ah[1] ),
    .Y(_05082_));
 sky130_fd_sc_hd__and4b_1 _09069_ (.A_N(_05057_),
    .B(_05071_),
    .C(_04971_),
    .D(_05016_),
    .X(_05083_));
 sky130_fd_sc_hd__nor2_1 _09070_ (.A(_05082_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__xor2_1 _09071_ (.A(_05016_),
    .B(_05067_),
    .X(_05085_));
 sky130_fd_sc_hd__nor2_1 _09072_ (.A(_05058_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__xnor2_1 _09073_ (.A(_05084_),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__xor2_1 _09074_ (.A(_05067_),
    .B(_05077_),
    .X(_05088_));
 sky130_fd_sc_hd__nand2_1 _09075_ (.A(\sbox1.ah[2] ),
    .B(_05088_),
    .Y(_05089_));
 sky130_fd_sc_hd__xnor2_1 _09076_ (.A(_05087_),
    .B(_05089_),
    .Y(_05090_));
 sky130_fd_sc_hd__xnor2_1 _09077_ (.A(_04877_),
    .B(_05090_),
    .Y(\sbox1.intermediate_to_invert_var[2] ));
 sky130_fd_sc_hd__inv_2 _09078_ (.A(\sbox1.ah[0] ),
    .Y(_05091_));
 sky130_fd_sc_hd__nor2_1 _09079_ (.A(_05091_),
    .B(_05071_),
    .Y(_05092_));
 sky130_fd_sc_hd__nand2_1 _09080_ (.A(\sbox1.ah[1] ),
    .B(_05088_),
    .Y(_05093_));
 sky130_fd_sc_hd__and2_1 _09081_ (.A(\sbox1.ah[3] ),
    .B(_05071_),
    .X(_05094_));
 sky130_fd_sc_hd__a21o_1 _09082_ (.A1(_05016_),
    .A2(_05058_),
    .B1(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__or2b_1 _09083_ (.A(_05085_),
    .B_N(\sbox1.ah[2] ),
    .X(_05096_));
 sky130_fd_sc_hd__xor2_1 _09084_ (.A(_05095_),
    .B(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__xnor2_1 _09085_ (.A(_05093_),
    .B(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__xnor2_1 _09086_ (.A(_05092_),
    .B(_05098_),
    .Y(\sbox1.intermediate_to_invert_var[1] ));
 sky130_fd_sc_hd__nand2_1 _09087_ (.A(\sbox1.ah[1] ),
    .B(_05067_),
    .Y(_05099_));
 sky130_fd_sc_hd__xnor2_1 _09088_ (.A(_05094_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__nor2_1 _09089_ (.A(\sbox1.ah[0] ),
    .B(_05074_),
    .Y(_05101_));
 sky130_fd_sc_hd__xnor2_1 _09090_ (.A(_05068_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__xnor2_1 _09091_ (.A(_05100_),
    .B(_05102_),
    .Y(\sbox1.intermediate_to_invert_var[0] ));
 sky130_fd_sc_hd__clkbuf_4 _09092_ (.A(_04367_),
    .X(_05103_));
 sky130_fd_sc_hd__clkbuf_4 _09093_ (.A(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__buf_2 _09094_ (.A(\sbox1.inversion_to_invert_var[2] ),
    .X(_05105_));
 sky130_fd_sc_hd__or3_1 _09095_ (.A(_05105_),
    .B(\sbox1.inversion_to_invert_var[3] ),
    .C(\sbox1.inversion_to_invert_var[0] ),
    .X(_05106_));
 sky130_fd_sc_hd__nand2_1 _09096_ (.A(_05105_),
    .B(\sbox1.inversion_to_invert_var[3] ),
    .Y(_05107_));
 sky130_fd_sc_hd__or2b_1 _09097_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B_N(\sbox1.inversion_to_invert_var[0] ),
    .X(_05108_));
 sky130_fd_sc_hd__nand3_2 _09098_ (.A(_05106_),
    .B(_05107_),
    .C(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__or2_2 _09099_ (.A(_05107_),
    .B(_05108_),
    .X(_05110_));
 sky130_fd_sc_hd__nand2_2 _09100_ (.A(_05109_),
    .B(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__nand2_1 _09101_ (.A(\sbox1.alph[0] ),
    .B(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__inv_2 _09102_ (.A(\sbox1.inversion_to_invert_var[3] ),
    .Y(_05113_));
 sky130_fd_sc_hd__xnor2_1 _09103_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B(\sbox1.inversion_to_invert_var[2] ),
    .Y(_05114_));
 sky130_fd_sc_hd__and2_1 _09104_ (.A(\sbox1.inversion_to_invert_var[3] ),
    .B(\sbox1.inversion_to_invert_var[0] ),
    .X(_05115_));
 sky130_fd_sc_hd__nand2_1 _09105_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B(_05105_),
    .Y(_05116_));
 sky130_fd_sc_hd__and3b_1 _09106_ (.A_N(\sbox1.inversion_to_invert_var[0] ),
    .B(_05105_),
    .C(\sbox1.inversion_to_invert_var[1] ),
    .X(_05117_));
 sky130_fd_sc_hd__a221oi_1 _09107_ (.A1(_05113_),
    .A2(_05114_),
    .B1(_05115_),
    .B2(_05116_),
    .C1(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__buf_2 _09108_ (.A(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__a21oi_1 _09109_ (.A1(_05109_),
    .A2(_05110_),
    .B1(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__and3_1 _09110_ (.A(_05109_),
    .B(_05110_),
    .C(_05118_),
    .X(_05121_));
 sky130_fd_sc_hd__o21a_1 _09111_ (.A1(_05120_),
    .A2(_05121_),
    .B1(\sbox1.alph[3] ),
    .X(_05122_));
 sky130_fd_sc_hd__xnor2_2 _09112_ (.A(_05112_),
    .B(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__nor2_1 _09113_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B(_05105_),
    .Y(_05124_));
 sky130_fd_sc_hd__o21ba_1 _09114_ (.A1(_05105_),
    .A2(\sbox1.inversion_to_invert_var[0] ),
    .B1_N(_05115_),
    .X(_05125_));
 sky130_fd_sc_hd__a211o_1 _09115_ (.A1(_05105_),
    .A2(\sbox1.inversion_to_invert_var[0] ),
    .B1(\sbox1.inversion_to_invert_var[3] ),
    .C1(\sbox1.inversion_to_invert_var[1] ),
    .X(_05126_));
 sky130_fd_sc_hd__o21a_2 _09116_ (.A1(_05124_),
    .A2(_05125_),
    .B1(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__nand2_1 _09117_ (.A(\sbox1.alph[1] ),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__and2b_1 _09118_ (.A_N(_05105_),
    .B(\sbox1.inversion_to_invert_var[0] ),
    .X(_05129_));
 sky130_fd_sc_hd__o21a_1 _09119_ (.A1(\sbox1.inversion_to_invert_var[1] ),
    .A2(_05105_),
    .B1(\sbox1.inversion_to_invert_var[3] ),
    .X(_05130_));
 sky130_fd_sc_hd__a2111o_1 _09120_ (.A1(_05113_),
    .A2(_05114_),
    .B1(_05117_),
    .C1(_05129_),
    .D1(_05130_),
    .X(_05131_));
 sky130_fd_sc_hd__or3b_1 _09121_ (.A(\sbox1.inversion_to_invert_var[1] ),
    .B(_05105_),
    .C_N(\sbox1.inversion_to_invert_var[3] ),
    .X(_05132_));
 sky130_fd_sc_hd__o221a_1 _09122_ (.A1(\sbox1.inversion_to_invert_var[3] ),
    .A2(_05114_),
    .B1(_05117_),
    .B2(_05129_),
    .C1(_05132_),
    .X(_05133_));
 sky130_fd_sc_hd__a21o_2 _09123_ (.A1(_05119_),
    .A2(_05131_),
    .B1(_05133_),
    .X(_05134_));
 sky130_fd_sc_hd__nand2_1 _09124_ (.A(\sbox1.alph[2] ),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__xnor2_2 _09125_ (.A(_05128_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__xnor2_4 _09126_ (.A(_05123_),
    .B(_05136_),
    .Y(_05137_));
 sky130_fd_sc_hd__nand2_1 _09127_ (.A(\sbox1.ah_reg[1] ),
    .B(_05119_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(\sbox1.ah_reg[3] ),
    .B(_05127_),
    .Y(_05139_));
 sky130_fd_sc_hd__xor2_2 _09129_ (.A(_05138_),
    .B(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__nand2_1 _09130_ (.A(\sbox1.ah_reg[2] ),
    .B(_05111_),
    .Y(_05141_));
 sky130_fd_sc_hd__or2b_1 _09131_ (.A(_05133_),
    .B_N(_05131_),
    .X(_05142_));
 sky130_fd_sc_hd__nand2_1 _09132_ (.A(\sbox1.ah_reg[0] ),
    .B(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__xnor2_2 _09133_ (.A(_05141_),
    .B(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__xnor2_4 _09134_ (.A(_05140_),
    .B(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__nand2_2 _09135_ (.A(\sbox1.alph[0] ),
    .B(_05142_),
    .Y(_05146_));
 sky130_fd_sc_hd__nand2_2 _09136_ (.A(\sbox1.alph[3] ),
    .B(_05127_),
    .Y(_05147_));
 sky130_fd_sc_hd__xor2_4 _09137_ (.A(_05146_),
    .B(_05147_),
    .X(_05148_));
 sky130_fd_sc_hd__nand2_1 _09138_ (.A(\sbox1.alph[1] ),
    .B(_05119_),
    .Y(_05149_));
 sky130_fd_sc_hd__nand2_1 _09139_ (.A(\sbox1.alph[2] ),
    .B(_05111_),
    .Y(_05150_));
 sky130_fd_sc_hd__xnor2_2 _09140_ (.A(_05149_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__xnor2_4 _09141_ (.A(_05148_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__xnor2_4 _09142_ (.A(_05145_),
    .B(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__xnor2_4 _09143_ (.A(_05137_),
    .B(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__and2_1 _09144_ (.A(_05109_),
    .B(_05110_),
    .X(_05155_));
 sky130_fd_sc_hd__o211a_1 _09145_ (.A1(\sbox1.ah_reg[0] ),
    .A2(_05155_),
    .B1(_05119_),
    .C1(\sbox1.ah_reg[3] ),
    .X(_05156_));
 sky130_fd_sc_hd__xnor2_1 _09146_ (.A(\sbox1.ah_reg[0] ),
    .B(\sbox1.ah_reg[3] ),
    .Y(_05157_));
 sky130_fd_sc_hd__a211oi_1 _09147_ (.A1(\sbox1.ah_reg[3] ),
    .A2(_05119_),
    .B1(_05157_),
    .C1(_05155_),
    .Y(_05158_));
 sky130_fd_sc_hd__nor2_2 _09148_ (.A(_05156_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand2_1 _09149_ (.A(\sbox1.ah_reg[1] ),
    .B(_05127_),
    .Y(_05160_));
 sky130_fd_sc_hd__nand2_1 _09150_ (.A(\sbox1.ah_reg[2] ),
    .B(_05134_),
    .Y(_05161_));
 sky130_fd_sc_hd__xnor2_2 _09151_ (.A(_05160_),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__xnor2_4 _09152_ (.A(_05159_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__nand2_2 _09153_ (.A(\sbox1.ah_reg[3] ),
    .B(_05134_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand2_1 _09154_ (.A(\sbox1.ah_reg[0] ),
    .B(_05119_),
    .Y(_05165_));
 sky130_fd_sc_hd__o211a_1 _09155_ (.A1(_05124_),
    .A2(_05125_),
    .B1(_05126_),
    .C1(\sbox1.ah_reg[2] ),
    .X(_05166_));
 sky130_fd_sc_hd__a21bo_1 _09156_ (.A1(_05109_),
    .A2(_05110_),
    .B1_N(\sbox1.ah_reg[1] ),
    .X(_05167_));
 sky130_fd_sc_hd__xnor2_1 _09157_ (.A(_05166_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__xnor2_2 _09158_ (.A(_05165_),
    .B(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__xnor2_4 _09159_ (.A(_05164_),
    .B(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__xor2_4 _09160_ (.A(_05163_),
    .B(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__xnor2_4 _09161_ (.A(_05154_),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__or2_1 _09162_ (.A(\sbox1.ah_reg[3] ),
    .B(\sbox1.ah_reg[2] ),
    .X(_05173_));
 sky130_fd_sc_hd__nand2_1 _09163_ (.A(\sbox1.ah_reg[3] ),
    .B(\sbox1.ah_reg[2] ),
    .Y(_05174_));
 sky130_fd_sc_hd__and3_2 _09164_ (.A(_05111_),
    .B(_05173_),
    .C(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__xor2_1 _09165_ (.A(\sbox1.ah_reg[2] ),
    .B(\sbox1.ah_reg[1] ),
    .X(_05176_));
 sky130_fd_sc_hd__o21ai_2 _09166_ (.A1(_05124_),
    .A2(_05125_),
    .B1(_05126_),
    .Y(_05177_));
 sky130_fd_sc_hd__a211oi_1 _09167_ (.A1(_05119_),
    .A2(_05176_),
    .B1(_05157_),
    .C1(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__o211a_1 _09168_ (.A1(_05177_),
    .A2(_05157_),
    .B1(_05176_),
    .C1(_05119_),
    .X(_05179_));
 sky130_fd_sc_hd__nor2_1 _09169_ (.A(_05178_),
    .B(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__nand2_1 _09170_ (.A(\sbox1.ah_reg[1] ),
    .B(_05142_),
    .Y(_05181_));
 sky130_fd_sc_hd__xnor2_2 _09171_ (.A(_05180_),
    .B(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__xnor2_4 _09172_ (.A(_05175_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__xnor2_4 _09173_ (.A(_05145_),
    .B(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__o21ai_2 _09174_ (.A1(_05120_),
    .A2(_05121_),
    .B1(\sbox1.alph[2] ),
    .Y(_05185_));
 sky130_fd_sc_hd__nand2_1 _09175_ (.A(\sbox1.alph[1] ),
    .B(_05134_),
    .Y(_05186_));
 sky130_fd_sc_hd__xnor2_2 _09176_ (.A(_05185_),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hd__o211ai_1 _09177_ (.A1(\sbox1.alph[0] ),
    .A2(_05177_),
    .B1(_05155_),
    .C1(\sbox1.alph[3] ),
    .Y(_05188_));
 sky130_fd_sc_hd__a211o_1 _09178_ (.A1(\sbox1.alph[3] ),
    .A2(_05155_),
    .B1(_05177_),
    .C1(\sbox1.alph[0] ),
    .X(_05189_));
 sky130_fd_sc_hd__o211a_1 _09179_ (.A1(\sbox1.alph[3] ),
    .A2(_05127_),
    .B1(_05188_),
    .C1(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__xnor2_4 _09180_ (.A(_05187_),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__xor2_2 _09181_ (.A(_05184_),
    .B(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__xnor2_2 _09182_ (.A(_05163_),
    .B(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__inv_2 _09183_ (.A(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__mux2_8 _09184_ (.A0(_05172_),
    .A1(_05194_),
    .S(_05060_),
    .X(_05195_));
 sky130_fd_sc_hd__clkbuf_8 _09185_ (.A(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__nor2_2 _09186_ (.A(_04369_),
    .B(_04946_),
    .Y(_05197_));
 sky130_fd_sc_hd__clkbuf_8 _09187_ (.A(_04617_),
    .X(_05198_));
 sky130_fd_sc_hd__nor2_1 _09188_ (.A(_05198_),
    .B(_04367_),
    .Y(_05199_));
 sky130_fd_sc_hd__clkbuf_4 _09189_ (.A(_05199_),
    .X(_05200_));
 sky130_fd_sc_hd__buf_4 _09190_ (.A(_04624_),
    .X(_05201_));
 sky130_fd_sc_hd__buf_4 _09191_ (.A(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__nor2_1 _09192_ (.A(_05202_),
    .B(_04367_),
    .Y(_05203_));
 sky130_fd_sc_hd__a22o_1 _09193_ (.A1(\sub1.data_o[19] ),
    .A2(_05200_),
    .B1(_05203_),
    .B2(\sub1.data_o[83] ),
    .X(_05204_));
 sky130_fd_sc_hd__a21o_1 _09194_ (.A1(\sub1.data_o[115] ),
    .A2(_05197_),
    .B1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__a31o_1 _09195_ (.A1(_05104_),
    .A2(_04946_),
    .A3(_05196_),
    .B1(_05205_),
    .X(_00000_));
 sky130_fd_sc_hd__nand2_2 _09196_ (.A(\sbox1.alph[3] ),
    .B(_05134_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_1 _09197_ (.A(\sbox1.alph[1] ),
    .B(_05111_),
    .Y(_05207_));
 sky130_fd_sc_hd__nand2_1 _09198_ (.A(\sbox1.alph[0] ),
    .B(_05119_),
    .Y(_05208_));
 sky130_fd_sc_hd__nand2_1 _09199_ (.A(\sbox1.alph[2] ),
    .B(_05127_),
    .Y(_05209_));
 sky130_fd_sc_hd__xor2_1 _09200_ (.A(_05208_),
    .B(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__xnor2_2 _09201_ (.A(_05207_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__xnor2_4 _09202_ (.A(_05206_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__xnor2_2 _09203_ (.A(_05170_),
    .B(_05192_),
    .Y(_05213_));
 sky130_fd_sc_hd__xor2_2 _09204_ (.A(_05212_),
    .B(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__xnor2_4 _09205_ (.A(_05163_),
    .B(_05184_),
    .Y(_05215_));
 sky130_fd_sc_hd__xnor2_2 _09206_ (.A(_05153_),
    .B(_05214_),
    .Y(_05216_));
 sky130_fd_sc_hd__xnor2_4 _09207_ (.A(_05215_),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__mux2_8 _09208_ (.A0(_05214_),
    .A1(_05217_),
    .S(_04649_),
    .X(_05218_));
 sky130_fd_sc_hd__buf_4 _09209_ (.A(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__a22o_1 _09210_ (.A1(\sub1.data_o[20] ),
    .A2(_05200_),
    .B1(_05203_),
    .B2(\sub1.data_o[84] ),
    .X(_05220_));
 sky130_fd_sc_hd__a21o_1 _09211_ (.A1(\sub1.data_o[116] ),
    .A2(_05197_),
    .B1(_05220_),
    .X(_05221_));
 sky130_fd_sc_hd__a31o_1 _09212_ (.A1(_05104_),
    .A2(_04946_),
    .A3(_05219_),
    .B1(_05221_),
    .X(_00001_));
 sky130_fd_sc_hd__xnor2_1 _09213_ (.A(_05170_),
    .B(_05191_),
    .Y(_05222_));
 sky130_fd_sc_hd__xnor2_2 _09214_ (.A(_05137_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__xnor2_4 _09215_ (.A(_05212_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__xnor2_4 _09216_ (.A(_05215_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__xnor2_4 _09217_ (.A(_05137_),
    .B(_05184_),
    .Y(_05226_));
 sky130_fd_sc_hd__mux2_8 _09218_ (.A0(_05225_),
    .A1(_05226_),
    .S(_05060_),
    .X(_05227_));
 sky130_fd_sc_hd__clkbuf_8 _09219_ (.A(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__a22o_1 _09220_ (.A1(\sub1.data_o[21] ),
    .A2(_05200_),
    .B1(_05203_),
    .B2(\sub1.data_o[85] ),
    .X(_05229_));
 sky130_fd_sc_hd__a21o_1 _09221_ (.A1(\sub1.data_o[117] ),
    .A2(_05197_),
    .B1(_05229_),
    .X(_05230_));
 sky130_fd_sc_hd__a31o_1 _09222_ (.A1(_05104_),
    .A2(_04946_),
    .A3(_05228_),
    .B1(_05230_),
    .X(_00002_));
 sky130_fd_sc_hd__nor2_1 _09223_ (.A(_05145_),
    .B(_05171_),
    .Y(_05231_));
 sky130_fd_sc_hd__a21o_1 _09224_ (.A1(_05145_),
    .A2(_05171_),
    .B1(_05060_),
    .X(_05232_));
 sky130_fd_sc_hd__xor2_4 _09225_ (.A(_05145_),
    .B(_05224_),
    .X(_05233_));
 sky130_fd_sc_hd__or2_1 _09226_ (.A(_04649_),
    .B(_05233_),
    .X(_05234_));
 sky130_fd_sc_hd__o21ai_4 _09227_ (.A1(_05231_),
    .A2(_05232_),
    .B1(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__clkbuf_8 _09228_ (.A(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__a22o_1 _09229_ (.A1(\sub1.data_o[22] ),
    .A2(_05200_),
    .B1(_05203_),
    .B2(\sub1.data_o[86] ),
    .X(_05237_));
 sky130_fd_sc_hd__a21o_1 _09230_ (.A1(\sub1.data_o[118] ),
    .A2(_05197_),
    .B1(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__a31o_1 _09231_ (.A1(_05104_),
    .A2(_04946_),
    .A3(_05236_),
    .B1(_05238_),
    .X(_00003_));
 sky130_fd_sc_hd__nor2_1 _09232_ (.A(_05193_),
    .B(_05224_),
    .Y(_05239_));
 sky130_fd_sc_hd__a21o_1 _09233_ (.A1(_05193_),
    .A2(_05224_),
    .B1(_05060_),
    .X(_05240_));
 sky130_fd_sc_hd__o21a_2 _09234_ (.A1(_05239_),
    .A2(_05240_),
    .B1(_05234_),
    .X(_05241_));
 sky130_fd_sc_hd__xnor2_4 _09235_ (.A(_05170_),
    .B(_05226_),
    .Y(_05242_));
 sky130_fd_sc_hd__xnor2_4 _09236_ (.A(_05233_),
    .B(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__xor2_4 _09237_ (.A(_05241_),
    .B(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__buf_6 _09238_ (.A(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__a22o_1 _09239_ (.A1(\sub1.data_o[23] ),
    .A2(_05200_),
    .B1(_05203_),
    .B2(\sub1.data_o[87] ),
    .X(_05246_));
 sky130_fd_sc_hd__a21o_1 _09240_ (.A1(\sub1.data_o[119] ),
    .A2(_05197_),
    .B1(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__a31o_1 _09241_ (.A1(_05104_),
    .A2(_04946_),
    .A3(_05245_),
    .B1(_05247_),
    .X(_00004_));
 sky130_fd_sc_hd__o31a_1 _09242_ (.A1(\ks1.state[1] ),
    .A2(_04723_),
    .A3(_04749_),
    .B1(_04737_),
    .X(_00005_));
 sky130_fd_sc_hd__nand2_1 _09243_ (.A(_04741_),
    .B(_04755_),
    .Y(_00006_));
 sky130_fd_sc_hd__clkbuf_4 _09244_ (.A(net130),
    .X(_05248_));
 sky130_fd_sc_hd__buf_2 _09245_ (.A(\fifo_bank_register.write_ptr[0] ),
    .X(_05249_));
 sky130_fd_sc_hd__buf_2 _09246_ (.A(\fifo_bank_register.write_ptr[1] ),
    .X(_05250_));
 sky130_fd_sc_hd__and3_1 _09247_ (.A(_05249_),
    .B(_05250_),
    .C(\fifo_bank_register.write_ptr[2] ),
    .X(_05251_));
 sky130_fd_sc_hd__a21oi_1 _09248_ (.A1(_05249_),
    .A2(_05250_),
    .B1(\fifo_bank_register.write_ptr[2] ),
    .Y(_05252_));
 sky130_fd_sc_hd__xnor2_2 _09249_ (.A(\fifo_bank_register.write_ptr[0] ),
    .B(\fifo_bank_register.write_ptr[1] ),
    .Y(_05253_));
 sky130_fd_sc_hd__inv_2 _09250_ (.A(\fifo_bank_register.write_ptr[3] ),
    .Y(_05254_));
 sky130_fd_sc_hd__a21o_1 _09251_ (.A1(_05252_),
    .A2(_05253_),
    .B1(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__o21ai_2 _09252_ (.A1(\fifo_bank_register.write_ptr[3] ),
    .A2(_05251_),
    .B1(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__nor2_1 _09253_ (.A(\fifo_bank_register.read_ptr[3] ),
    .B(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__xor2_2 _09254_ (.A(\fifo_bank_register.read_ptr[0] ),
    .B(_05249_),
    .X(_05258_));
 sky130_fd_sc_hd__a21bo_1 _09255_ (.A1(\fifo_bank_register.read_ptr[3] ),
    .A2(_05256_),
    .B1_N(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__mux2_1 _09256_ (.A0(\fifo_bank_register.write_ptr[3] ),
    .A1(_05255_),
    .S(_05253_),
    .X(_05260_));
 sky130_fd_sc_hd__xnor2_1 _09257_ (.A(\fifo_bank_register.read_ptr[1] ),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__buf_2 _09258_ (.A(\fifo_bank_register.read_ptr[2] ),
    .X(_05262_));
 sky130_fd_sc_hd__a21oi_1 _09259_ (.A1(\fifo_bank_register.write_ptr[3] ),
    .A2(_05253_),
    .B1(_05252_),
    .Y(_05263_));
 sky130_fd_sc_hd__mux2_1 _09260_ (.A0(_05263_),
    .A1(\fifo_bank_register.write_ptr[3] ),
    .S(_05251_),
    .X(_05264_));
 sky130_fd_sc_hd__xor2_1 _09261_ (.A(_05262_),
    .B(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__o41a_4 _09262_ (.A1(_05257_),
    .A2(_05259_),
    .A3(_05261_),
    .A4(_05265_),
    .B1(net258),
    .X(_05266_));
 sky130_fd_sc_hd__and3b_1 _09263_ (.A_N(_05250_),
    .B(_05249_),
    .C(net597),
    .X(_05267_));
 sky130_fd_sc_hd__and4b_1 _09264_ (.A_N(\fifo_bank_register.write_ptr[2] ),
    .B(\fifo_bank_register.write_ptr[3] ),
    .C(_05266_),
    .D(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__buf_4 _09265_ (.A(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__clkbuf_4 _09266_ (.A(_05269_),
    .X(_05270_));
 sky130_fd_sc_hd__mux2_1 _09267_ (.A0(\fifo_bank_register.bank[9][0] ),
    .A1(_05248_),
    .S(_05270_),
    .X(_05271_));
 sky130_fd_sc_hd__clkbuf_1 _09268_ (.A(_05271_),
    .X(_00008_));
 sky130_fd_sc_hd__clkbuf_4 _09269_ (.A(net169),
    .X(_05272_));
 sky130_fd_sc_hd__mux2_1 _09270_ (.A0(\fifo_bank_register.bank[9][1] ),
    .A1(_05272_),
    .S(_05270_),
    .X(_05273_));
 sky130_fd_sc_hd__clkbuf_1 _09271_ (.A(_05273_),
    .X(_00009_));
 sky130_fd_sc_hd__buf_2 _09272_ (.A(net180),
    .X(_05274_));
 sky130_fd_sc_hd__mux2_1 _09273_ (.A0(\fifo_bank_register.bank[9][2] ),
    .A1(_05274_),
    .S(_05270_),
    .X(_05275_));
 sky130_fd_sc_hd__clkbuf_1 _09274_ (.A(_05275_),
    .X(_00010_));
 sky130_fd_sc_hd__clkbuf_4 _09275_ (.A(net191),
    .X(_05276_));
 sky130_fd_sc_hd__mux2_1 _09276_ (.A0(\fifo_bank_register.bank[9][3] ),
    .A1(_05276_),
    .S(_05270_),
    .X(_05277_));
 sky130_fd_sc_hd__clkbuf_1 _09277_ (.A(_05277_),
    .X(_00011_));
 sky130_fd_sc_hd__buf_2 _09278_ (.A(net202),
    .X(_05278_));
 sky130_fd_sc_hd__mux2_1 _09279_ (.A0(\fifo_bank_register.bank[9][4] ),
    .A1(_05278_),
    .S(_05270_),
    .X(_05279_));
 sky130_fd_sc_hd__clkbuf_1 _09280_ (.A(_05279_),
    .X(_00012_));
 sky130_fd_sc_hd__buf_2 _09281_ (.A(net213),
    .X(_05280_));
 sky130_fd_sc_hd__mux2_1 _09282_ (.A0(\fifo_bank_register.bank[9][5] ),
    .A1(_05280_),
    .S(_05270_),
    .X(_05281_));
 sky130_fd_sc_hd__clkbuf_1 _09283_ (.A(_05281_),
    .X(_00013_));
 sky130_fd_sc_hd__clkbuf_4 _09284_ (.A(net224),
    .X(_05282_));
 sky130_fd_sc_hd__mux2_1 _09285_ (.A0(\fifo_bank_register.bank[9][6] ),
    .A1(_05282_),
    .S(_05270_),
    .X(_05283_));
 sky130_fd_sc_hd__clkbuf_1 _09286_ (.A(_05283_),
    .X(_00014_));
 sky130_fd_sc_hd__clkbuf_4 _09287_ (.A(net235),
    .X(_05284_));
 sky130_fd_sc_hd__mux2_1 _09288_ (.A0(\fifo_bank_register.bank[9][7] ),
    .A1(_05284_),
    .S(_05270_),
    .X(_05285_));
 sky130_fd_sc_hd__clkbuf_1 _09289_ (.A(_05285_),
    .X(_00015_));
 sky130_fd_sc_hd__clkbuf_4 _09290_ (.A(net246),
    .X(_05286_));
 sky130_fd_sc_hd__mux2_1 _09291_ (.A0(\fifo_bank_register.bank[9][8] ),
    .A1(_05286_),
    .S(_05270_),
    .X(_05287_));
 sky130_fd_sc_hd__clkbuf_1 _09292_ (.A(_05287_),
    .X(_00016_));
 sky130_fd_sc_hd__buf_2 _09293_ (.A(net257),
    .X(_05288_));
 sky130_fd_sc_hd__mux2_1 _09294_ (.A0(\fifo_bank_register.bank[9][9] ),
    .A1(_05288_),
    .S(_05270_),
    .X(_05289_));
 sky130_fd_sc_hd__clkbuf_1 _09295_ (.A(_05289_),
    .X(_00017_));
 sky130_fd_sc_hd__clkbuf_4 _09296_ (.A(net141),
    .X(_05290_));
 sky130_fd_sc_hd__buf_4 _09297_ (.A(_05269_),
    .X(_05291_));
 sky130_fd_sc_hd__mux2_1 _09298_ (.A0(\fifo_bank_register.bank[9][10] ),
    .A1(_05290_),
    .S(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_1 _09299_ (.A(_05292_),
    .X(_00018_));
 sky130_fd_sc_hd__buf_2 _09300_ (.A(net152),
    .X(_05293_));
 sky130_fd_sc_hd__mux2_1 _09301_ (.A0(\fifo_bank_register.bank[9][11] ),
    .A1(_05293_),
    .S(_05291_),
    .X(_05294_));
 sky130_fd_sc_hd__clkbuf_1 _09302_ (.A(_05294_),
    .X(_00019_));
 sky130_fd_sc_hd__buf_2 _09303_ (.A(net161),
    .X(_05295_));
 sky130_fd_sc_hd__mux2_1 _09304_ (.A0(\fifo_bank_register.bank[9][12] ),
    .A1(_05295_),
    .S(_05291_),
    .X(_05296_));
 sky130_fd_sc_hd__clkbuf_1 _09305_ (.A(_05296_),
    .X(_00020_));
 sky130_fd_sc_hd__buf_2 _09306_ (.A(net162),
    .X(_05297_));
 sky130_fd_sc_hd__mux2_1 _09307_ (.A0(\fifo_bank_register.bank[9][13] ),
    .A1(_05297_),
    .S(_05291_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_1 _09308_ (.A(_05298_),
    .X(_00021_));
 sky130_fd_sc_hd__buf_2 _09309_ (.A(net163),
    .X(_05299_));
 sky130_fd_sc_hd__mux2_1 _09310_ (.A0(\fifo_bank_register.bank[9][14] ),
    .A1(_05299_),
    .S(_05291_),
    .X(_05300_));
 sky130_fd_sc_hd__clkbuf_1 _09311_ (.A(_05300_),
    .X(_00022_));
 sky130_fd_sc_hd__buf_2 _09312_ (.A(net164),
    .X(_05301_));
 sky130_fd_sc_hd__mux2_1 _09313_ (.A0(\fifo_bank_register.bank[9][15] ),
    .A1(_05301_),
    .S(_05291_),
    .X(_05302_));
 sky130_fd_sc_hd__clkbuf_1 _09314_ (.A(_05302_),
    .X(_00023_));
 sky130_fd_sc_hd__buf_2 _09315_ (.A(net165),
    .X(_05303_));
 sky130_fd_sc_hd__mux2_1 _09316_ (.A0(\fifo_bank_register.bank[9][16] ),
    .A1(_05303_),
    .S(_05291_),
    .X(_05304_));
 sky130_fd_sc_hd__clkbuf_1 _09317_ (.A(_05304_),
    .X(_00024_));
 sky130_fd_sc_hd__clkbuf_4 _09318_ (.A(net166),
    .X(_05305_));
 sky130_fd_sc_hd__mux2_1 _09319_ (.A0(\fifo_bank_register.bank[9][17] ),
    .A1(_05305_),
    .S(_05291_),
    .X(_05306_));
 sky130_fd_sc_hd__clkbuf_1 _09320_ (.A(_05306_),
    .X(_00025_));
 sky130_fd_sc_hd__buf_2 _09321_ (.A(net167),
    .X(_05307_));
 sky130_fd_sc_hd__mux2_1 _09322_ (.A0(\fifo_bank_register.bank[9][18] ),
    .A1(_05307_),
    .S(_05291_),
    .X(_05308_));
 sky130_fd_sc_hd__clkbuf_1 _09323_ (.A(_05308_),
    .X(_00026_));
 sky130_fd_sc_hd__buf_2 _09324_ (.A(net168),
    .X(_05309_));
 sky130_fd_sc_hd__mux2_1 _09325_ (.A0(\fifo_bank_register.bank[9][19] ),
    .A1(_05309_),
    .S(_05291_),
    .X(_05310_));
 sky130_fd_sc_hd__clkbuf_1 _09326_ (.A(_05310_),
    .X(_00027_));
 sky130_fd_sc_hd__clkbuf_4 _09327_ (.A(net170),
    .X(_05311_));
 sky130_fd_sc_hd__buf_6 _09328_ (.A(_05268_),
    .X(_05312_));
 sky130_fd_sc_hd__buf_4 _09329_ (.A(_05312_),
    .X(_05313_));
 sky130_fd_sc_hd__mux2_1 _09330_ (.A0(\fifo_bank_register.bank[9][20] ),
    .A1(_05311_),
    .S(_05313_),
    .X(_05314_));
 sky130_fd_sc_hd__clkbuf_1 _09331_ (.A(_05314_),
    .X(_00028_));
 sky130_fd_sc_hd__clkbuf_2 _09332_ (.A(net171),
    .X(_05315_));
 sky130_fd_sc_hd__mux2_1 _09333_ (.A0(\fifo_bank_register.bank[9][21] ),
    .A1(_05315_),
    .S(_05313_),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_1 _09334_ (.A(_05316_),
    .X(_00029_));
 sky130_fd_sc_hd__buf_2 _09335_ (.A(net172),
    .X(_05317_));
 sky130_fd_sc_hd__mux2_1 _09336_ (.A0(\fifo_bank_register.bank[9][22] ),
    .A1(_05317_),
    .S(_05313_),
    .X(_05318_));
 sky130_fd_sc_hd__clkbuf_1 _09337_ (.A(_05318_),
    .X(_00030_));
 sky130_fd_sc_hd__buf_2 _09338_ (.A(net173),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _09339_ (.A0(\fifo_bank_register.bank[9][23] ),
    .A1(_05319_),
    .S(_05313_),
    .X(_05320_));
 sky130_fd_sc_hd__clkbuf_1 _09340_ (.A(_05320_),
    .X(_00031_));
 sky130_fd_sc_hd__clkbuf_4 _09341_ (.A(net174),
    .X(_05321_));
 sky130_fd_sc_hd__mux2_1 _09342_ (.A0(\fifo_bank_register.bank[9][24] ),
    .A1(_05321_),
    .S(_05313_),
    .X(_05322_));
 sky130_fd_sc_hd__clkbuf_1 _09343_ (.A(_05322_),
    .X(_00032_));
 sky130_fd_sc_hd__buf_2 _09344_ (.A(net175),
    .X(_05323_));
 sky130_fd_sc_hd__mux2_1 _09345_ (.A0(\fifo_bank_register.bank[9][25] ),
    .A1(_05323_),
    .S(_05313_),
    .X(_05324_));
 sky130_fd_sc_hd__clkbuf_1 _09346_ (.A(_05324_),
    .X(_00033_));
 sky130_fd_sc_hd__buf_2 _09347_ (.A(net176),
    .X(_05325_));
 sky130_fd_sc_hd__mux2_1 _09348_ (.A0(\fifo_bank_register.bank[9][26] ),
    .A1(_05325_),
    .S(_05313_),
    .X(_05326_));
 sky130_fd_sc_hd__clkbuf_1 _09349_ (.A(_05326_),
    .X(_00034_));
 sky130_fd_sc_hd__clkbuf_4 _09350_ (.A(net177),
    .X(_05327_));
 sky130_fd_sc_hd__mux2_1 _09351_ (.A0(\fifo_bank_register.bank[9][27] ),
    .A1(_05327_),
    .S(_05313_),
    .X(_05328_));
 sky130_fd_sc_hd__clkbuf_1 _09352_ (.A(_05328_),
    .X(_00035_));
 sky130_fd_sc_hd__clkbuf_4 _09353_ (.A(net178),
    .X(_05329_));
 sky130_fd_sc_hd__mux2_1 _09354_ (.A0(\fifo_bank_register.bank[9][28] ),
    .A1(_05329_),
    .S(_05313_),
    .X(_05330_));
 sky130_fd_sc_hd__clkbuf_1 _09355_ (.A(_05330_),
    .X(_00036_));
 sky130_fd_sc_hd__buf_2 _09356_ (.A(net179),
    .X(_05331_));
 sky130_fd_sc_hd__mux2_1 _09357_ (.A0(\fifo_bank_register.bank[9][29] ),
    .A1(_05331_),
    .S(_05313_),
    .X(_05332_));
 sky130_fd_sc_hd__clkbuf_1 _09358_ (.A(_05332_),
    .X(_00037_));
 sky130_fd_sc_hd__clkbuf_4 _09359_ (.A(net181),
    .X(_05333_));
 sky130_fd_sc_hd__buf_4 _09360_ (.A(_05312_),
    .X(_05334_));
 sky130_fd_sc_hd__mux2_1 _09361_ (.A0(\fifo_bank_register.bank[9][30] ),
    .A1(_05333_),
    .S(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__clkbuf_1 _09362_ (.A(_05335_),
    .X(_00038_));
 sky130_fd_sc_hd__clkbuf_4 _09363_ (.A(net182),
    .X(_05336_));
 sky130_fd_sc_hd__mux2_1 _09364_ (.A0(\fifo_bank_register.bank[9][31] ),
    .A1(_05336_),
    .S(_05334_),
    .X(_05337_));
 sky130_fd_sc_hd__clkbuf_1 _09365_ (.A(_05337_),
    .X(_00039_));
 sky130_fd_sc_hd__buf_2 _09366_ (.A(net183),
    .X(_05338_));
 sky130_fd_sc_hd__mux2_1 _09367_ (.A0(\fifo_bank_register.bank[9][32] ),
    .A1(_05338_),
    .S(_05334_),
    .X(_05339_));
 sky130_fd_sc_hd__clkbuf_1 _09368_ (.A(_05339_),
    .X(_00040_));
 sky130_fd_sc_hd__clkbuf_4 _09369_ (.A(net184),
    .X(_05340_));
 sky130_fd_sc_hd__mux2_1 _09370_ (.A0(\fifo_bank_register.bank[9][33] ),
    .A1(_05340_),
    .S(_05334_),
    .X(_05341_));
 sky130_fd_sc_hd__clkbuf_1 _09371_ (.A(_05341_),
    .X(_00041_));
 sky130_fd_sc_hd__clkbuf_4 _09372_ (.A(net185),
    .X(_05342_));
 sky130_fd_sc_hd__mux2_1 _09373_ (.A0(\fifo_bank_register.bank[9][34] ),
    .A1(_05342_),
    .S(_05334_),
    .X(_05343_));
 sky130_fd_sc_hd__clkbuf_1 _09374_ (.A(_05343_),
    .X(_00042_));
 sky130_fd_sc_hd__buf_2 _09375_ (.A(net186),
    .X(_05344_));
 sky130_fd_sc_hd__mux2_1 _09376_ (.A0(\fifo_bank_register.bank[9][35] ),
    .A1(_05344_),
    .S(_05334_),
    .X(_05345_));
 sky130_fd_sc_hd__clkbuf_1 _09377_ (.A(_05345_),
    .X(_00043_));
 sky130_fd_sc_hd__buf_2 _09378_ (.A(net187),
    .X(_05346_));
 sky130_fd_sc_hd__mux2_1 _09379_ (.A0(\fifo_bank_register.bank[9][36] ),
    .A1(_05346_),
    .S(_05334_),
    .X(_05347_));
 sky130_fd_sc_hd__clkbuf_1 _09380_ (.A(_05347_),
    .X(_00044_));
 sky130_fd_sc_hd__buf_2 _09381_ (.A(net188),
    .X(_05348_));
 sky130_fd_sc_hd__mux2_1 _09382_ (.A0(\fifo_bank_register.bank[9][37] ),
    .A1(_05348_),
    .S(_05334_),
    .X(_05349_));
 sky130_fd_sc_hd__clkbuf_1 _09383_ (.A(_05349_),
    .X(_00045_));
 sky130_fd_sc_hd__clkbuf_4 _09384_ (.A(net189),
    .X(_05350_));
 sky130_fd_sc_hd__mux2_1 _09385_ (.A0(\fifo_bank_register.bank[9][38] ),
    .A1(_05350_),
    .S(_05334_),
    .X(_05351_));
 sky130_fd_sc_hd__clkbuf_1 _09386_ (.A(_05351_),
    .X(_00046_));
 sky130_fd_sc_hd__clkbuf_4 _09387_ (.A(net190),
    .X(_05352_));
 sky130_fd_sc_hd__mux2_1 _09388_ (.A0(\fifo_bank_register.bank[9][39] ),
    .A1(_05352_),
    .S(_05334_),
    .X(_05353_));
 sky130_fd_sc_hd__clkbuf_1 _09389_ (.A(_05353_),
    .X(_00047_));
 sky130_fd_sc_hd__buf_2 _09390_ (.A(net192),
    .X(_05354_));
 sky130_fd_sc_hd__buf_4 _09391_ (.A(_05312_),
    .X(_05355_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(\fifo_bank_register.bank[9][40] ),
    .A1(_05354_),
    .S(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__clkbuf_1 _09393_ (.A(_05356_),
    .X(_00048_));
 sky130_fd_sc_hd__buf_2 _09394_ (.A(net193),
    .X(_05357_));
 sky130_fd_sc_hd__mux2_1 _09395_ (.A0(\fifo_bank_register.bank[9][41] ),
    .A1(_05357_),
    .S(_05355_),
    .X(_05358_));
 sky130_fd_sc_hd__clkbuf_1 _09396_ (.A(_05358_),
    .X(_00049_));
 sky130_fd_sc_hd__clkbuf_4 _09397_ (.A(net194),
    .X(_05359_));
 sky130_fd_sc_hd__mux2_1 _09398_ (.A0(\fifo_bank_register.bank[9][42] ),
    .A1(_05359_),
    .S(_05355_),
    .X(_05360_));
 sky130_fd_sc_hd__clkbuf_1 _09399_ (.A(_05360_),
    .X(_00050_));
 sky130_fd_sc_hd__buf_2 _09400_ (.A(net195),
    .X(_05361_));
 sky130_fd_sc_hd__mux2_1 _09401_ (.A0(\fifo_bank_register.bank[9][43] ),
    .A1(_05361_),
    .S(_05355_),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_1 _09402_ (.A(_05362_),
    .X(_00051_));
 sky130_fd_sc_hd__buf_2 _09403_ (.A(net196),
    .X(_05363_));
 sky130_fd_sc_hd__mux2_1 _09404_ (.A0(\fifo_bank_register.bank[9][44] ),
    .A1(_05363_),
    .S(_05355_),
    .X(_05364_));
 sky130_fd_sc_hd__clkbuf_1 _09405_ (.A(_05364_),
    .X(_00052_));
 sky130_fd_sc_hd__clkbuf_4 _09406_ (.A(net197),
    .X(_05365_));
 sky130_fd_sc_hd__mux2_1 _09407_ (.A0(\fifo_bank_register.bank[9][45] ),
    .A1(_05365_),
    .S(_05355_),
    .X(_05366_));
 sky130_fd_sc_hd__clkbuf_1 _09408_ (.A(_05366_),
    .X(_00053_));
 sky130_fd_sc_hd__clkbuf_4 _09409_ (.A(net198),
    .X(_05367_));
 sky130_fd_sc_hd__mux2_1 _09410_ (.A0(\fifo_bank_register.bank[9][46] ),
    .A1(_05367_),
    .S(_05355_),
    .X(_05368_));
 sky130_fd_sc_hd__clkbuf_1 _09411_ (.A(_05368_),
    .X(_00054_));
 sky130_fd_sc_hd__buf_4 _09412_ (.A(net199),
    .X(_05369_));
 sky130_fd_sc_hd__mux2_1 _09413_ (.A0(\fifo_bank_register.bank[9][47] ),
    .A1(_05369_),
    .S(_05355_),
    .X(_05370_));
 sky130_fd_sc_hd__clkbuf_1 _09414_ (.A(_05370_),
    .X(_00055_));
 sky130_fd_sc_hd__buf_4 _09415_ (.A(net200),
    .X(_05371_));
 sky130_fd_sc_hd__mux2_1 _09416_ (.A0(\fifo_bank_register.bank[9][48] ),
    .A1(_05371_),
    .S(_05355_),
    .X(_05372_));
 sky130_fd_sc_hd__clkbuf_1 _09417_ (.A(_05372_),
    .X(_00056_));
 sky130_fd_sc_hd__clkbuf_4 _09418_ (.A(net201),
    .X(_05373_));
 sky130_fd_sc_hd__mux2_1 _09419_ (.A0(\fifo_bank_register.bank[9][49] ),
    .A1(_05373_),
    .S(_05355_),
    .X(_05374_));
 sky130_fd_sc_hd__clkbuf_1 _09420_ (.A(_05374_),
    .X(_00057_));
 sky130_fd_sc_hd__buf_2 _09421_ (.A(net203),
    .X(_05375_));
 sky130_fd_sc_hd__buf_4 _09422_ (.A(_05312_),
    .X(_05376_));
 sky130_fd_sc_hd__mux2_1 _09423_ (.A0(\fifo_bank_register.bank[9][50] ),
    .A1(_05375_),
    .S(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__clkbuf_1 _09424_ (.A(_05377_),
    .X(_00058_));
 sky130_fd_sc_hd__buf_2 _09425_ (.A(net204),
    .X(_05378_));
 sky130_fd_sc_hd__mux2_1 _09426_ (.A0(\fifo_bank_register.bank[9][51] ),
    .A1(_05378_),
    .S(_05376_),
    .X(_05379_));
 sky130_fd_sc_hd__clkbuf_1 _09427_ (.A(_05379_),
    .X(_00059_));
 sky130_fd_sc_hd__clkbuf_4 _09428_ (.A(net205),
    .X(_05380_));
 sky130_fd_sc_hd__mux2_1 _09429_ (.A0(\fifo_bank_register.bank[9][52] ),
    .A1(_05380_),
    .S(_05376_),
    .X(_05381_));
 sky130_fd_sc_hd__clkbuf_1 _09430_ (.A(_05381_),
    .X(_00060_));
 sky130_fd_sc_hd__clkbuf_4 _09431_ (.A(net206),
    .X(_05382_));
 sky130_fd_sc_hd__mux2_1 _09432_ (.A0(\fifo_bank_register.bank[9][53] ),
    .A1(_05382_),
    .S(_05376_),
    .X(_05383_));
 sky130_fd_sc_hd__clkbuf_1 _09433_ (.A(_05383_),
    .X(_00061_));
 sky130_fd_sc_hd__buf_2 _09434_ (.A(net207),
    .X(_05384_));
 sky130_fd_sc_hd__mux2_1 _09435_ (.A0(\fifo_bank_register.bank[9][54] ),
    .A1(_05384_),
    .S(_05376_),
    .X(_05385_));
 sky130_fd_sc_hd__clkbuf_1 _09436_ (.A(_05385_),
    .X(_00062_));
 sky130_fd_sc_hd__clkbuf_4 _09437_ (.A(net208),
    .X(_05386_));
 sky130_fd_sc_hd__mux2_1 _09438_ (.A0(\fifo_bank_register.bank[9][55] ),
    .A1(_05386_),
    .S(_05376_),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _09439_ (.A(_05387_),
    .X(_00063_));
 sky130_fd_sc_hd__buf_2 _09440_ (.A(net209),
    .X(_05388_));
 sky130_fd_sc_hd__mux2_1 _09441_ (.A0(\fifo_bank_register.bank[9][56] ),
    .A1(_05388_),
    .S(_05376_),
    .X(_05389_));
 sky130_fd_sc_hd__clkbuf_1 _09442_ (.A(_05389_),
    .X(_00064_));
 sky130_fd_sc_hd__clkbuf_4 _09443_ (.A(net210),
    .X(_05390_));
 sky130_fd_sc_hd__mux2_1 _09444_ (.A0(\fifo_bank_register.bank[9][57] ),
    .A1(_05390_),
    .S(_05376_),
    .X(_05391_));
 sky130_fd_sc_hd__clkbuf_1 _09445_ (.A(_05391_),
    .X(_00065_));
 sky130_fd_sc_hd__clkbuf_4 _09446_ (.A(net211),
    .X(_05392_));
 sky130_fd_sc_hd__mux2_1 _09447_ (.A0(\fifo_bank_register.bank[9][58] ),
    .A1(_05392_),
    .S(_05376_),
    .X(_05393_));
 sky130_fd_sc_hd__clkbuf_1 _09448_ (.A(_05393_),
    .X(_00066_));
 sky130_fd_sc_hd__buf_2 _09449_ (.A(net212),
    .X(_05394_));
 sky130_fd_sc_hd__mux2_1 _09450_ (.A0(\fifo_bank_register.bank[9][59] ),
    .A1(_05394_),
    .S(_05376_),
    .X(_05395_));
 sky130_fd_sc_hd__clkbuf_1 _09451_ (.A(_05395_),
    .X(_00067_));
 sky130_fd_sc_hd__buf_2 _09452_ (.A(net214),
    .X(_05396_));
 sky130_fd_sc_hd__buf_4 _09453_ (.A(_05312_),
    .X(_05397_));
 sky130_fd_sc_hd__mux2_1 _09454_ (.A0(\fifo_bank_register.bank[9][60] ),
    .A1(_05396_),
    .S(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__clkbuf_1 _09455_ (.A(_05398_),
    .X(_00068_));
 sky130_fd_sc_hd__clkbuf_4 _09456_ (.A(net215),
    .X(_05399_));
 sky130_fd_sc_hd__mux2_1 _09457_ (.A0(\fifo_bank_register.bank[9][61] ),
    .A1(_05399_),
    .S(_05397_),
    .X(_05400_));
 sky130_fd_sc_hd__clkbuf_1 _09458_ (.A(_05400_),
    .X(_00069_));
 sky130_fd_sc_hd__buf_2 _09459_ (.A(net216),
    .X(_05401_));
 sky130_fd_sc_hd__mux2_1 _09460_ (.A0(\fifo_bank_register.bank[9][62] ),
    .A1(_05401_),
    .S(_05397_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _09461_ (.A(_05402_),
    .X(_00070_));
 sky130_fd_sc_hd__clkbuf_4 _09462_ (.A(net217),
    .X(_05403_));
 sky130_fd_sc_hd__mux2_1 _09463_ (.A0(\fifo_bank_register.bank[9][63] ),
    .A1(_05403_),
    .S(_05397_),
    .X(_05404_));
 sky130_fd_sc_hd__clkbuf_1 _09464_ (.A(_05404_),
    .X(_00071_));
 sky130_fd_sc_hd__clkbuf_4 _09465_ (.A(net218),
    .X(_05405_));
 sky130_fd_sc_hd__mux2_1 _09466_ (.A0(\fifo_bank_register.bank[9][64] ),
    .A1(_05405_),
    .S(_05397_),
    .X(_05406_));
 sky130_fd_sc_hd__clkbuf_1 _09467_ (.A(_05406_),
    .X(_00072_));
 sky130_fd_sc_hd__buf_2 _09468_ (.A(net219),
    .X(_05407_));
 sky130_fd_sc_hd__mux2_1 _09469_ (.A0(\fifo_bank_register.bank[9][65] ),
    .A1(_05407_),
    .S(_05397_),
    .X(_05408_));
 sky130_fd_sc_hd__clkbuf_1 _09470_ (.A(_05408_),
    .X(_00073_));
 sky130_fd_sc_hd__buf_2 _09471_ (.A(net220),
    .X(_05409_));
 sky130_fd_sc_hd__mux2_1 _09472_ (.A0(\fifo_bank_register.bank[9][66] ),
    .A1(_05409_),
    .S(_05397_),
    .X(_05410_));
 sky130_fd_sc_hd__clkbuf_1 _09473_ (.A(_05410_),
    .X(_00074_));
 sky130_fd_sc_hd__buf_2 _09474_ (.A(net221),
    .X(_05411_));
 sky130_fd_sc_hd__mux2_1 _09475_ (.A0(\fifo_bank_register.bank[9][67] ),
    .A1(_05411_),
    .S(_05397_),
    .X(_05412_));
 sky130_fd_sc_hd__clkbuf_1 _09476_ (.A(_05412_),
    .X(_00075_));
 sky130_fd_sc_hd__buf_2 _09477_ (.A(net222),
    .X(_05413_));
 sky130_fd_sc_hd__mux2_1 _09478_ (.A0(\fifo_bank_register.bank[9][68] ),
    .A1(_05413_),
    .S(_05397_),
    .X(_05414_));
 sky130_fd_sc_hd__clkbuf_1 _09479_ (.A(_05414_),
    .X(_00076_));
 sky130_fd_sc_hd__clkbuf_4 _09480_ (.A(net223),
    .X(_05415_));
 sky130_fd_sc_hd__mux2_1 _09481_ (.A0(\fifo_bank_register.bank[9][69] ),
    .A1(_05415_),
    .S(_05397_),
    .X(_05416_));
 sky130_fd_sc_hd__clkbuf_1 _09482_ (.A(_05416_),
    .X(_00077_));
 sky130_fd_sc_hd__clkbuf_4 _09483_ (.A(net225),
    .X(_05417_));
 sky130_fd_sc_hd__buf_4 _09484_ (.A(_05312_),
    .X(_05418_));
 sky130_fd_sc_hd__mux2_1 _09485_ (.A0(\fifo_bank_register.bank[9][70] ),
    .A1(_05417_),
    .S(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__clkbuf_1 _09486_ (.A(_05419_),
    .X(_00078_));
 sky130_fd_sc_hd__buf_2 _09487_ (.A(net226),
    .X(_05420_));
 sky130_fd_sc_hd__mux2_1 _09488_ (.A0(\fifo_bank_register.bank[9][71] ),
    .A1(_05420_),
    .S(_05418_),
    .X(_05421_));
 sky130_fd_sc_hd__clkbuf_1 _09489_ (.A(_05421_),
    .X(_00079_));
 sky130_fd_sc_hd__buf_2 _09490_ (.A(net227),
    .X(_05422_));
 sky130_fd_sc_hd__mux2_1 _09491_ (.A0(\fifo_bank_register.bank[9][72] ),
    .A1(_05422_),
    .S(_05418_),
    .X(_05423_));
 sky130_fd_sc_hd__clkbuf_1 _09492_ (.A(_05423_),
    .X(_00080_));
 sky130_fd_sc_hd__buf_2 _09493_ (.A(net228),
    .X(_05424_));
 sky130_fd_sc_hd__mux2_1 _09494_ (.A0(\fifo_bank_register.bank[9][73] ),
    .A1(_05424_),
    .S(_05418_),
    .X(_05425_));
 sky130_fd_sc_hd__clkbuf_1 _09495_ (.A(_05425_),
    .X(_00081_));
 sky130_fd_sc_hd__buf_2 _09496_ (.A(net229),
    .X(_05426_));
 sky130_fd_sc_hd__mux2_1 _09497_ (.A0(\fifo_bank_register.bank[9][74] ),
    .A1(_05426_),
    .S(_05418_),
    .X(_05427_));
 sky130_fd_sc_hd__clkbuf_1 _09498_ (.A(_05427_),
    .X(_00082_));
 sky130_fd_sc_hd__clkbuf_4 _09499_ (.A(net230),
    .X(_05428_));
 sky130_fd_sc_hd__mux2_1 _09500_ (.A0(\fifo_bank_register.bank[9][75] ),
    .A1(_05428_),
    .S(_05418_),
    .X(_05429_));
 sky130_fd_sc_hd__clkbuf_1 _09501_ (.A(_05429_),
    .X(_00083_));
 sky130_fd_sc_hd__clkbuf_4 _09502_ (.A(net231),
    .X(_05430_));
 sky130_fd_sc_hd__mux2_1 _09503_ (.A0(\fifo_bank_register.bank[9][76] ),
    .A1(_05430_),
    .S(_05418_),
    .X(_05431_));
 sky130_fd_sc_hd__clkbuf_1 _09504_ (.A(_05431_),
    .X(_00084_));
 sky130_fd_sc_hd__clkbuf_4 _09505_ (.A(net232),
    .X(_05432_));
 sky130_fd_sc_hd__mux2_1 _09506_ (.A0(\fifo_bank_register.bank[9][77] ),
    .A1(_05432_),
    .S(_05418_),
    .X(_05433_));
 sky130_fd_sc_hd__clkbuf_1 _09507_ (.A(_05433_),
    .X(_00085_));
 sky130_fd_sc_hd__clkbuf_4 _09508_ (.A(net233),
    .X(_05434_));
 sky130_fd_sc_hd__mux2_1 _09509_ (.A0(\fifo_bank_register.bank[9][78] ),
    .A1(_05434_),
    .S(_05418_),
    .X(_05435_));
 sky130_fd_sc_hd__clkbuf_1 _09510_ (.A(_05435_),
    .X(_00086_));
 sky130_fd_sc_hd__buf_2 _09511_ (.A(net234),
    .X(_05436_));
 sky130_fd_sc_hd__mux2_1 _09512_ (.A0(\fifo_bank_register.bank[9][79] ),
    .A1(_05436_),
    .S(_05418_),
    .X(_05437_));
 sky130_fd_sc_hd__clkbuf_1 _09513_ (.A(_05437_),
    .X(_00087_));
 sky130_fd_sc_hd__clkbuf_4 _09514_ (.A(net236),
    .X(_05438_));
 sky130_fd_sc_hd__buf_4 _09515_ (.A(_05312_),
    .X(_05439_));
 sky130_fd_sc_hd__mux2_1 _09516_ (.A0(\fifo_bank_register.bank[9][80] ),
    .A1(_05438_),
    .S(_05439_),
    .X(_05440_));
 sky130_fd_sc_hd__clkbuf_1 _09517_ (.A(_05440_),
    .X(_00088_));
 sky130_fd_sc_hd__clkbuf_4 _09518_ (.A(net237),
    .X(_05441_));
 sky130_fd_sc_hd__mux2_1 _09519_ (.A0(\fifo_bank_register.bank[9][81] ),
    .A1(_05441_),
    .S(_05439_),
    .X(_05442_));
 sky130_fd_sc_hd__clkbuf_1 _09520_ (.A(_05442_),
    .X(_00089_));
 sky130_fd_sc_hd__clkbuf_4 _09521_ (.A(net238),
    .X(_05443_));
 sky130_fd_sc_hd__mux2_1 _09522_ (.A0(\fifo_bank_register.bank[9][82] ),
    .A1(_05443_),
    .S(_05439_),
    .X(_05444_));
 sky130_fd_sc_hd__clkbuf_1 _09523_ (.A(_05444_),
    .X(_00090_));
 sky130_fd_sc_hd__clkbuf_4 _09524_ (.A(net239),
    .X(_05445_));
 sky130_fd_sc_hd__mux2_1 _09525_ (.A0(\fifo_bank_register.bank[9][83] ),
    .A1(_05445_),
    .S(_05439_),
    .X(_05446_));
 sky130_fd_sc_hd__clkbuf_1 _09526_ (.A(_05446_),
    .X(_00091_));
 sky130_fd_sc_hd__clkbuf_4 _09527_ (.A(net240),
    .X(_05447_));
 sky130_fd_sc_hd__mux2_1 _09528_ (.A0(\fifo_bank_register.bank[9][84] ),
    .A1(_05447_),
    .S(_05439_),
    .X(_05448_));
 sky130_fd_sc_hd__clkbuf_1 _09529_ (.A(_05448_),
    .X(_00092_));
 sky130_fd_sc_hd__clkbuf_4 _09530_ (.A(net241),
    .X(_05449_));
 sky130_fd_sc_hd__mux2_1 _09531_ (.A0(\fifo_bank_register.bank[9][85] ),
    .A1(_05449_),
    .S(_05439_),
    .X(_05450_));
 sky130_fd_sc_hd__clkbuf_1 _09532_ (.A(_05450_),
    .X(_00093_));
 sky130_fd_sc_hd__clkbuf_4 _09533_ (.A(net242),
    .X(_05451_));
 sky130_fd_sc_hd__mux2_1 _09534_ (.A0(\fifo_bank_register.bank[9][86] ),
    .A1(_05451_),
    .S(_05439_),
    .X(_05452_));
 sky130_fd_sc_hd__clkbuf_1 _09535_ (.A(_05452_),
    .X(_00094_));
 sky130_fd_sc_hd__clkbuf_4 _09536_ (.A(net243),
    .X(_05453_));
 sky130_fd_sc_hd__mux2_1 _09537_ (.A0(\fifo_bank_register.bank[9][87] ),
    .A1(_05453_),
    .S(_05439_),
    .X(_05454_));
 sky130_fd_sc_hd__clkbuf_1 _09538_ (.A(_05454_),
    .X(_00095_));
 sky130_fd_sc_hd__buf_2 _09539_ (.A(net244),
    .X(_05455_));
 sky130_fd_sc_hd__mux2_1 _09540_ (.A0(\fifo_bank_register.bank[9][88] ),
    .A1(_05455_),
    .S(_05439_),
    .X(_05456_));
 sky130_fd_sc_hd__clkbuf_1 _09541_ (.A(_05456_),
    .X(_00096_));
 sky130_fd_sc_hd__buf_2 _09542_ (.A(net245),
    .X(_05457_));
 sky130_fd_sc_hd__mux2_1 _09543_ (.A0(\fifo_bank_register.bank[9][89] ),
    .A1(_05457_),
    .S(_05439_),
    .X(_05458_));
 sky130_fd_sc_hd__clkbuf_1 _09544_ (.A(_05458_),
    .X(_00097_));
 sky130_fd_sc_hd__clkbuf_4 _09545_ (.A(net247),
    .X(_05459_));
 sky130_fd_sc_hd__buf_4 _09546_ (.A(_05312_),
    .X(_05460_));
 sky130_fd_sc_hd__mux2_1 _09547_ (.A0(\fifo_bank_register.bank[9][90] ),
    .A1(_05459_),
    .S(_05460_),
    .X(_05461_));
 sky130_fd_sc_hd__clkbuf_1 _09548_ (.A(_05461_),
    .X(_00098_));
 sky130_fd_sc_hd__buf_2 _09549_ (.A(net248),
    .X(_05462_));
 sky130_fd_sc_hd__mux2_1 _09550_ (.A0(\fifo_bank_register.bank[9][91] ),
    .A1(_05462_),
    .S(_05460_),
    .X(_05463_));
 sky130_fd_sc_hd__clkbuf_1 _09551_ (.A(_05463_),
    .X(_00099_));
 sky130_fd_sc_hd__buf_2 _09552_ (.A(net249),
    .X(_05464_));
 sky130_fd_sc_hd__mux2_1 _09553_ (.A0(\fifo_bank_register.bank[9][92] ),
    .A1(_05464_),
    .S(_05460_),
    .X(_05465_));
 sky130_fd_sc_hd__clkbuf_1 _09554_ (.A(_05465_),
    .X(_00100_));
 sky130_fd_sc_hd__buf_2 _09555_ (.A(net250),
    .X(_05466_));
 sky130_fd_sc_hd__mux2_1 _09556_ (.A0(\fifo_bank_register.bank[9][93] ),
    .A1(_05466_),
    .S(_05460_),
    .X(_05467_));
 sky130_fd_sc_hd__clkbuf_1 _09557_ (.A(_05467_),
    .X(_00101_));
 sky130_fd_sc_hd__clkbuf_4 _09558_ (.A(net251),
    .X(_05468_));
 sky130_fd_sc_hd__mux2_1 _09559_ (.A0(\fifo_bank_register.bank[9][94] ),
    .A1(_05468_),
    .S(_05460_),
    .X(_05469_));
 sky130_fd_sc_hd__clkbuf_1 _09560_ (.A(_05469_),
    .X(_00102_));
 sky130_fd_sc_hd__clkbuf_4 _09561_ (.A(net252),
    .X(_05470_));
 sky130_fd_sc_hd__mux2_1 _09562_ (.A0(\fifo_bank_register.bank[9][95] ),
    .A1(_05470_),
    .S(_05460_),
    .X(_05471_));
 sky130_fd_sc_hd__clkbuf_1 _09563_ (.A(_05471_),
    .X(_00103_));
 sky130_fd_sc_hd__clkbuf_4 _09564_ (.A(net253),
    .X(_05472_));
 sky130_fd_sc_hd__mux2_1 _09565_ (.A0(\fifo_bank_register.bank[9][96] ),
    .A1(_05472_),
    .S(_05460_),
    .X(_05473_));
 sky130_fd_sc_hd__clkbuf_1 _09566_ (.A(_05473_),
    .X(_00104_));
 sky130_fd_sc_hd__buf_2 _09567_ (.A(net254),
    .X(_05474_));
 sky130_fd_sc_hd__mux2_1 _09568_ (.A0(\fifo_bank_register.bank[9][97] ),
    .A1(_05474_),
    .S(_05460_),
    .X(_05475_));
 sky130_fd_sc_hd__clkbuf_1 _09569_ (.A(_05475_),
    .X(_00105_));
 sky130_fd_sc_hd__buf_2 _09570_ (.A(net255),
    .X(_05476_));
 sky130_fd_sc_hd__mux2_1 _09571_ (.A0(\fifo_bank_register.bank[9][98] ),
    .A1(_05476_),
    .S(_05460_),
    .X(_05477_));
 sky130_fd_sc_hd__clkbuf_1 _09572_ (.A(_05477_),
    .X(_00106_));
 sky130_fd_sc_hd__buf_2 _09573_ (.A(net256),
    .X(_05478_));
 sky130_fd_sc_hd__mux2_1 _09574_ (.A0(\fifo_bank_register.bank[9][99] ),
    .A1(_05478_),
    .S(_05460_),
    .X(_05479_));
 sky130_fd_sc_hd__clkbuf_1 _09575_ (.A(_05479_),
    .X(_00107_));
 sky130_fd_sc_hd__buf_2 _09576_ (.A(net131),
    .X(_05480_));
 sky130_fd_sc_hd__buf_4 _09577_ (.A(_05312_),
    .X(_05481_));
 sky130_fd_sc_hd__mux2_1 _09578_ (.A0(\fifo_bank_register.bank[9][100] ),
    .A1(_05480_),
    .S(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__clkbuf_1 _09579_ (.A(_05482_),
    .X(_00108_));
 sky130_fd_sc_hd__buf_2 _09580_ (.A(net132),
    .X(_05483_));
 sky130_fd_sc_hd__mux2_1 _09581_ (.A0(\fifo_bank_register.bank[9][101] ),
    .A1(_05483_),
    .S(_05481_),
    .X(_05484_));
 sky130_fd_sc_hd__clkbuf_1 _09582_ (.A(_05484_),
    .X(_00109_));
 sky130_fd_sc_hd__buf_2 _09583_ (.A(net133),
    .X(_05485_));
 sky130_fd_sc_hd__mux2_1 _09584_ (.A0(\fifo_bank_register.bank[9][102] ),
    .A1(_05485_),
    .S(_05481_),
    .X(_05486_));
 sky130_fd_sc_hd__clkbuf_1 _09585_ (.A(_05486_),
    .X(_00110_));
 sky130_fd_sc_hd__buf_2 _09586_ (.A(net134),
    .X(_05487_));
 sky130_fd_sc_hd__mux2_1 _09587_ (.A0(\fifo_bank_register.bank[9][103] ),
    .A1(_05487_),
    .S(_05481_),
    .X(_05488_));
 sky130_fd_sc_hd__clkbuf_1 _09588_ (.A(_05488_),
    .X(_00111_));
 sky130_fd_sc_hd__buf_2 _09589_ (.A(net135),
    .X(_05489_));
 sky130_fd_sc_hd__mux2_1 _09590_ (.A0(\fifo_bank_register.bank[9][104] ),
    .A1(_05489_),
    .S(_05481_),
    .X(_05490_));
 sky130_fd_sc_hd__clkbuf_1 _09591_ (.A(_05490_),
    .X(_00112_));
 sky130_fd_sc_hd__buf_2 _09592_ (.A(net136),
    .X(_05491_));
 sky130_fd_sc_hd__mux2_1 _09593_ (.A0(\fifo_bank_register.bank[9][105] ),
    .A1(_05491_),
    .S(_05481_),
    .X(_05492_));
 sky130_fd_sc_hd__clkbuf_1 _09594_ (.A(_05492_),
    .X(_00113_));
 sky130_fd_sc_hd__buf_2 _09595_ (.A(net137),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_1 _09596_ (.A0(\fifo_bank_register.bank[9][106] ),
    .A1(_05493_),
    .S(_05481_),
    .X(_05494_));
 sky130_fd_sc_hd__clkbuf_1 _09597_ (.A(_05494_),
    .X(_00114_));
 sky130_fd_sc_hd__buf_2 _09598_ (.A(net138),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _09599_ (.A0(\fifo_bank_register.bank[9][107] ),
    .A1(_05495_),
    .S(_05481_),
    .X(_05496_));
 sky130_fd_sc_hd__clkbuf_1 _09600_ (.A(_05496_),
    .X(_00115_));
 sky130_fd_sc_hd__buf_2 _09601_ (.A(net139),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _09602_ (.A0(\fifo_bank_register.bank[9][108] ),
    .A1(_05497_),
    .S(_05481_),
    .X(_05498_));
 sky130_fd_sc_hd__clkbuf_1 _09603_ (.A(_05498_),
    .X(_00116_));
 sky130_fd_sc_hd__buf_2 _09604_ (.A(net140),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _09605_ (.A0(\fifo_bank_register.bank[9][109] ),
    .A1(_05499_),
    .S(_05481_),
    .X(_05500_));
 sky130_fd_sc_hd__clkbuf_1 _09606_ (.A(_05500_),
    .X(_00117_));
 sky130_fd_sc_hd__buf_2 _09607_ (.A(net142),
    .X(_05501_));
 sky130_fd_sc_hd__buf_4 _09608_ (.A(_05312_),
    .X(_05502_));
 sky130_fd_sc_hd__mux2_1 _09609_ (.A0(\fifo_bank_register.bank[9][110] ),
    .A1(_05501_),
    .S(_05502_),
    .X(_05503_));
 sky130_fd_sc_hd__clkbuf_1 _09610_ (.A(_05503_),
    .X(_00118_));
 sky130_fd_sc_hd__buf_2 _09611_ (.A(net143),
    .X(_05504_));
 sky130_fd_sc_hd__mux2_1 _09612_ (.A0(\fifo_bank_register.bank[9][111] ),
    .A1(_05504_),
    .S(_05502_),
    .X(_05505_));
 sky130_fd_sc_hd__clkbuf_1 _09613_ (.A(_05505_),
    .X(_00119_));
 sky130_fd_sc_hd__buf_2 _09614_ (.A(net144),
    .X(_05506_));
 sky130_fd_sc_hd__mux2_1 _09615_ (.A0(\fifo_bank_register.bank[9][112] ),
    .A1(_05506_),
    .S(_05502_),
    .X(_05507_));
 sky130_fd_sc_hd__clkbuf_1 _09616_ (.A(_05507_),
    .X(_00120_));
 sky130_fd_sc_hd__buf_2 _09617_ (.A(net145),
    .X(_05508_));
 sky130_fd_sc_hd__mux2_1 _09618_ (.A0(\fifo_bank_register.bank[9][113] ),
    .A1(_05508_),
    .S(_05502_),
    .X(_05509_));
 sky130_fd_sc_hd__clkbuf_1 _09619_ (.A(_05509_),
    .X(_00121_));
 sky130_fd_sc_hd__buf_2 _09620_ (.A(net146),
    .X(_05510_));
 sky130_fd_sc_hd__mux2_1 _09621_ (.A0(\fifo_bank_register.bank[9][114] ),
    .A1(_05510_),
    .S(_05502_),
    .X(_05511_));
 sky130_fd_sc_hd__clkbuf_1 _09622_ (.A(_05511_),
    .X(_00122_));
 sky130_fd_sc_hd__buf_2 _09623_ (.A(net147),
    .X(_05512_));
 sky130_fd_sc_hd__mux2_1 _09624_ (.A0(\fifo_bank_register.bank[9][115] ),
    .A1(_05512_),
    .S(_05502_),
    .X(_05513_));
 sky130_fd_sc_hd__clkbuf_1 _09625_ (.A(_05513_),
    .X(_00123_));
 sky130_fd_sc_hd__buf_2 _09626_ (.A(net148),
    .X(_05514_));
 sky130_fd_sc_hd__mux2_1 _09627_ (.A0(\fifo_bank_register.bank[9][116] ),
    .A1(_05514_),
    .S(_05502_),
    .X(_05515_));
 sky130_fd_sc_hd__clkbuf_1 _09628_ (.A(_05515_),
    .X(_00124_));
 sky130_fd_sc_hd__buf_2 _09629_ (.A(net149),
    .X(_05516_));
 sky130_fd_sc_hd__mux2_1 _09630_ (.A0(\fifo_bank_register.bank[9][117] ),
    .A1(_05516_),
    .S(_05502_),
    .X(_05517_));
 sky130_fd_sc_hd__clkbuf_1 _09631_ (.A(_05517_),
    .X(_00125_));
 sky130_fd_sc_hd__clkbuf_4 _09632_ (.A(net150),
    .X(_05518_));
 sky130_fd_sc_hd__mux2_1 _09633_ (.A0(\fifo_bank_register.bank[9][118] ),
    .A1(_05518_),
    .S(_05502_),
    .X(_05519_));
 sky130_fd_sc_hd__clkbuf_1 _09634_ (.A(_05519_),
    .X(_00126_));
 sky130_fd_sc_hd__clkbuf_4 _09635_ (.A(net151),
    .X(_05520_));
 sky130_fd_sc_hd__mux2_1 _09636_ (.A0(\fifo_bank_register.bank[9][119] ),
    .A1(_05520_),
    .S(_05502_),
    .X(_05521_));
 sky130_fd_sc_hd__clkbuf_1 _09637_ (.A(_05521_),
    .X(_00127_));
 sky130_fd_sc_hd__clkbuf_4 _09638_ (.A(net153),
    .X(_05522_));
 sky130_fd_sc_hd__mux2_1 _09639_ (.A0(\fifo_bank_register.bank[9][120] ),
    .A1(_05522_),
    .S(_05269_),
    .X(_05523_));
 sky130_fd_sc_hd__clkbuf_1 _09640_ (.A(_05523_),
    .X(_00128_));
 sky130_fd_sc_hd__buf_4 _09641_ (.A(net154),
    .X(_05524_));
 sky130_fd_sc_hd__mux2_1 _09642_ (.A0(\fifo_bank_register.bank[9][121] ),
    .A1(_05524_),
    .S(_05269_),
    .X(_05525_));
 sky130_fd_sc_hd__clkbuf_1 _09643_ (.A(_05525_),
    .X(_00129_));
 sky130_fd_sc_hd__clkbuf_2 _09644_ (.A(net155),
    .X(_05526_));
 sky130_fd_sc_hd__mux2_1 _09645_ (.A0(\fifo_bank_register.bank[9][122] ),
    .A1(_05526_),
    .S(_05269_),
    .X(_05527_));
 sky130_fd_sc_hd__clkbuf_1 _09646_ (.A(_05527_),
    .X(_00130_));
 sky130_fd_sc_hd__clkbuf_4 _09647_ (.A(net156),
    .X(_05528_));
 sky130_fd_sc_hd__mux2_1 _09648_ (.A0(\fifo_bank_register.bank[9][123] ),
    .A1(_05528_),
    .S(_05269_),
    .X(_05529_));
 sky130_fd_sc_hd__clkbuf_1 _09649_ (.A(_05529_),
    .X(_00131_));
 sky130_fd_sc_hd__clkbuf_4 _09650_ (.A(net157),
    .X(_05530_));
 sky130_fd_sc_hd__mux2_1 _09651_ (.A0(\fifo_bank_register.bank[9][124] ),
    .A1(_05530_),
    .S(_05269_),
    .X(_05531_));
 sky130_fd_sc_hd__clkbuf_1 _09652_ (.A(_05531_),
    .X(_00132_));
 sky130_fd_sc_hd__clkbuf_4 _09653_ (.A(net158),
    .X(_05532_));
 sky130_fd_sc_hd__mux2_1 _09654_ (.A0(\fifo_bank_register.bank[9][125] ),
    .A1(_05532_),
    .S(_05269_),
    .X(_05533_));
 sky130_fd_sc_hd__clkbuf_1 _09655_ (.A(_05533_),
    .X(_00133_));
 sky130_fd_sc_hd__clkbuf_4 _09656_ (.A(net159),
    .X(_05534_));
 sky130_fd_sc_hd__mux2_1 _09657_ (.A0(\fifo_bank_register.bank[9][126] ),
    .A1(_05534_),
    .S(_05269_),
    .X(_05535_));
 sky130_fd_sc_hd__clkbuf_1 _09658_ (.A(_05535_),
    .X(_00134_));
 sky130_fd_sc_hd__clkbuf_4 _09659_ (.A(net160),
    .X(_05536_));
 sky130_fd_sc_hd__mux2_1 _09660_ (.A0(\fifo_bank_register.bank[9][127] ),
    .A1(_05536_),
    .S(_05269_),
    .X(_05537_));
 sky130_fd_sc_hd__clkbuf_1 _09661_ (.A(_05537_),
    .X(_00135_));
 sky130_fd_sc_hd__nor2_1 _09662_ (.A(\addroundkey_round[0] ),
    .B(_04644_),
    .Y(_05538_));
 sky130_fd_sc_hd__a211o_1 _09663_ (.A1(\addroundkey_round[0] ),
    .A2(_04637_),
    .B1(_04723_),
    .C1(_05538_),
    .X(_00136_));
 sky130_fd_sc_hd__xor2_1 _09664_ (.A(\addroundkey_round[0] ),
    .B(\addroundkey_round[1] ),
    .X(_05539_));
 sky130_fd_sc_hd__a32o_1 _09665_ (.A1(\addroundkey_round[1] ),
    .A2(_04637_),
    .A3(_04642_),
    .B1(_04749_),
    .B2(_05539_),
    .X(_00137_));
 sky130_fd_sc_hd__and3_1 _09666_ (.A(\addroundkey_round[0] ),
    .B(\addroundkey_round[1] ),
    .C(\addroundkey_round[2] ),
    .X(_05540_));
 sky130_fd_sc_hd__a21oi_1 _09667_ (.A1(\addroundkey_round[0] ),
    .A2(\addroundkey_round[1] ),
    .B1(\addroundkey_round[2] ),
    .Y(_05541_));
 sky130_fd_sc_hd__nor3_2 _09668_ (.A(_04644_),
    .B(_05540_),
    .C(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__a31o_1 _09669_ (.A1(\addroundkey_round[2] ),
    .A2(_04637_),
    .A3(_04642_),
    .B1(_05542_),
    .X(_00138_));
 sky130_fd_sc_hd__xnor2_1 _09670_ (.A(\addroundkey_round[3] ),
    .B(_05540_),
    .Y(_05543_));
 sky130_fd_sc_hd__nor2_1 _09671_ (.A(_04644_),
    .B(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__a31o_1 _09672_ (.A1(\addroundkey_round[3] ),
    .A2(_04637_),
    .A3(_04642_),
    .B1(_05544_),
    .X(_00139_));
 sky130_fd_sc_hd__or2_1 _09673_ (.A(_05152_),
    .B(_05242_),
    .X(_05545_));
 sky130_fd_sc_hd__a21oi_1 _09674_ (.A1(_05152_),
    .A2(_05242_),
    .B1(_05060_),
    .Y(_05546_));
 sky130_fd_sc_hd__a2bb2o_4 _09675_ (.A1_N(_04649_),
    .A2_N(_05153_),
    .B1(_05545_),
    .B2(_05546_),
    .X(_05547_));
 sky130_fd_sc_hd__buf_4 _09676_ (.A(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__mux2_1 _09677_ (.A0(\sub1.data_o[120] ),
    .A1(_05548_),
    .S(_04891_),
    .X(_05549_));
 sky130_fd_sc_hd__clkbuf_1 _09678_ (.A(_05549_),
    .X(_00140_));
 sky130_fd_sc_hd__nor2_1 _09679_ (.A(_05154_),
    .B(_05243_),
    .Y(_05550_));
 sky130_fd_sc_hd__a21o_1 _09680_ (.A1(_05154_),
    .A2(_05243_),
    .B1(_05060_),
    .X(_05551_));
 sky130_fd_sc_hd__o22a_2 _09681_ (.A1(_04649_),
    .A2(_05184_),
    .B1(_05550_),
    .B2(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__xnor2_4 _09682_ (.A(_05170_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__buf_4 _09683_ (.A(_05553_),
    .X(_05554_));
 sky130_fd_sc_hd__mux2_1 _09684_ (.A0(\sub1.data_o[121] ),
    .A1(_05554_),
    .S(_04891_),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_1 _09685_ (.A(_05555_),
    .X(_00141_));
 sky130_fd_sc_hd__xnor2_1 _09686_ (.A(_05153_),
    .B(_05243_),
    .Y(_05556_));
 sky130_fd_sc_hd__xnor2_1 _09687_ (.A(_05191_),
    .B(_05556_),
    .Y(_05557_));
 sky130_fd_sc_hd__mux2_1 _09688_ (.A0(_05213_),
    .A1(_05557_),
    .S(_04649_),
    .X(_05558_));
 sky130_fd_sc_hd__buf_6 _09689_ (.A(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__buf_4 _09690_ (.A(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__mux2_1 _09691_ (.A0(\sub1.data_o[122] ),
    .A1(_05560_),
    .S(_04891_),
    .X(_05561_));
 sky130_fd_sc_hd__clkbuf_1 _09692_ (.A(_05561_),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _09693_ (.A0(\sub1.data_o[123] ),
    .A1(_05196_),
    .S(_04891_),
    .X(_05562_));
 sky130_fd_sc_hd__clkbuf_1 _09694_ (.A(_05562_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _09695_ (.A0(\sub1.data_o[124] ),
    .A1(_05219_),
    .S(_04891_),
    .X(_05563_));
 sky130_fd_sc_hd__clkbuf_1 _09696_ (.A(_05563_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _09697_ (.A0(\sub1.data_o[125] ),
    .A1(_05228_),
    .S(_04891_),
    .X(_05564_));
 sky130_fd_sc_hd__clkbuf_1 _09698_ (.A(_05564_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _09699_ (.A0(\sub1.data_o[126] ),
    .A1(_05236_),
    .S(_04891_),
    .X(_05565_));
 sky130_fd_sc_hd__clkbuf_1 _09700_ (.A(_05565_),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _09701_ (.A0(\sub1.data_o[127] ),
    .A1(_05245_),
    .S(_04891_),
    .X(_05566_));
 sky130_fd_sc_hd__clkbuf_1 _09702_ (.A(_05566_),
    .X(_00147_));
 sky130_fd_sc_hd__buf_4 _09703_ (.A(_04609_),
    .X(_05567_));
 sky130_fd_sc_hd__clkbuf_4 _09704_ (.A(_05567_),
    .X(_05568_));
 sky130_fd_sc_hd__a31o_1 _09705_ (.A1(addroundkey_ready_o),
    .A2(_05568_),
    .A3(_04618_),
    .B1(net388),
    .X(_05569_));
 sky130_fd_sc_hd__and2b_1 _09706_ (.A_N(net258),
    .B(_05569_),
    .X(_05570_));
 sky130_fd_sc_hd__clkbuf_1 _09707_ (.A(_05570_),
    .X(_00148_));
 sky130_fd_sc_hd__nand2_1 _09708_ (.A(_05198_),
    .B(_04629_),
    .Y(_05571_));
 sky130_fd_sc_hd__xor2_1 _09709_ (.A(_04613_),
    .B(_04627_),
    .X(_05572_));
 sky130_fd_sc_hd__nor2_1 _09710_ (.A(_05568_),
    .B(net258),
    .Y(_05573_));
 sky130_fd_sc_hd__a32o_1 _09711_ (.A1(_04619_),
    .A2(_05571_),
    .A3(_05572_),
    .B1(_05573_),
    .B2(_04613_),
    .X(_00149_));
 sky130_fd_sc_hd__clkbuf_4 _09712_ (.A(_04625_),
    .X(_05574_));
 sky130_fd_sc_hd__clkbuf_4 _09713_ (.A(_05574_),
    .X(_05575_));
 sky130_fd_sc_hd__clkbuf_4 _09714_ (.A(_04626_),
    .X(_05576_));
 sky130_fd_sc_hd__nand2_1 _09715_ (.A(_04613_),
    .B(_05576_),
    .Y(_05577_));
 sky130_fd_sc_hd__a21o_1 _09716_ (.A1(_05575_),
    .A2(_05577_),
    .B1(_04629_),
    .X(_05578_));
 sky130_fd_sc_hd__xor2_1 _09717_ (.A(\round[1] ),
    .B(_04613_),
    .X(_05579_));
 sky130_fd_sc_hd__xnor2_1 _09718_ (.A(_05578_),
    .B(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__a21oi_1 _09719_ (.A1(_05198_),
    .A2(net258),
    .B1(_05568_),
    .Y(_05581_));
 sky130_fd_sc_hd__or2_1 _09720_ (.A(\round[1] ),
    .B(net258),
    .X(_05582_));
 sky130_fd_sc_hd__a22o_1 _09721_ (.A1(_04619_),
    .A2(_05580_),
    .B1(_05581_),
    .B2(_05582_),
    .X(_00150_));
 sky130_fd_sc_hd__and2_1 _09722_ (.A(_04617_),
    .B(\mix1.ready_o ),
    .X(_05583_));
 sky130_fd_sc_hd__buf_2 _09723_ (.A(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__buf_4 _09724_ (.A(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_4 _09725_ (.A(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__nor2_1 _09726_ (.A(_04614_),
    .B(_05575_),
    .Y(_05587_));
 sky130_fd_sc_hd__or3_1 _09727_ (.A(\round[1] ),
    .B(_04613_),
    .C(_05574_),
    .X(_05588_));
 sky130_fd_sc_hd__and2_1 _09728_ (.A(\round[2] ),
    .B(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__and3_1 _09729_ (.A(\round[1] ),
    .B(_04613_),
    .C(\round[2] ),
    .X(_05590_));
 sky130_fd_sc_hd__a21oi_1 _09730_ (.A1(\round[1] ),
    .A2(_04613_),
    .B1(\round[2] ),
    .Y(_05591_));
 sky130_fd_sc_hd__o21ai_1 _09731_ (.A1(_05590_),
    .A2(_05591_),
    .B1(_05586_),
    .Y(_05592_));
 sky130_fd_sc_hd__o31a_1 _09732_ (.A1(_05586_),
    .A2(_05587_),
    .A3(_05589_),
    .B1(_05592_),
    .X(_05593_));
 sky130_fd_sc_hd__a32o_1 _09733_ (.A1(_05568_),
    .A2(_04623_),
    .A3(_05593_),
    .B1(_05573_),
    .B2(\round[2] ),
    .X(_00151_));
 sky130_fd_sc_hd__o21ai_1 _09734_ (.A1(\round[3] ),
    .A2(_05590_),
    .B1(_05586_),
    .Y(_05594_));
 sky130_fd_sc_hd__a21oi_1 _09735_ (.A1(\round[3] ),
    .A2(_05590_),
    .B1(_05594_),
    .Y(_05595_));
 sky130_fd_sc_hd__or3b_1 _09736_ (.A(_05588_),
    .B(\round[2] ),
    .C_N(\round[3] ),
    .X(_05596_));
 sky130_fd_sc_hd__o211a_1 _09737_ (.A1(\round[3] ),
    .A2(_05587_),
    .B1(_05596_),
    .C1(_05576_),
    .X(_05597_));
 sky130_fd_sc_hd__buf_4 _09738_ (.A(_05202_),
    .X(_05598_));
 sky130_fd_sc_hd__o21ai_1 _09739_ (.A1(_05598_),
    .A2(addroundkey_ready_o),
    .B1(_04618_),
    .Y(_05599_));
 sky130_fd_sc_hd__o211a_1 _09740_ (.A1(_05595_),
    .A2(_05597_),
    .B1(_05599_),
    .C1(_05568_),
    .X(_05600_));
 sky130_fd_sc_hd__o32a_1 _09741_ (.A1(\round[3] ),
    .A2(_05568_),
    .A3(net258),
    .B1(_05581_),
    .B2(_05600_),
    .X(_00152_));
 sky130_fd_sc_hd__nor2_1 _09742_ (.A(_04624_),
    .B(_04615_),
    .Y(_05601_));
 sky130_fd_sc_hd__buf_4 _09743_ (.A(_05601_),
    .X(_05602_));
 sky130_fd_sc_hd__buf_4 _09744_ (.A(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__clkbuf_4 _09745_ (.A(_05603_),
    .X(_05604_));
 sky130_fd_sc_hd__mux2_1 _09746_ (.A0(net1),
    .A1(\mix1.data_o[0] ),
    .S(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__clkbuf_4 _09747_ (.A(_04900_),
    .X(_05606_));
 sky130_fd_sc_hd__clkbuf_4 _09748_ (.A(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__buf_4 _09749_ (.A(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__buf_4 _09750_ (.A(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__clkbuf_4 _09751_ (.A(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__mux2_1 _09752_ (.A0(\sub1.data_o[0] ),
    .A1(_05605_),
    .S(_05610_),
    .X(_05611_));
 sky130_fd_sc_hd__or2_1 _09753_ (.A(_04618_),
    .B(_04629_),
    .X(_05612_));
 sky130_fd_sc_hd__buf_4 _09754_ (.A(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__o21ai_4 _09755_ (.A1(_04627_),
    .A2(_05613_),
    .B1(_04609_),
    .Y(_05614_));
 sky130_fd_sc_hd__clkbuf_4 _09756_ (.A(_05614_),
    .X(_05615_));
 sky130_fd_sc_hd__nor2_2 _09757_ (.A(_04618_),
    .B(_04629_),
    .Y(_05616_));
 sky130_fd_sc_hd__buf_4 _09758_ (.A(_05616_),
    .X(_05617_));
 sky130_fd_sc_hd__clkbuf_4 _09759_ (.A(_05617_),
    .X(_05618_));
 sky130_fd_sc_hd__nand2_4 _09760_ (.A(_04625_),
    .B(_05616_),
    .Y(_05619_));
 sky130_fd_sc_hd__clkbuf_4 _09761_ (.A(_05619_),
    .X(_05620_));
 sky130_fd_sc_hd__clkbuf_4 _09762_ (.A(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__a32o_1 _09763_ (.A1(\mix1.data_o[0] ),
    .A2(_05586_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[0] ),
    .X(_05622_));
 sky130_fd_sc_hd__buf_6 _09764_ (.A(_04609_),
    .X(_05623_));
 sky130_fd_sc_hd__a22o_2 _09765_ (.A1(_05611_),
    .A2(_05615_),
    .B1(_05622_),
    .B2(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__buf_4 _09766_ (.A(_04639_),
    .X(_05625_));
 sky130_fd_sc_hd__mux2_1 _09767_ (.A0(net130),
    .A1(\ks1.key_reg[0] ),
    .S(_05625_),
    .X(_05626_));
 sky130_fd_sc_hd__xor2_1 _09768_ (.A(_05624_),
    .B(_05626_),
    .X(_05627_));
 sky130_fd_sc_hd__mux2_1 _09769_ (.A0(\addroundkey_data_o[0] ),
    .A1(_05627_),
    .S(next_addroundkey_ready_o),
    .X(_05628_));
 sky130_fd_sc_hd__clkbuf_1 _09770_ (.A(_05628_),
    .X(_00153_));
 sky130_fd_sc_hd__clkbuf_4 _09771_ (.A(_05615_),
    .X(_05629_));
 sky130_fd_sc_hd__mux2_1 _09772_ (.A0(net40),
    .A1(\mix1.data_o[1] ),
    .S(_05604_),
    .X(_05630_));
 sky130_fd_sc_hd__mux2_1 _09773_ (.A0(\sub1.data_o[1] ),
    .A1(_05630_),
    .S(_05610_),
    .X(_05631_));
 sky130_fd_sc_hd__a32o_1 _09774_ (.A1(\mix1.data_o[1] ),
    .A2(_05586_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[1] ),
    .X(_05632_));
 sky130_fd_sc_hd__clkbuf_4 _09775_ (.A(_05567_),
    .X(_05633_));
 sky130_fd_sc_hd__a22o_1 _09776_ (.A1(_05629_),
    .A2(_05631_),
    .B1(_05632_),
    .B2(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__mux2_2 _09777_ (.A0(net169),
    .A1(\ks1.key_reg[1] ),
    .S(_05625_),
    .X(_05635_));
 sky130_fd_sc_hd__xor2_1 _09778_ (.A(_05634_),
    .B(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__mux2_1 _09779_ (.A0(\addroundkey_data_o[1] ),
    .A1(_05636_),
    .S(next_addroundkey_ready_o),
    .X(_05637_));
 sky130_fd_sc_hd__clkbuf_1 _09780_ (.A(_05637_),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _09781_ (.A0(net51),
    .A1(\mix1.data_o[2] ),
    .S(_05604_),
    .X(_05638_));
 sky130_fd_sc_hd__mux2_1 _09782_ (.A0(\sub1.data_o[2] ),
    .A1(_05638_),
    .S(_05610_),
    .X(_05639_));
 sky130_fd_sc_hd__a32o_1 _09783_ (.A1(\mix1.data_o[2] ),
    .A2(_05586_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[2] ),
    .X(_05640_));
 sky130_fd_sc_hd__a22o_1 _09784_ (.A1(_05629_),
    .A2(_05639_),
    .B1(_05640_),
    .B2(_05633_),
    .X(_05641_));
 sky130_fd_sc_hd__mux2_2 _09785_ (.A0(net180),
    .A1(\ks1.key_reg[2] ),
    .S(_05625_),
    .X(_05642_));
 sky130_fd_sc_hd__xor2_1 _09786_ (.A(_05641_),
    .B(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(\addroundkey_data_o[2] ),
    .A1(_05643_),
    .S(next_addroundkey_ready_o),
    .X(_05644_));
 sky130_fd_sc_hd__clkbuf_1 _09788_ (.A(_05644_),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _09789_ (.A0(net62),
    .A1(\mix1.data_o[3] ),
    .S(_05604_),
    .X(_05645_));
 sky130_fd_sc_hd__mux2_1 _09790_ (.A0(\sub1.data_o[3] ),
    .A1(_05645_),
    .S(_05610_),
    .X(_05646_));
 sky130_fd_sc_hd__a32o_1 _09791_ (.A1(\mix1.data_o[3] ),
    .A2(_05586_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[3] ),
    .X(_05647_));
 sky130_fd_sc_hd__a22o_1 _09792_ (.A1(_05629_),
    .A2(_05646_),
    .B1(_05647_),
    .B2(_05633_),
    .X(_05648_));
 sky130_fd_sc_hd__mux2_1 _09793_ (.A0(net191),
    .A1(\ks1.key_reg[3] ),
    .S(_05625_),
    .X(_05649_));
 sky130_fd_sc_hd__xor2_1 _09794_ (.A(_05648_),
    .B(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__mux2_1 _09795_ (.A0(\addroundkey_data_o[3] ),
    .A1(_05650_),
    .S(next_addroundkey_ready_o),
    .X(_05651_));
 sky130_fd_sc_hd__clkbuf_1 _09796_ (.A(_05651_),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _09797_ (.A0(net73),
    .A1(\mix1.data_o[4] ),
    .S(_05604_),
    .X(_05652_));
 sky130_fd_sc_hd__mux2_1 _09798_ (.A0(\sub1.data_o[4] ),
    .A1(_05652_),
    .S(_05610_),
    .X(_05653_));
 sky130_fd_sc_hd__a32o_1 _09799_ (.A1(\mix1.data_o[4] ),
    .A2(_05586_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[4] ),
    .X(_05654_));
 sky130_fd_sc_hd__a22o_1 _09800_ (.A1(_05629_),
    .A2(_05653_),
    .B1(_05654_),
    .B2(_05633_),
    .X(_05655_));
 sky130_fd_sc_hd__mux2_1 _09801_ (.A0(net202),
    .A1(\ks1.key_reg[4] ),
    .S(_05625_),
    .X(_05656_));
 sky130_fd_sc_hd__xor2_1 _09802_ (.A(_05655_),
    .B(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__mux2_1 _09803_ (.A0(\addroundkey_data_o[4] ),
    .A1(_05657_),
    .S(next_addroundkey_ready_o),
    .X(_05658_));
 sky130_fd_sc_hd__clkbuf_1 _09804_ (.A(_05658_),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _09805_ (.A0(net84),
    .A1(\mix1.data_o[5] ),
    .S(_05604_),
    .X(_05659_));
 sky130_fd_sc_hd__mux2_1 _09806_ (.A0(\sub1.data_o[5] ),
    .A1(_05659_),
    .S(_05610_),
    .X(_05660_));
 sky130_fd_sc_hd__a32o_1 _09807_ (.A1(\mix1.data_o[5] ),
    .A2(_05586_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[5] ),
    .X(_05661_));
 sky130_fd_sc_hd__a22o_1 _09808_ (.A1(_05629_),
    .A2(_05660_),
    .B1(_05661_),
    .B2(_05633_),
    .X(_05662_));
 sky130_fd_sc_hd__mux2_2 _09809_ (.A0(net213),
    .A1(\ks1.key_reg[5] ),
    .S(_05625_),
    .X(_05663_));
 sky130_fd_sc_hd__xor2_1 _09810_ (.A(_05662_),
    .B(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__mux2_1 _09811_ (.A0(\addroundkey_data_o[5] ),
    .A1(_05664_),
    .S(next_addroundkey_ready_o),
    .X(_05665_));
 sky130_fd_sc_hd__clkbuf_1 _09812_ (.A(_05665_),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _09813_ (.A0(net95),
    .A1(\mix1.data_o[6] ),
    .S(_05604_),
    .X(_05666_));
 sky130_fd_sc_hd__mux2_1 _09814_ (.A0(\sub1.data_o[6] ),
    .A1(_05666_),
    .S(_05610_),
    .X(_05667_));
 sky130_fd_sc_hd__a32o_1 _09815_ (.A1(\mix1.data_o[6] ),
    .A2(_05586_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[6] ),
    .X(_05668_));
 sky130_fd_sc_hd__a22o_1 _09816_ (.A1(_05629_),
    .A2(_05667_),
    .B1(_05668_),
    .B2(_05633_),
    .X(_05669_));
 sky130_fd_sc_hd__mux2_1 _09817_ (.A0(net224),
    .A1(\ks1.key_reg[6] ),
    .S(_05625_),
    .X(_05670_));
 sky130_fd_sc_hd__xor2_1 _09818_ (.A(_05669_),
    .B(_05670_),
    .X(_05671_));
 sky130_fd_sc_hd__mux2_1 _09819_ (.A0(\addroundkey_data_o[6] ),
    .A1(_05671_),
    .S(next_addroundkey_ready_o),
    .X(_05672_));
 sky130_fd_sc_hd__clkbuf_1 _09820_ (.A(_05672_),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _09821_ (.A0(net106),
    .A1(\mix1.data_o[7] ),
    .S(_05604_),
    .X(_05673_));
 sky130_fd_sc_hd__mux2_1 _09822_ (.A0(\sub1.data_o[7] ),
    .A1(_05673_),
    .S(_05610_),
    .X(_05674_));
 sky130_fd_sc_hd__clkbuf_4 _09823_ (.A(_05584_),
    .X(_05675_));
 sky130_fd_sc_hd__buf_4 _09824_ (.A(_05675_),
    .X(_05676_));
 sky130_fd_sc_hd__clkbuf_4 _09825_ (.A(_05676_),
    .X(_05677_));
 sky130_fd_sc_hd__a32o_1 _09826_ (.A1(\mix1.data_o[7] ),
    .A2(_05677_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[7] ),
    .X(_05678_));
 sky130_fd_sc_hd__a22o_1 _09827_ (.A1(_05629_),
    .A2(_05674_),
    .B1(_05678_),
    .B2(_05633_),
    .X(_05679_));
 sky130_fd_sc_hd__mux2_1 _09828_ (.A0(net235),
    .A1(\ks1.key_reg[7] ),
    .S(_05625_),
    .X(_05680_));
 sky130_fd_sc_hd__xor2_1 _09829_ (.A(_05679_),
    .B(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__mux2_1 _09830_ (.A0(\addroundkey_data_o[7] ),
    .A1(_05681_),
    .S(next_addroundkey_ready_o),
    .X(_05682_));
 sky130_fd_sc_hd__clkbuf_1 _09831_ (.A(_05682_),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _09832_ (.A0(net117),
    .A1(\mix1.data_o[8] ),
    .S(_05604_),
    .X(_05683_));
 sky130_fd_sc_hd__mux2_1 _09833_ (.A0(\sub1.data_o[8] ),
    .A1(_05683_),
    .S(_05610_),
    .X(_05684_));
 sky130_fd_sc_hd__a32o_1 _09834_ (.A1(\mix1.data_o[8] ),
    .A2(_05677_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[8] ),
    .X(_05685_));
 sky130_fd_sc_hd__a22o_1 _09835_ (.A1(_05629_),
    .A2(_05684_),
    .B1(_05685_),
    .B2(_05633_),
    .X(_05686_));
 sky130_fd_sc_hd__mux2_1 _09836_ (.A0(net246),
    .A1(\ks1.key_reg[8] ),
    .S(_05625_),
    .X(_05687_));
 sky130_fd_sc_hd__xor2_1 _09837_ (.A(_05686_),
    .B(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__mux2_1 _09838_ (.A0(\addroundkey_data_o[8] ),
    .A1(_05688_),
    .S(next_addroundkey_ready_o),
    .X(_05689_));
 sky130_fd_sc_hd__clkbuf_1 _09839_ (.A(_05689_),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _09840_ (.A0(net128),
    .A1(\mix1.data_o[9] ),
    .S(_05604_),
    .X(_05690_));
 sky130_fd_sc_hd__mux2_1 _09841_ (.A0(\sub1.data_o[9] ),
    .A1(_05690_),
    .S(_05610_),
    .X(_05691_));
 sky130_fd_sc_hd__a32o_1 _09842_ (.A1(\mix1.data_o[9] ),
    .A2(_05677_),
    .A3(_05618_),
    .B1(_05621_),
    .B2(\sub1.data_o[9] ),
    .X(_05692_));
 sky130_fd_sc_hd__a22o_1 _09843_ (.A1(_05629_),
    .A2(_05691_),
    .B1(_05692_),
    .B2(_05633_),
    .X(_05693_));
 sky130_fd_sc_hd__mux2_2 _09844_ (.A0(net257),
    .A1(\ks1.key_reg[9] ),
    .S(_05625_),
    .X(_05694_));
 sky130_fd_sc_hd__xor2_1 _09845_ (.A(_05693_),
    .B(_05694_),
    .X(_05695_));
 sky130_fd_sc_hd__buf_4 _09846_ (.A(_04640_),
    .X(_05696_));
 sky130_fd_sc_hd__buf_4 _09847_ (.A(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__mux2_1 _09848_ (.A0(\addroundkey_data_o[9] ),
    .A1(_05695_),
    .S(_05697_),
    .X(_05698_));
 sky130_fd_sc_hd__clkbuf_1 _09849_ (.A(_05698_),
    .X(_00162_));
 sky130_fd_sc_hd__buf_4 _09850_ (.A(_05603_),
    .X(_05699_));
 sky130_fd_sc_hd__mux2_1 _09851_ (.A0(net12),
    .A1(\mix1.data_o[10] ),
    .S(_05699_),
    .X(_05700_));
 sky130_fd_sc_hd__buf_4 _09852_ (.A(_05609_),
    .X(_05701_));
 sky130_fd_sc_hd__mux2_1 _09853_ (.A0(\sub1.data_o[10] ),
    .A1(_05700_),
    .S(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__clkbuf_4 _09854_ (.A(_05617_),
    .X(_05703_));
 sky130_fd_sc_hd__clkbuf_4 _09855_ (.A(_05620_),
    .X(_05704_));
 sky130_fd_sc_hd__a32o_1 _09856_ (.A1(\mix1.data_o[10] ),
    .A2(_05677_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[10] ),
    .X(_05705_));
 sky130_fd_sc_hd__a22o_1 _09857_ (.A1(_05629_),
    .A2(_05702_),
    .B1(_05705_),
    .B2(_05633_),
    .X(_05706_));
 sky130_fd_sc_hd__clkbuf_4 _09858_ (.A(_04638_),
    .X(_05707_));
 sky130_fd_sc_hd__buf_4 _09859_ (.A(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__mux2_1 _09860_ (.A0(net141),
    .A1(\ks1.key_reg[10] ),
    .S(_05708_),
    .X(_05709_));
 sky130_fd_sc_hd__xor2_1 _09861_ (.A(_05706_),
    .B(_05709_),
    .X(_05710_));
 sky130_fd_sc_hd__mux2_1 _09862_ (.A0(\addroundkey_data_o[10] ),
    .A1(_05710_),
    .S(_05697_),
    .X(_05711_));
 sky130_fd_sc_hd__clkbuf_1 _09863_ (.A(_05711_),
    .X(_00163_));
 sky130_fd_sc_hd__clkbuf_4 _09864_ (.A(_05615_),
    .X(_05712_));
 sky130_fd_sc_hd__mux2_1 _09865_ (.A0(net23),
    .A1(\mix1.data_o[11] ),
    .S(_05699_),
    .X(_05713_));
 sky130_fd_sc_hd__mux2_1 _09866_ (.A0(\sub1.data_o[11] ),
    .A1(_05713_),
    .S(_05701_),
    .X(_05714_));
 sky130_fd_sc_hd__a32o_1 _09867_ (.A1(\mix1.data_o[11] ),
    .A2(_05677_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[11] ),
    .X(_05715_));
 sky130_fd_sc_hd__clkbuf_4 _09868_ (.A(_05567_),
    .X(_05716_));
 sky130_fd_sc_hd__a22o_1 _09869_ (.A1(_05712_),
    .A2(_05714_),
    .B1(_05715_),
    .B2(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__mux2_1 _09870_ (.A0(net152),
    .A1(\ks1.key_reg[11] ),
    .S(_05708_),
    .X(_05718_));
 sky130_fd_sc_hd__xor2_1 _09871_ (.A(_05717_),
    .B(_05718_),
    .X(_05719_));
 sky130_fd_sc_hd__mux2_1 _09872_ (.A0(\addroundkey_data_o[11] ),
    .A1(_05719_),
    .S(_05697_),
    .X(_05720_));
 sky130_fd_sc_hd__clkbuf_1 _09873_ (.A(_05720_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _09874_ (.A0(net32),
    .A1(\mix1.data_o[12] ),
    .S(_05699_),
    .X(_05721_));
 sky130_fd_sc_hd__mux2_1 _09875_ (.A0(\sub1.data_o[12] ),
    .A1(_05721_),
    .S(_05701_),
    .X(_05722_));
 sky130_fd_sc_hd__a32o_1 _09876_ (.A1(\mix1.data_o[12] ),
    .A2(_05677_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[12] ),
    .X(_05723_));
 sky130_fd_sc_hd__a22o_1 _09877_ (.A1(_05712_),
    .A2(_05722_),
    .B1(_05723_),
    .B2(_05716_),
    .X(_05724_));
 sky130_fd_sc_hd__mux2_1 _09878_ (.A0(net161),
    .A1(\ks1.key_reg[12] ),
    .S(_05708_),
    .X(_05725_));
 sky130_fd_sc_hd__xor2_1 _09879_ (.A(_05724_),
    .B(_05725_),
    .X(_05726_));
 sky130_fd_sc_hd__mux2_1 _09880_ (.A0(\addroundkey_data_o[12] ),
    .A1(_05726_),
    .S(_05697_),
    .X(_05727_));
 sky130_fd_sc_hd__clkbuf_1 _09881_ (.A(_05727_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(net33),
    .A1(\mix1.data_o[13] ),
    .S(_05699_),
    .X(_05728_));
 sky130_fd_sc_hd__mux2_1 _09883_ (.A0(\sub1.data_o[13] ),
    .A1(_05728_),
    .S(_05701_),
    .X(_05729_));
 sky130_fd_sc_hd__a32o_1 _09884_ (.A1(\mix1.data_o[13] ),
    .A2(_05677_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[13] ),
    .X(_05730_));
 sky130_fd_sc_hd__a22o_1 _09885_ (.A1(_05712_),
    .A2(_05729_),
    .B1(_05730_),
    .B2(_05716_),
    .X(_05731_));
 sky130_fd_sc_hd__mux2_2 _09886_ (.A0(net162),
    .A1(\ks1.key_reg[13] ),
    .S(_05708_),
    .X(_05732_));
 sky130_fd_sc_hd__xor2_1 _09887_ (.A(_05731_),
    .B(_05732_),
    .X(_05733_));
 sky130_fd_sc_hd__mux2_1 _09888_ (.A0(\addroundkey_data_o[13] ),
    .A1(_05733_),
    .S(_05697_),
    .X(_05734_));
 sky130_fd_sc_hd__clkbuf_1 _09889_ (.A(_05734_),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _09890_ (.A0(net34),
    .A1(\mix1.data_o[14] ),
    .S(_05699_),
    .X(_05735_));
 sky130_fd_sc_hd__mux2_1 _09891_ (.A0(\sub1.data_o[14] ),
    .A1(_05735_),
    .S(_05701_),
    .X(_05736_));
 sky130_fd_sc_hd__a32o_1 _09892_ (.A1(\mix1.data_o[14] ),
    .A2(_05677_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[14] ),
    .X(_05737_));
 sky130_fd_sc_hd__a22o_1 _09893_ (.A1(_05712_),
    .A2(_05736_),
    .B1(_05737_),
    .B2(_05716_),
    .X(_05738_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(net163),
    .A1(\ks1.key_reg[14] ),
    .S(_05708_),
    .X(_05739_));
 sky130_fd_sc_hd__xor2_1 _09895_ (.A(_05738_),
    .B(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__mux2_1 _09896_ (.A0(\addroundkey_data_o[14] ),
    .A1(_05740_),
    .S(_05697_),
    .X(_05741_));
 sky130_fd_sc_hd__clkbuf_1 _09897_ (.A(_05741_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _09898_ (.A0(net35),
    .A1(\mix1.data_o[15] ),
    .S(_05699_),
    .X(_05742_));
 sky130_fd_sc_hd__mux2_1 _09899_ (.A0(\sub1.data_o[15] ),
    .A1(_05742_),
    .S(_05701_),
    .X(_05743_));
 sky130_fd_sc_hd__a32o_1 _09900_ (.A1(\mix1.data_o[15] ),
    .A2(_05677_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[15] ),
    .X(_05744_));
 sky130_fd_sc_hd__a22o_1 _09901_ (.A1(_05712_),
    .A2(_05743_),
    .B1(_05744_),
    .B2(_05716_),
    .X(_05745_));
 sky130_fd_sc_hd__mux2_1 _09902_ (.A0(net164),
    .A1(\ks1.key_reg[15] ),
    .S(_05708_),
    .X(_05746_));
 sky130_fd_sc_hd__xor2_1 _09903_ (.A(_05745_),
    .B(_05746_),
    .X(_05747_));
 sky130_fd_sc_hd__mux2_1 _09904_ (.A0(\addroundkey_data_o[15] ),
    .A1(_05747_),
    .S(_05697_),
    .X(_05748_));
 sky130_fd_sc_hd__clkbuf_1 _09905_ (.A(_05748_),
    .X(_00168_));
 sky130_fd_sc_hd__buf_4 _09906_ (.A(_05601_),
    .X(_05749_));
 sky130_fd_sc_hd__mux2_1 _09907_ (.A0(net36),
    .A1(\mix1.data_o[16] ),
    .S(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__buf_4 _09908_ (.A(_05607_),
    .X(_05751_));
 sky130_fd_sc_hd__mux2_1 _09909_ (.A0(\sub1.data_o[16] ),
    .A1(_05750_),
    .S(_05751_),
    .X(_05752_));
 sky130_fd_sc_hd__clkbuf_4 _09910_ (.A(_05613_),
    .X(_05753_));
 sky130_fd_sc_hd__buf_2 _09911_ (.A(\sub1.ready_o ),
    .X(_05754_));
 sky130_fd_sc_hd__a31o_1 _09912_ (.A1(_05201_),
    .A2(_05754_),
    .A3(\sub1.data_o[16] ),
    .B1(_05585_),
    .X(_05755_));
 sky130_fd_sc_hd__a21o_1 _09913_ (.A1(_05575_),
    .A2(_05752_),
    .B1(_05755_),
    .X(_05756_));
 sky130_fd_sc_hd__buf_8 _09914_ (.A(_05616_),
    .X(_05757_));
 sky130_fd_sc_hd__buf_4 _09915_ (.A(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__o21a_1 _09916_ (.A1(\mix1.data_o[16] ),
    .A2(_05576_),
    .B1(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__a221o_1 _09917_ (.A1(\sub1.data_o[16] ),
    .A2(_05753_),
    .B1(_05756_),
    .B2(_05759_),
    .C1(_04611_),
    .X(_05760_));
 sky130_fd_sc_hd__o21ai_1 _09918_ (.A1(_05568_),
    .A2(_05752_),
    .B1(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__buf_4 _09919_ (.A(_05707_),
    .X(_05762_));
 sky130_fd_sc_hd__mux2_4 _09920_ (.A0(net165),
    .A1(\ks1.key_reg[16] ),
    .S(_05762_),
    .X(_05763_));
 sky130_fd_sc_hd__xnor2_1 _09921_ (.A(_05761_),
    .B(_05763_),
    .Y(_05764_));
 sky130_fd_sc_hd__mux2_1 _09922_ (.A0(\addroundkey_data_o[16] ),
    .A1(_05764_),
    .S(_05697_),
    .X(_05765_));
 sky130_fd_sc_hd__clkbuf_1 _09923_ (.A(_05765_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _09924_ (.A0(net37),
    .A1(\mix1.data_o[17] ),
    .S(_05749_),
    .X(_05766_));
 sky130_fd_sc_hd__mux2_1 _09925_ (.A0(\sub1.data_o[17] ),
    .A1(_05766_),
    .S(_05751_),
    .X(_05767_));
 sky130_fd_sc_hd__a31o_1 _09926_ (.A1(_05201_),
    .A2(_05754_),
    .A3(\sub1.data_o[17] ),
    .B1(_05585_),
    .X(_05768_));
 sky130_fd_sc_hd__a21o_1 _09927_ (.A1(_05575_),
    .A2(_05767_),
    .B1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__o21a_1 _09928_ (.A1(\mix1.data_o[17] ),
    .A2(_05576_),
    .B1(_05758_),
    .X(_05770_));
 sky130_fd_sc_hd__a221o_1 _09929_ (.A1(\sub1.data_o[17] ),
    .A2(_05753_),
    .B1(_05769_),
    .B2(_05770_),
    .C1(_04611_),
    .X(_05771_));
 sky130_fd_sc_hd__o21ai_1 _09930_ (.A1(_05568_),
    .A2(_05767_),
    .B1(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__mux2_2 _09931_ (.A0(net166),
    .A1(\ks1.key_reg[17] ),
    .S(_05762_),
    .X(_05773_));
 sky130_fd_sc_hd__xnor2_1 _09932_ (.A(_05772_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__mux2_1 _09933_ (.A0(\addroundkey_data_o[17] ),
    .A1(_05774_),
    .S(_05697_),
    .X(_05775_));
 sky130_fd_sc_hd__clkbuf_1 _09934_ (.A(_05775_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _09935_ (.A0(net38),
    .A1(\mix1.data_o[18] ),
    .S(_05749_),
    .X(_05776_));
 sky130_fd_sc_hd__mux2_1 _09936_ (.A0(\sub1.data_o[18] ),
    .A1(_05776_),
    .S(_05751_),
    .X(_05777_));
 sky130_fd_sc_hd__a31o_1 _09937_ (.A1(_05201_),
    .A2(_05754_),
    .A3(\sub1.data_o[18] ),
    .B1(_05585_),
    .X(_05778_));
 sky130_fd_sc_hd__a21o_1 _09938_ (.A1(_05575_),
    .A2(_05777_),
    .B1(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__o21a_1 _09939_ (.A1(\mix1.data_o[18] ),
    .A2(_05576_),
    .B1(_05758_),
    .X(_05780_));
 sky130_fd_sc_hd__a221o_1 _09940_ (.A1(\sub1.data_o[18] ),
    .A2(_05753_),
    .B1(_05779_),
    .B2(_05780_),
    .C1(_04611_),
    .X(_05781_));
 sky130_fd_sc_hd__o21ai_1 _09941_ (.A1(_05568_),
    .A2(_05777_),
    .B1(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__mux2_2 _09942_ (.A0(net167),
    .A1(\ks1.key_reg[18] ),
    .S(_05762_),
    .X(_05783_));
 sky130_fd_sc_hd__xnor2_1 _09943_ (.A(_05782_),
    .B(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__mux2_1 _09944_ (.A0(\addroundkey_data_o[18] ),
    .A1(_05784_),
    .S(_05697_),
    .X(_05785_));
 sky130_fd_sc_hd__clkbuf_1 _09945_ (.A(_05785_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _09946_ (.A0(net39),
    .A1(\mix1.data_o[19] ),
    .S(_05699_),
    .X(_05786_));
 sky130_fd_sc_hd__mux2_1 _09947_ (.A0(\sub1.data_o[19] ),
    .A1(_05786_),
    .S(_05701_),
    .X(_05787_));
 sky130_fd_sc_hd__a32o_1 _09948_ (.A1(\mix1.data_o[19] ),
    .A2(_05677_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[19] ),
    .X(_05788_));
 sky130_fd_sc_hd__a22o_1 _09949_ (.A1(_05712_),
    .A2(_05787_),
    .B1(_05788_),
    .B2(_05716_),
    .X(_05789_));
 sky130_fd_sc_hd__mux2_1 _09950_ (.A0(net168),
    .A1(\ks1.key_reg[19] ),
    .S(_05708_),
    .X(_05790_));
 sky130_fd_sc_hd__xor2_1 _09951_ (.A(_05789_),
    .B(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__buf_4 _09952_ (.A(_04640_),
    .X(_05792_));
 sky130_fd_sc_hd__buf_4 _09953_ (.A(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__mux2_1 _09954_ (.A0(\addroundkey_data_o[19] ),
    .A1(_05791_),
    .S(_05793_),
    .X(_05794_));
 sky130_fd_sc_hd__clkbuf_1 _09955_ (.A(_05794_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _09956_ (.A0(net41),
    .A1(\mix1.data_o[20] ),
    .S(_05699_),
    .X(_05795_));
 sky130_fd_sc_hd__mux2_1 _09957_ (.A0(\sub1.data_o[20] ),
    .A1(_05795_),
    .S(_05701_),
    .X(_05796_));
 sky130_fd_sc_hd__clkbuf_4 _09958_ (.A(_05676_),
    .X(_05797_));
 sky130_fd_sc_hd__a32o_1 _09959_ (.A1(\mix1.data_o[20] ),
    .A2(_05797_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[20] ),
    .X(_05798_));
 sky130_fd_sc_hd__a22o_1 _09960_ (.A1(_05712_),
    .A2(_05796_),
    .B1(_05798_),
    .B2(_05716_),
    .X(_05799_));
 sky130_fd_sc_hd__mux2_1 _09961_ (.A0(net170),
    .A1(\ks1.key_reg[20] ),
    .S(_05708_),
    .X(_05800_));
 sky130_fd_sc_hd__xor2_1 _09962_ (.A(_05799_),
    .B(_05800_),
    .X(_05801_));
 sky130_fd_sc_hd__mux2_1 _09963_ (.A0(\addroundkey_data_o[20] ),
    .A1(_05801_),
    .S(_05793_),
    .X(_05802_));
 sky130_fd_sc_hd__clkbuf_1 _09964_ (.A(_05802_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _09965_ (.A0(net42),
    .A1(\mix1.data_o[21] ),
    .S(_05699_),
    .X(_05803_));
 sky130_fd_sc_hd__mux2_1 _09966_ (.A0(\sub1.data_o[21] ),
    .A1(_05803_),
    .S(_05701_),
    .X(_05804_));
 sky130_fd_sc_hd__a32o_1 _09967_ (.A1(\mix1.data_o[21] ),
    .A2(_05797_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[21] ),
    .X(_05805_));
 sky130_fd_sc_hd__a22o_1 _09968_ (.A1(_05712_),
    .A2(_05804_),
    .B1(_05805_),
    .B2(_05716_),
    .X(_05806_));
 sky130_fd_sc_hd__mux2_2 _09969_ (.A0(net171),
    .A1(\ks1.key_reg[21] ),
    .S(_05708_),
    .X(_05807_));
 sky130_fd_sc_hd__xor2_1 _09970_ (.A(_05806_),
    .B(_05807_),
    .X(_05808_));
 sky130_fd_sc_hd__mux2_1 _09971_ (.A0(\addroundkey_data_o[21] ),
    .A1(_05808_),
    .S(_05793_),
    .X(_05809_));
 sky130_fd_sc_hd__clkbuf_1 _09972_ (.A(_05809_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _09973_ (.A0(net43),
    .A1(\mix1.data_o[22] ),
    .S(_05699_),
    .X(_05810_));
 sky130_fd_sc_hd__mux2_1 _09974_ (.A0(\sub1.data_o[22] ),
    .A1(_05810_),
    .S(_05701_),
    .X(_05811_));
 sky130_fd_sc_hd__a32o_1 _09975_ (.A1(\mix1.data_o[22] ),
    .A2(_05797_),
    .A3(_05703_),
    .B1(_05704_),
    .B2(\sub1.data_o[22] ),
    .X(_05812_));
 sky130_fd_sc_hd__a22o_1 _09976_ (.A1(_05712_),
    .A2(_05811_),
    .B1(_05812_),
    .B2(_05716_),
    .X(_05813_));
 sky130_fd_sc_hd__mux2_4 _09977_ (.A0(net172),
    .A1(\ks1.key_reg[22] ),
    .S(_05708_),
    .X(_05814_));
 sky130_fd_sc_hd__xor2_1 _09978_ (.A(_05813_),
    .B(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__mux2_1 _09979_ (.A0(\addroundkey_data_o[22] ),
    .A1(_05815_),
    .S(_05793_),
    .X(_05816_));
 sky130_fd_sc_hd__clkbuf_1 _09980_ (.A(_05816_),
    .X(_00175_));
 sky130_fd_sc_hd__buf_4 _09981_ (.A(_05603_),
    .X(_05817_));
 sky130_fd_sc_hd__mux2_1 _09982_ (.A0(net44),
    .A1(\mix1.data_o[23] ),
    .S(_05817_),
    .X(_05818_));
 sky130_fd_sc_hd__clkbuf_4 _09983_ (.A(_05609_),
    .X(_05819_));
 sky130_fd_sc_hd__mux2_1 _09984_ (.A0(\sub1.data_o[23] ),
    .A1(_05818_),
    .S(_05819_),
    .X(_05820_));
 sky130_fd_sc_hd__buf_2 _09985_ (.A(_05757_),
    .X(_05821_));
 sky130_fd_sc_hd__buf_2 _09986_ (.A(_05620_),
    .X(_05822_));
 sky130_fd_sc_hd__a32o_1 _09987_ (.A1(\mix1.data_o[23] ),
    .A2(_05797_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[23] ),
    .X(_05823_));
 sky130_fd_sc_hd__a22o_1 _09988_ (.A1(_05712_),
    .A2(_05820_),
    .B1(_05823_),
    .B2(_05716_),
    .X(_05824_));
 sky130_fd_sc_hd__buf_4 _09989_ (.A(_05707_),
    .X(_05825_));
 sky130_fd_sc_hd__mux2_4 _09990_ (.A0(net173),
    .A1(\ks1.key_reg[23] ),
    .S(_05825_),
    .X(_05826_));
 sky130_fd_sc_hd__xor2_1 _09991_ (.A(_05824_),
    .B(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__mux2_1 _09992_ (.A0(\addroundkey_data_o[23] ),
    .A1(_05827_),
    .S(_05793_),
    .X(_05828_));
 sky130_fd_sc_hd__clkbuf_1 _09993_ (.A(_05828_),
    .X(_00176_));
 sky130_fd_sc_hd__clkbuf_4 _09994_ (.A(_05615_),
    .X(_05829_));
 sky130_fd_sc_hd__mux2_1 _09995_ (.A0(net45),
    .A1(\mix1.data_o[24] ),
    .S(_05817_),
    .X(_05830_));
 sky130_fd_sc_hd__mux2_1 _09996_ (.A0(\sub1.data_o[24] ),
    .A1(_05830_),
    .S(_05819_),
    .X(_05831_));
 sky130_fd_sc_hd__a32o_1 _09997_ (.A1(\mix1.data_o[24] ),
    .A2(_05797_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[24] ),
    .X(_05832_));
 sky130_fd_sc_hd__clkbuf_4 _09998_ (.A(_04609_),
    .X(_05833_));
 sky130_fd_sc_hd__a22o_1 _09999_ (.A1(_05829_),
    .A2(_05831_),
    .B1(_05832_),
    .B2(_05833_),
    .X(_05834_));
 sky130_fd_sc_hd__mux2_1 _10000_ (.A0(net174),
    .A1(\ks1.key_reg[24] ),
    .S(_05825_),
    .X(_05835_));
 sky130_fd_sc_hd__xor2_1 _10001_ (.A(_05834_),
    .B(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__mux2_1 _10002_ (.A0(\addroundkey_data_o[24] ),
    .A1(_05836_),
    .S(_05793_),
    .X(_05837_));
 sky130_fd_sc_hd__clkbuf_1 _10003_ (.A(_05837_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _10004_ (.A0(net46),
    .A1(\mix1.data_o[25] ),
    .S(_05817_),
    .X(_05838_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(\sub1.data_o[25] ),
    .A1(_05838_),
    .S(_05819_),
    .X(_05839_));
 sky130_fd_sc_hd__a32o_1 _10006_ (.A1(\mix1.data_o[25] ),
    .A2(_05797_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[25] ),
    .X(_05840_));
 sky130_fd_sc_hd__a22o_1 _10007_ (.A1(_05829_),
    .A2(_05839_),
    .B1(_05840_),
    .B2(_05833_),
    .X(_05841_));
 sky130_fd_sc_hd__mux2_1 _10008_ (.A0(net175),
    .A1(\ks1.key_reg[25] ),
    .S(_05825_),
    .X(_05842_));
 sky130_fd_sc_hd__xor2_1 _10009_ (.A(_05841_),
    .B(_05842_),
    .X(_05843_));
 sky130_fd_sc_hd__mux2_1 _10010_ (.A0(\addroundkey_data_o[25] ),
    .A1(_05843_),
    .S(_05793_),
    .X(_05844_));
 sky130_fd_sc_hd__clkbuf_1 _10011_ (.A(_05844_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _10012_ (.A0(net47),
    .A1(\mix1.data_o[26] ),
    .S(_05817_),
    .X(_05845_));
 sky130_fd_sc_hd__mux2_1 _10013_ (.A0(\sub1.data_o[26] ),
    .A1(_05845_),
    .S(_05819_),
    .X(_05846_));
 sky130_fd_sc_hd__a32o_1 _10014_ (.A1(\mix1.data_o[26] ),
    .A2(_05797_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[26] ),
    .X(_05847_));
 sky130_fd_sc_hd__a22o_1 _10015_ (.A1(_05829_),
    .A2(_05846_),
    .B1(_05847_),
    .B2(_05833_),
    .X(_05848_));
 sky130_fd_sc_hd__mux2_2 _10016_ (.A0(net176),
    .A1(\ks1.key_reg[26] ),
    .S(_05825_),
    .X(_05849_));
 sky130_fd_sc_hd__xor2_1 _10017_ (.A(_05848_),
    .B(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__mux2_1 _10018_ (.A0(\addroundkey_data_o[26] ),
    .A1(_05850_),
    .S(_05793_),
    .X(_05851_));
 sky130_fd_sc_hd__clkbuf_1 _10019_ (.A(_05851_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _10020_ (.A0(net48),
    .A1(\mix1.data_o[27] ),
    .S(_05817_),
    .X(_05852_));
 sky130_fd_sc_hd__mux2_1 _10021_ (.A0(\sub1.data_o[27] ),
    .A1(_05852_),
    .S(_05819_),
    .X(_05853_));
 sky130_fd_sc_hd__a32o_1 _10022_ (.A1(\mix1.data_o[27] ),
    .A2(_05797_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[27] ),
    .X(_05854_));
 sky130_fd_sc_hd__a22o_1 _10023_ (.A1(_05829_),
    .A2(_05853_),
    .B1(_05854_),
    .B2(_05833_),
    .X(_05855_));
 sky130_fd_sc_hd__mux2_1 _10024_ (.A0(net177),
    .A1(\ks1.key_reg[27] ),
    .S(_05825_),
    .X(_05856_));
 sky130_fd_sc_hd__xor2_1 _10025_ (.A(_05855_),
    .B(_05856_),
    .X(_05857_));
 sky130_fd_sc_hd__mux2_1 _10026_ (.A0(\addroundkey_data_o[27] ),
    .A1(_05857_),
    .S(_05793_),
    .X(_05858_));
 sky130_fd_sc_hd__clkbuf_1 _10027_ (.A(_05858_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _10028_ (.A0(net49),
    .A1(\mix1.data_o[28] ),
    .S(_05817_),
    .X(_05859_));
 sky130_fd_sc_hd__mux2_1 _10029_ (.A0(\sub1.data_o[28] ),
    .A1(_05859_),
    .S(_05819_),
    .X(_05860_));
 sky130_fd_sc_hd__a32o_1 _10030_ (.A1(\mix1.data_o[28] ),
    .A2(_05797_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[28] ),
    .X(_05861_));
 sky130_fd_sc_hd__a22o_1 _10031_ (.A1(_05829_),
    .A2(_05860_),
    .B1(_05861_),
    .B2(_05833_),
    .X(_05862_));
 sky130_fd_sc_hd__mux2_2 _10032_ (.A0(net178),
    .A1(\ks1.key_reg[28] ),
    .S(_05825_),
    .X(_05863_));
 sky130_fd_sc_hd__xor2_1 _10033_ (.A(_05862_),
    .B(_05863_),
    .X(_05864_));
 sky130_fd_sc_hd__mux2_1 _10034_ (.A0(\addroundkey_data_o[28] ),
    .A1(_05864_),
    .S(_05793_),
    .X(_05865_));
 sky130_fd_sc_hd__clkbuf_1 _10035_ (.A(_05865_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _10036_ (.A0(net50),
    .A1(\mix1.data_o[29] ),
    .S(_05817_),
    .X(_05866_));
 sky130_fd_sc_hd__mux2_1 _10037_ (.A0(\sub1.data_o[29] ),
    .A1(_05866_),
    .S(_05819_),
    .X(_05867_));
 sky130_fd_sc_hd__a32o_1 _10038_ (.A1(\mix1.data_o[29] ),
    .A2(_05797_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[29] ),
    .X(_05868_));
 sky130_fd_sc_hd__a22o_1 _10039_ (.A1(_05829_),
    .A2(_05867_),
    .B1(_05868_),
    .B2(_05833_),
    .X(_05869_));
 sky130_fd_sc_hd__mux2_2 _10040_ (.A0(net179),
    .A1(\ks1.key_reg[29] ),
    .S(_05825_),
    .X(_05870_));
 sky130_fd_sc_hd__xor2_1 _10041_ (.A(_05869_),
    .B(_05870_),
    .X(_05871_));
 sky130_fd_sc_hd__buf_4 _10042_ (.A(_05792_),
    .X(_05872_));
 sky130_fd_sc_hd__mux2_1 _10043_ (.A0(\addroundkey_data_o[29] ),
    .A1(_05871_),
    .S(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__clkbuf_1 _10044_ (.A(_05873_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _10045_ (.A0(net52),
    .A1(\mix1.data_o[30] ),
    .S(_05817_),
    .X(_05874_));
 sky130_fd_sc_hd__mux2_1 _10046_ (.A0(\sub1.data_o[30] ),
    .A1(_05874_),
    .S(_05819_),
    .X(_05875_));
 sky130_fd_sc_hd__clkbuf_4 _10047_ (.A(_05585_),
    .X(_05876_));
 sky130_fd_sc_hd__a32o_1 _10048_ (.A1(\mix1.data_o[30] ),
    .A2(_05876_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[30] ),
    .X(_05877_));
 sky130_fd_sc_hd__a22o_1 _10049_ (.A1(_05829_),
    .A2(_05875_),
    .B1(_05877_),
    .B2(_05833_),
    .X(_05878_));
 sky130_fd_sc_hd__mux2_2 _10050_ (.A0(net181),
    .A1(\ks1.key_reg[30] ),
    .S(_05825_),
    .X(_05879_));
 sky130_fd_sc_hd__xor2_1 _10051_ (.A(_05878_),
    .B(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__mux2_1 _10052_ (.A0(\addroundkey_data_o[30] ),
    .A1(_05880_),
    .S(_05872_),
    .X(_05881_));
 sky130_fd_sc_hd__clkbuf_1 _10053_ (.A(_05881_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _10054_ (.A0(net53),
    .A1(\mix1.data_o[31] ),
    .S(_05817_),
    .X(_05882_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(\sub1.data_o[31] ),
    .A1(_05882_),
    .S(_05819_),
    .X(_05883_));
 sky130_fd_sc_hd__a32o_1 _10056_ (.A1(\mix1.data_o[31] ),
    .A2(_05876_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[31] ),
    .X(_05884_));
 sky130_fd_sc_hd__a22o_1 _10057_ (.A1(_05829_),
    .A2(_05883_),
    .B1(_05884_),
    .B2(_05833_),
    .X(_05885_));
 sky130_fd_sc_hd__mux2_2 _10058_ (.A0(net182),
    .A1(\ks1.key_reg[31] ),
    .S(_05825_),
    .X(_05886_));
 sky130_fd_sc_hd__xor2_1 _10059_ (.A(_05885_),
    .B(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__mux2_1 _10060_ (.A0(\addroundkey_data_o[31] ),
    .A1(_05887_),
    .S(_05872_),
    .X(_05888_));
 sky130_fd_sc_hd__clkbuf_1 _10061_ (.A(_05888_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _10062_ (.A0(net54),
    .A1(\mix1.data_o[32] ),
    .S(_05749_),
    .X(_05889_));
 sky130_fd_sc_hd__mux2_1 _10063_ (.A0(\sub1.data_o[32] ),
    .A1(_05889_),
    .S(_05751_),
    .X(_05890_));
 sky130_fd_sc_hd__a31o_1 _10064_ (.A1(_05201_),
    .A2(_05754_),
    .A3(\sub1.data_o[32] ),
    .B1(_05585_),
    .X(_05891_));
 sky130_fd_sc_hd__a21o_1 _10065_ (.A1(_05575_),
    .A2(_05890_),
    .B1(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__o21a_1 _10066_ (.A1(\mix1.data_o[32] ),
    .A2(_05576_),
    .B1(_05758_),
    .X(_05893_));
 sky130_fd_sc_hd__a221o_1 _10067_ (.A1(\sub1.data_o[32] ),
    .A2(_05753_),
    .B1(_05892_),
    .B2(_05893_),
    .C1(_04611_),
    .X(_05894_));
 sky130_fd_sc_hd__o21ai_4 _10068_ (.A1(_05568_),
    .A2(_05890_),
    .B1(_05894_),
    .Y(_05895_));
 sky130_fd_sc_hd__mux2_2 _10069_ (.A0(net183),
    .A1(\ks1.key_reg[32] ),
    .S(_05762_),
    .X(_05896_));
 sky130_fd_sc_hd__xnor2_1 _10070_ (.A(_05895_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__mux2_1 _10071_ (.A0(\addroundkey_data_o[32] ),
    .A1(_05897_),
    .S(_05872_),
    .X(_05898_));
 sky130_fd_sc_hd__clkbuf_1 _10072_ (.A(_05898_),
    .X(_00185_));
 sky130_fd_sc_hd__clkbuf_8 _10073_ (.A(_05567_),
    .X(_05899_));
 sky130_fd_sc_hd__mux2_1 _10074_ (.A0(net55),
    .A1(\mix1.data_o[33] ),
    .S(_05749_),
    .X(_05900_));
 sky130_fd_sc_hd__mux2_1 _10075_ (.A0(\sub1.data_o[33] ),
    .A1(_05900_),
    .S(_05751_),
    .X(_05901_));
 sky130_fd_sc_hd__buf_2 _10076_ (.A(_05584_),
    .X(_05902_));
 sky130_fd_sc_hd__a31o_1 _10077_ (.A1(_05201_),
    .A2(_05754_),
    .A3(\sub1.data_o[33] ),
    .B1(_05902_),
    .X(_05903_));
 sky130_fd_sc_hd__a21o_1 _10078_ (.A1(_05575_),
    .A2(_05901_),
    .B1(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__o21a_1 _10079_ (.A1(\mix1.data_o[33] ),
    .A2(_05576_),
    .B1(_05758_),
    .X(_05905_));
 sky130_fd_sc_hd__a221o_1 _10080_ (.A1(\sub1.data_o[33] ),
    .A2(_05753_),
    .B1(_05904_),
    .B2(_05905_),
    .C1(_04611_),
    .X(_05906_));
 sky130_fd_sc_hd__o21ai_4 _10081_ (.A1(_05899_),
    .A2(_05901_),
    .B1(_05906_),
    .Y(_05907_));
 sky130_fd_sc_hd__mux2_1 _10082_ (.A0(net184),
    .A1(\ks1.key_reg[33] ),
    .S(_05762_),
    .X(_05908_));
 sky130_fd_sc_hd__xnor2_1 _10083_ (.A(_05907_),
    .B(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__mux2_1 _10084_ (.A0(\addroundkey_data_o[33] ),
    .A1(_05909_),
    .S(_05872_),
    .X(_05910_));
 sky130_fd_sc_hd__clkbuf_1 _10085_ (.A(_05910_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _10086_ (.A0(net56),
    .A1(\mix1.data_o[34] ),
    .S(_05749_),
    .X(_05911_));
 sky130_fd_sc_hd__mux2_1 _10087_ (.A0(\sub1.data_o[34] ),
    .A1(_05911_),
    .S(_05751_),
    .X(_05912_));
 sky130_fd_sc_hd__clkbuf_4 _10088_ (.A(_04624_),
    .X(_05913_));
 sky130_fd_sc_hd__a31o_1 _10089_ (.A1(_05913_),
    .A2(_05754_),
    .A3(\sub1.data_o[34] ),
    .B1(_05902_),
    .X(_05914_));
 sky130_fd_sc_hd__a21o_1 _10090_ (.A1(_05575_),
    .A2(_05912_),
    .B1(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__clkbuf_4 _10091_ (.A(_05757_),
    .X(_05916_));
 sky130_fd_sc_hd__o21a_1 _10092_ (.A1(\mix1.data_o[34] ),
    .A2(_05576_),
    .B1(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__a221o_1 _10093_ (.A1(\sub1.data_o[34] ),
    .A2(_05753_),
    .B1(_05915_),
    .B2(_05917_),
    .C1(_04611_),
    .X(_05918_));
 sky130_fd_sc_hd__o21ai_2 _10094_ (.A1(_05899_),
    .A2(_05912_),
    .B1(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__buf_4 _10095_ (.A(_05707_),
    .X(_05920_));
 sky130_fd_sc_hd__mux2_4 _10096_ (.A0(net185),
    .A1(\ks1.key_reg[34] ),
    .S(_05920_),
    .X(_05921_));
 sky130_fd_sc_hd__xnor2_1 _10097_ (.A(_05919_),
    .B(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__mux2_1 _10098_ (.A0(\addroundkey_data_o[34] ),
    .A1(_05922_),
    .S(_05872_),
    .X(_05923_));
 sky130_fd_sc_hd__clkbuf_1 _10099_ (.A(_05923_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _10100_ (.A0(net57),
    .A1(\mix1.data_o[35] ),
    .S(_05749_),
    .X(_05924_));
 sky130_fd_sc_hd__mux2_1 _10101_ (.A0(\sub1.data_o[35] ),
    .A1(_05924_),
    .S(_05751_),
    .X(_05925_));
 sky130_fd_sc_hd__a31o_1 _10102_ (.A1(_05913_),
    .A2(_05754_),
    .A3(\sub1.data_o[35] ),
    .B1(_05902_),
    .X(_05926_));
 sky130_fd_sc_hd__a21o_1 _10103_ (.A1(_05575_),
    .A2(_05925_),
    .B1(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__o21a_1 _10104_ (.A1(\mix1.data_o[35] ),
    .A2(_05576_),
    .B1(_05916_),
    .X(_05928_));
 sky130_fd_sc_hd__a221o_1 _10105_ (.A1(\sub1.data_o[35] ),
    .A2(_05753_),
    .B1(_05927_),
    .B2(_05928_),
    .C1(_04611_),
    .X(_05929_));
 sky130_fd_sc_hd__o21ai_2 _10106_ (.A1(_05899_),
    .A2(_05925_),
    .B1(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__mux2_2 _10107_ (.A0(net186),
    .A1(\ks1.key_reg[35] ),
    .S(_05920_),
    .X(_05931_));
 sky130_fd_sc_hd__xnor2_1 _10108_ (.A(_05930_),
    .B(_05931_),
    .Y(_05932_));
 sky130_fd_sc_hd__mux2_1 _10109_ (.A0(\addroundkey_data_o[35] ),
    .A1(_05932_),
    .S(_05872_),
    .X(_05933_));
 sky130_fd_sc_hd__clkbuf_1 _10110_ (.A(_05933_),
    .X(_00188_));
 sky130_fd_sc_hd__clkbuf_4 _10111_ (.A(_05602_),
    .X(_05934_));
 sky130_fd_sc_hd__mux2_1 _10112_ (.A0(net58),
    .A1(\mix1.data_o[36] ),
    .S(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__buf_4 _10113_ (.A(_05608_),
    .X(_05936_));
 sky130_fd_sc_hd__mux2_1 _10114_ (.A0(\sub1.data_o[36] ),
    .A1(_05935_),
    .S(_05936_),
    .X(_05937_));
 sky130_fd_sc_hd__a31o_1 _10115_ (.A1(_05913_),
    .A2(_05754_),
    .A3(\sub1.data_o[36] ),
    .B1(_05902_),
    .X(_05938_));
 sky130_fd_sc_hd__a21o_1 _10116_ (.A1(_05575_),
    .A2(_05937_),
    .B1(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__o21a_1 _10117_ (.A1(\mix1.data_o[36] ),
    .A2(_05576_),
    .B1(_05916_),
    .X(_05940_));
 sky130_fd_sc_hd__clkbuf_4 _10118_ (.A(_04610_),
    .X(_05941_));
 sky130_fd_sc_hd__a221o_1 _10119_ (.A1(\sub1.data_o[36] ),
    .A2(_05753_),
    .B1(_05939_),
    .B2(_05940_),
    .C1(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__o21ai_4 _10120_ (.A1(_05899_),
    .A2(_05937_),
    .B1(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__mux2_2 _10121_ (.A0(net187),
    .A1(\ks1.key_reg[36] ),
    .S(_05920_),
    .X(_05944_));
 sky130_fd_sc_hd__xnor2_1 _10122_ (.A(_05943_),
    .B(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__mux2_1 _10123_ (.A0(\addroundkey_data_o[36] ),
    .A1(_05945_),
    .S(_05872_),
    .X(_05946_));
 sky130_fd_sc_hd__clkbuf_1 _10124_ (.A(_05946_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _10125_ (.A0(net59),
    .A1(\mix1.data_o[37] ),
    .S(_05934_),
    .X(_05947_));
 sky130_fd_sc_hd__mux2_1 _10126_ (.A0(\sub1.data_o[37] ),
    .A1(_05947_),
    .S(_05936_),
    .X(_05948_));
 sky130_fd_sc_hd__clkbuf_4 _10127_ (.A(_05574_),
    .X(_05949_));
 sky130_fd_sc_hd__a31o_1 _10128_ (.A1(_05913_),
    .A2(_05754_),
    .A3(\sub1.data_o[37] ),
    .B1(_05902_),
    .X(_05950_));
 sky130_fd_sc_hd__a21o_1 _10129_ (.A1(_05949_),
    .A2(_05948_),
    .B1(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__clkbuf_4 _10130_ (.A(_04626_),
    .X(_05952_));
 sky130_fd_sc_hd__o21a_1 _10131_ (.A1(\mix1.data_o[37] ),
    .A2(_05952_),
    .B1(_05916_),
    .X(_05953_));
 sky130_fd_sc_hd__a221o_1 _10132_ (.A1(\sub1.data_o[37] ),
    .A2(_05753_),
    .B1(_05951_),
    .B2(_05953_),
    .C1(_05941_),
    .X(_05954_));
 sky130_fd_sc_hd__o21ai_1 _10133_ (.A1(_05899_),
    .A2(_05948_),
    .B1(_05954_),
    .Y(_05955_));
 sky130_fd_sc_hd__mux2_4 _10134_ (.A0(net188),
    .A1(\ks1.key_reg[37] ),
    .S(_05920_),
    .X(_05956_));
 sky130_fd_sc_hd__xnor2_1 _10135_ (.A(_05955_),
    .B(_05956_),
    .Y(_05957_));
 sky130_fd_sc_hd__mux2_1 _10136_ (.A0(\addroundkey_data_o[37] ),
    .A1(_05957_),
    .S(_05872_),
    .X(_05958_));
 sky130_fd_sc_hd__clkbuf_1 _10137_ (.A(_05958_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _10138_ (.A0(net60),
    .A1(\mix1.data_o[38] ),
    .S(_05934_),
    .X(_05959_));
 sky130_fd_sc_hd__mux2_1 _10139_ (.A0(\sub1.data_o[38] ),
    .A1(_05959_),
    .S(_05936_),
    .X(_05960_));
 sky130_fd_sc_hd__a31o_1 _10140_ (.A1(_05913_),
    .A2(_05754_),
    .A3(\sub1.data_o[38] ),
    .B1(_05902_),
    .X(_05961_));
 sky130_fd_sc_hd__a21o_1 _10141_ (.A1(_05949_),
    .A2(_05960_),
    .B1(_05961_),
    .X(_05962_));
 sky130_fd_sc_hd__o21a_1 _10142_ (.A1(\mix1.data_o[38] ),
    .A2(_05952_),
    .B1(_05916_),
    .X(_05963_));
 sky130_fd_sc_hd__a221o_1 _10143_ (.A1(\sub1.data_o[38] ),
    .A2(_05753_),
    .B1(_05962_),
    .B2(_05963_),
    .C1(_05941_),
    .X(_05964_));
 sky130_fd_sc_hd__o21ai_2 _10144_ (.A1(_05899_),
    .A2(_05960_),
    .B1(_05964_),
    .Y(_05965_));
 sky130_fd_sc_hd__mux2_4 _10145_ (.A0(net189),
    .A1(\ks1.key_reg[38] ),
    .S(_05920_),
    .X(_05966_));
 sky130_fd_sc_hd__xnor2_1 _10146_ (.A(_05965_),
    .B(_05966_),
    .Y(_05967_));
 sky130_fd_sc_hd__mux2_1 _10147_ (.A0(\addroundkey_data_o[38] ),
    .A1(_05967_),
    .S(_05872_),
    .X(_05968_));
 sky130_fd_sc_hd__clkbuf_1 _10148_ (.A(_05968_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _10149_ (.A0(net61),
    .A1(\mix1.data_o[39] ),
    .S(_05934_),
    .X(_05969_));
 sky130_fd_sc_hd__mux2_1 _10150_ (.A0(\sub1.data_o[39] ),
    .A1(_05969_),
    .S(_05936_),
    .X(_05970_));
 sky130_fd_sc_hd__clkbuf_4 _10151_ (.A(_05613_),
    .X(_05971_));
 sky130_fd_sc_hd__clkbuf_4 _10152_ (.A(\sub1.ready_o ),
    .X(_05972_));
 sky130_fd_sc_hd__a31o_1 _10153_ (.A1(_05913_),
    .A2(_05972_),
    .A3(\sub1.data_o[39] ),
    .B1(_05902_),
    .X(_05973_));
 sky130_fd_sc_hd__a21o_1 _10154_ (.A1(_05949_),
    .A2(_05970_),
    .B1(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__o21a_1 _10155_ (.A1(\mix1.data_o[39] ),
    .A2(_05952_),
    .B1(_05916_),
    .X(_05975_));
 sky130_fd_sc_hd__a221o_1 _10156_ (.A1(\sub1.data_o[39] ),
    .A2(_05971_),
    .B1(_05974_),
    .B2(_05975_),
    .C1(_05941_),
    .X(_05976_));
 sky130_fd_sc_hd__o21ai_4 _10157_ (.A1(_05899_),
    .A2(_05970_),
    .B1(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__mux2_1 _10158_ (.A0(net190),
    .A1(\ks1.key_reg[39] ),
    .S(_05920_),
    .X(_05978_));
 sky130_fd_sc_hd__xnor2_1 _10159_ (.A(_05977_),
    .B(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__buf_4 _10160_ (.A(_05792_),
    .X(_05980_));
 sky130_fd_sc_hd__mux2_1 _10161_ (.A0(\addroundkey_data_o[39] ),
    .A1(_05979_),
    .S(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__clkbuf_1 _10162_ (.A(_05981_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _10163_ (.A0(net63),
    .A1(\mix1.data_o[40] ),
    .S(_05817_),
    .X(_05982_));
 sky130_fd_sc_hd__mux2_1 _10164_ (.A0(\sub1.data_o[40] ),
    .A1(_05982_),
    .S(_05819_),
    .X(_05983_));
 sky130_fd_sc_hd__a32o_1 _10165_ (.A1(\mix1.data_o[40] ),
    .A2(_05876_),
    .A3(_05821_),
    .B1(_05822_),
    .B2(\sub1.data_o[40] ),
    .X(_05984_));
 sky130_fd_sc_hd__a22o_1 _10166_ (.A1(_05829_),
    .A2(_05983_),
    .B1(_05984_),
    .B2(_05833_),
    .X(_05985_));
 sky130_fd_sc_hd__mux2_1 _10167_ (.A0(net192),
    .A1(\ks1.key_reg[40] ),
    .S(_05825_),
    .X(_05986_));
 sky130_fd_sc_hd__xor2_1 _10168_ (.A(_05985_),
    .B(_05986_),
    .X(_05987_));
 sky130_fd_sc_hd__mux2_1 _10169_ (.A0(\addroundkey_data_o[40] ),
    .A1(_05987_),
    .S(_05980_),
    .X(_05988_));
 sky130_fd_sc_hd__clkbuf_1 _10170_ (.A(_05988_),
    .X(_00193_));
 sky130_fd_sc_hd__buf_4 _10171_ (.A(_05603_),
    .X(_05989_));
 sky130_fd_sc_hd__mux2_1 _10172_ (.A0(net64),
    .A1(\mix1.data_o[41] ),
    .S(_05989_),
    .X(_05990_));
 sky130_fd_sc_hd__clkbuf_4 _10173_ (.A(_05609_),
    .X(_05991_));
 sky130_fd_sc_hd__mux2_1 _10174_ (.A0(\sub1.data_o[41] ),
    .A1(_05990_),
    .S(_05991_),
    .X(_05992_));
 sky130_fd_sc_hd__buf_2 _10175_ (.A(_05757_),
    .X(_05993_));
 sky130_fd_sc_hd__buf_2 _10176_ (.A(_05620_),
    .X(_05994_));
 sky130_fd_sc_hd__a32o_1 _10177_ (.A1(\mix1.data_o[41] ),
    .A2(_05876_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[41] ),
    .X(_05995_));
 sky130_fd_sc_hd__a22o_1 _10178_ (.A1(_05829_),
    .A2(_05992_),
    .B1(_05995_),
    .B2(_05833_),
    .X(_05996_));
 sky130_fd_sc_hd__buf_4 _10179_ (.A(_05707_),
    .X(_05997_));
 sky130_fd_sc_hd__mux2_1 _10180_ (.A0(net193),
    .A1(\ks1.key_reg[41] ),
    .S(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__xor2_1 _10181_ (.A(_05996_),
    .B(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__mux2_1 _10182_ (.A0(\addroundkey_data_o[41] ),
    .A1(_05999_),
    .S(_05980_),
    .X(_06000_));
 sky130_fd_sc_hd__clkbuf_1 _10183_ (.A(_06000_),
    .X(_00194_));
 sky130_fd_sc_hd__buf_2 _10184_ (.A(_05615_),
    .X(_06001_));
 sky130_fd_sc_hd__mux2_1 _10185_ (.A0(net65),
    .A1(\mix1.data_o[42] ),
    .S(_05989_),
    .X(_06002_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(\sub1.data_o[42] ),
    .A1(_06002_),
    .S(_05991_),
    .X(_06003_));
 sky130_fd_sc_hd__a32o_1 _10187_ (.A1(\mix1.data_o[42] ),
    .A2(_05876_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[42] ),
    .X(_06004_));
 sky130_fd_sc_hd__clkbuf_4 _10188_ (.A(_04609_),
    .X(_06005_));
 sky130_fd_sc_hd__a22o_1 _10189_ (.A1(_06001_),
    .A2(_06003_),
    .B1(_06004_),
    .B2(_06005_),
    .X(_06006_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(net194),
    .A1(\ks1.key_reg[42] ),
    .S(_05997_),
    .X(_06007_));
 sky130_fd_sc_hd__xor2_1 _10191_ (.A(_06006_),
    .B(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(\addroundkey_data_o[42] ),
    .A1(_06008_),
    .S(_05980_),
    .X(_06009_));
 sky130_fd_sc_hd__clkbuf_1 _10193_ (.A(_06009_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _10194_ (.A0(net66),
    .A1(\mix1.data_o[43] ),
    .S(_05989_),
    .X(_06010_));
 sky130_fd_sc_hd__mux2_1 _10195_ (.A0(\sub1.data_o[43] ),
    .A1(_06010_),
    .S(_05991_),
    .X(_06011_));
 sky130_fd_sc_hd__a32o_1 _10196_ (.A1(\mix1.data_o[43] ),
    .A2(_05876_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[43] ),
    .X(_06012_));
 sky130_fd_sc_hd__a22o_1 _10197_ (.A1(_06001_),
    .A2(_06011_),
    .B1(_06012_),
    .B2(_06005_),
    .X(_06013_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(net195),
    .A1(\ks1.key_reg[43] ),
    .S(_05997_),
    .X(_06014_));
 sky130_fd_sc_hd__xor2_1 _10199_ (.A(_06013_),
    .B(_06014_),
    .X(_06015_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(\addroundkey_data_o[43] ),
    .A1(_06015_),
    .S(_05980_),
    .X(_06016_));
 sky130_fd_sc_hd__clkbuf_1 _10201_ (.A(_06016_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(net67),
    .A1(\mix1.data_o[44] ),
    .S(_05989_),
    .X(_06017_));
 sky130_fd_sc_hd__mux2_1 _10203_ (.A0(\sub1.data_o[44] ),
    .A1(_06017_),
    .S(_05991_),
    .X(_06018_));
 sky130_fd_sc_hd__a32o_1 _10204_ (.A1(\mix1.data_o[44] ),
    .A2(_05876_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[44] ),
    .X(_06019_));
 sky130_fd_sc_hd__a22o_1 _10205_ (.A1(_06001_),
    .A2(_06018_),
    .B1(_06019_),
    .B2(_06005_),
    .X(_06020_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(net196),
    .A1(\ks1.key_reg[44] ),
    .S(_05997_),
    .X(_06021_));
 sky130_fd_sc_hd__xor2_1 _10207_ (.A(_06020_),
    .B(_06021_),
    .X(_06022_));
 sky130_fd_sc_hd__mux2_1 _10208_ (.A0(\addroundkey_data_o[44] ),
    .A1(_06022_),
    .S(_05980_),
    .X(_06023_));
 sky130_fd_sc_hd__clkbuf_1 _10209_ (.A(_06023_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _10210_ (.A0(net68),
    .A1(\mix1.data_o[45] ),
    .S(_05989_),
    .X(_06024_));
 sky130_fd_sc_hd__mux2_1 _10211_ (.A0(\sub1.data_o[45] ),
    .A1(_06024_),
    .S(_05991_),
    .X(_06025_));
 sky130_fd_sc_hd__a32o_1 _10212_ (.A1(\mix1.data_o[45] ),
    .A2(_05876_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[45] ),
    .X(_06026_));
 sky130_fd_sc_hd__a22o_1 _10213_ (.A1(_06001_),
    .A2(_06025_),
    .B1(_06026_),
    .B2(_06005_),
    .X(_06027_));
 sky130_fd_sc_hd__mux2_1 _10214_ (.A0(net197),
    .A1(\ks1.key_reg[45] ),
    .S(_05997_),
    .X(_06028_));
 sky130_fd_sc_hd__xor2_1 _10215_ (.A(_06027_),
    .B(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__mux2_1 _10216_ (.A0(\addroundkey_data_o[45] ),
    .A1(_06029_),
    .S(_05980_),
    .X(_06030_));
 sky130_fd_sc_hd__clkbuf_1 _10217_ (.A(_06030_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _10218_ (.A0(net69),
    .A1(\mix1.data_o[46] ),
    .S(_05989_),
    .X(_06031_));
 sky130_fd_sc_hd__mux2_1 _10219_ (.A0(\sub1.data_o[46] ),
    .A1(_06031_),
    .S(_05991_),
    .X(_06032_));
 sky130_fd_sc_hd__a32o_1 _10220_ (.A1(\mix1.data_o[46] ),
    .A2(_05876_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[46] ),
    .X(_06033_));
 sky130_fd_sc_hd__a22o_1 _10221_ (.A1(_06001_),
    .A2(_06032_),
    .B1(_06033_),
    .B2(_06005_),
    .X(_06034_));
 sky130_fd_sc_hd__mux2_1 _10222_ (.A0(net198),
    .A1(\ks1.key_reg[46] ),
    .S(_05997_),
    .X(_06035_));
 sky130_fd_sc_hd__xor2_1 _10223_ (.A(_06034_),
    .B(_06035_),
    .X(_06036_));
 sky130_fd_sc_hd__mux2_1 _10224_ (.A0(\addroundkey_data_o[46] ),
    .A1(_06036_),
    .S(_05980_),
    .X(_06037_));
 sky130_fd_sc_hd__clkbuf_1 _10225_ (.A(_06037_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _10226_ (.A0(net70),
    .A1(\mix1.data_o[47] ),
    .S(_05989_),
    .X(_06038_));
 sky130_fd_sc_hd__mux2_1 _10227_ (.A0(\sub1.data_o[47] ),
    .A1(_06038_),
    .S(_05991_),
    .X(_06039_));
 sky130_fd_sc_hd__a32o_1 _10228_ (.A1(\mix1.data_o[47] ),
    .A2(_05876_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[47] ),
    .X(_06040_));
 sky130_fd_sc_hd__a22o_1 _10229_ (.A1(_06001_),
    .A2(_06039_),
    .B1(_06040_),
    .B2(_06005_),
    .X(_06041_));
 sky130_fd_sc_hd__mux2_1 _10230_ (.A0(net199),
    .A1(\ks1.key_reg[47] ),
    .S(_05997_),
    .X(_06042_));
 sky130_fd_sc_hd__xor2_1 _10231_ (.A(_06041_),
    .B(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__mux2_1 _10232_ (.A0(\addroundkey_data_o[47] ),
    .A1(_06043_),
    .S(_05980_),
    .X(_06044_));
 sky130_fd_sc_hd__clkbuf_1 _10233_ (.A(_06044_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _10234_ (.A0(net71),
    .A1(\mix1.data_o[48] ),
    .S(_05934_),
    .X(_06045_));
 sky130_fd_sc_hd__mux2_1 _10235_ (.A0(\sub1.data_o[48] ),
    .A1(_06045_),
    .S(_05936_),
    .X(_06046_));
 sky130_fd_sc_hd__a31o_1 _10236_ (.A1(_05913_),
    .A2(_05972_),
    .A3(\sub1.data_o[48] ),
    .B1(_05902_),
    .X(_06047_));
 sky130_fd_sc_hd__a21o_1 _10237_ (.A1(_05949_),
    .A2(_06046_),
    .B1(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__o21a_1 _10238_ (.A1(\mix1.data_o[48] ),
    .A2(_05952_),
    .B1(_05916_),
    .X(_06049_));
 sky130_fd_sc_hd__a221o_1 _10239_ (.A1(\sub1.data_o[48] ),
    .A2(_05971_),
    .B1(_06048_),
    .B2(_06049_),
    .C1(_05941_),
    .X(_06050_));
 sky130_fd_sc_hd__o21ai_4 _10240_ (.A1(_05899_),
    .A2(_06046_),
    .B1(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__mux2_1 _10241_ (.A0(net200),
    .A1(\ks1.key_reg[48] ),
    .S(_05920_),
    .X(_06052_));
 sky130_fd_sc_hd__xnor2_1 _10242_ (.A(_06051_),
    .B(_06052_),
    .Y(_06053_));
 sky130_fd_sc_hd__mux2_1 _10243_ (.A0(\addroundkey_data_o[48] ),
    .A1(_06053_),
    .S(_05980_),
    .X(_06054_));
 sky130_fd_sc_hd__clkbuf_1 _10244_ (.A(_06054_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _10245_ (.A0(net72),
    .A1(\mix1.data_o[49] ),
    .S(_05934_),
    .X(_06055_));
 sky130_fd_sc_hd__mux2_1 _10246_ (.A0(\sub1.data_o[49] ),
    .A1(_06055_),
    .S(_05936_),
    .X(_06056_));
 sky130_fd_sc_hd__a31o_1 _10247_ (.A1(_05913_),
    .A2(_05972_),
    .A3(\sub1.data_o[49] ),
    .B1(_05902_),
    .X(_06057_));
 sky130_fd_sc_hd__a21o_1 _10248_ (.A1(_05949_),
    .A2(_06056_),
    .B1(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__o21a_1 _10249_ (.A1(\mix1.data_o[49] ),
    .A2(_05952_),
    .B1(_05916_),
    .X(_06059_));
 sky130_fd_sc_hd__a221o_1 _10250_ (.A1(\sub1.data_o[49] ),
    .A2(_05971_),
    .B1(_06058_),
    .B2(_06059_),
    .C1(_05941_),
    .X(_06060_));
 sky130_fd_sc_hd__o21ai_1 _10251_ (.A1(_05899_),
    .A2(_06056_),
    .B1(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__mux2_4 _10252_ (.A0(net201),
    .A1(\ks1.key_reg[49] ),
    .S(_05920_),
    .X(_06062_));
 sky130_fd_sc_hd__xnor2_1 _10253_ (.A(_06061_),
    .B(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__clkbuf_8 _10254_ (.A(_05792_),
    .X(_06064_));
 sky130_fd_sc_hd__mux2_1 _10255_ (.A0(\addroundkey_data_o[49] ),
    .A1(_06063_),
    .S(_06064_),
    .X(_06065_));
 sky130_fd_sc_hd__clkbuf_1 _10256_ (.A(_06065_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _10257_ (.A0(net74),
    .A1(\mix1.data_o[50] ),
    .S(_05934_),
    .X(_06066_));
 sky130_fd_sc_hd__mux2_1 _10258_ (.A0(\sub1.data_o[50] ),
    .A1(_06066_),
    .S(_05936_),
    .X(_06067_));
 sky130_fd_sc_hd__a31o_1 _10259_ (.A1(_05913_),
    .A2(_05972_),
    .A3(\sub1.data_o[50] ),
    .B1(_05902_),
    .X(_06068_));
 sky130_fd_sc_hd__a21o_1 _10260_ (.A1(_05949_),
    .A2(_06067_),
    .B1(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__o21a_1 _10261_ (.A1(\mix1.data_o[50] ),
    .A2(_05952_),
    .B1(_05916_),
    .X(_06070_));
 sky130_fd_sc_hd__a221o_1 _10262_ (.A1(\sub1.data_o[50] ),
    .A2(_05971_),
    .B1(_06069_),
    .B2(_06070_),
    .C1(_05941_),
    .X(_06071_));
 sky130_fd_sc_hd__o21ai_1 _10263_ (.A1(_05899_),
    .A2(_06067_),
    .B1(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__mux2_2 _10264_ (.A0(net203),
    .A1(\ks1.key_reg[50] ),
    .S(_05920_),
    .X(_06073_));
 sky130_fd_sc_hd__xnor2_1 _10265_ (.A(_06072_),
    .B(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__mux2_1 _10266_ (.A0(\addroundkey_data_o[50] ),
    .A1(_06074_),
    .S(_06064_),
    .X(_06075_));
 sky130_fd_sc_hd__clkbuf_1 _10267_ (.A(_06075_),
    .X(_00203_));
 sky130_fd_sc_hd__clkbuf_8 _10268_ (.A(_05567_),
    .X(_06076_));
 sky130_fd_sc_hd__mux2_1 _10269_ (.A0(net75),
    .A1(\mix1.data_o[51] ),
    .S(_05934_),
    .X(_06077_));
 sky130_fd_sc_hd__mux2_1 _10270_ (.A0(\sub1.data_o[51] ),
    .A1(_06077_),
    .S(_05936_),
    .X(_06078_));
 sky130_fd_sc_hd__clkbuf_4 _10271_ (.A(_05584_),
    .X(_06079_));
 sky130_fd_sc_hd__a31o_1 _10272_ (.A1(_05913_),
    .A2(_05972_),
    .A3(\sub1.data_o[51] ),
    .B1(_06079_),
    .X(_06080_));
 sky130_fd_sc_hd__a21o_1 _10273_ (.A1(_05949_),
    .A2(_06078_),
    .B1(_06080_),
    .X(_06081_));
 sky130_fd_sc_hd__o21a_1 _10274_ (.A1(\mix1.data_o[51] ),
    .A2(_05952_),
    .B1(_05916_),
    .X(_06082_));
 sky130_fd_sc_hd__a221o_1 _10275_ (.A1(\sub1.data_o[51] ),
    .A2(_05971_),
    .B1(_06081_),
    .B2(_06082_),
    .C1(_05941_),
    .X(_06083_));
 sky130_fd_sc_hd__o21ai_1 _10276_ (.A1(_06076_),
    .A2(_06078_),
    .B1(_06083_),
    .Y(_06084_));
 sky130_fd_sc_hd__mux2_4 _10277_ (.A0(net204),
    .A1(\ks1.key_reg[51] ),
    .S(_05920_),
    .X(_06085_));
 sky130_fd_sc_hd__xnor2_1 _10278_ (.A(_06084_),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__mux2_1 _10279_ (.A0(\addroundkey_data_o[51] ),
    .A1(_06086_),
    .S(_06064_),
    .X(_06087_));
 sky130_fd_sc_hd__clkbuf_1 _10280_ (.A(_06087_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _10281_ (.A0(net76),
    .A1(\mix1.data_o[52] ),
    .S(_05934_),
    .X(_06088_));
 sky130_fd_sc_hd__mux2_1 _10282_ (.A0(\sub1.data_o[52] ),
    .A1(_06088_),
    .S(_05936_),
    .X(_06089_));
 sky130_fd_sc_hd__clkbuf_4 _10283_ (.A(_04624_),
    .X(_06090_));
 sky130_fd_sc_hd__a31o_1 _10284_ (.A1(_06090_),
    .A2(_05972_),
    .A3(\sub1.data_o[52] ),
    .B1(_06079_),
    .X(_06091_));
 sky130_fd_sc_hd__a21o_1 _10285_ (.A1(_05949_),
    .A2(_06089_),
    .B1(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_4 _10286_ (.A(_05757_),
    .X(_06093_));
 sky130_fd_sc_hd__o21a_1 _10287_ (.A1(\mix1.data_o[52] ),
    .A2(_05952_),
    .B1(_06093_),
    .X(_06094_));
 sky130_fd_sc_hd__a221o_1 _10288_ (.A1(\sub1.data_o[52] ),
    .A2(_05971_),
    .B1(_06092_),
    .B2(_06094_),
    .C1(_05941_),
    .X(_06095_));
 sky130_fd_sc_hd__o21ai_4 _10289_ (.A1(_06076_),
    .A2(_06089_),
    .B1(_06095_),
    .Y(_06096_));
 sky130_fd_sc_hd__clkbuf_8 _10290_ (.A(_05707_),
    .X(_06097_));
 sky130_fd_sc_hd__mux2_1 _10291_ (.A0(net205),
    .A1(\ks1.key_reg[52] ),
    .S(_06097_),
    .X(_06098_));
 sky130_fd_sc_hd__xnor2_1 _10292_ (.A(_06096_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__mux2_1 _10293_ (.A0(\addroundkey_data_o[52] ),
    .A1(_06099_),
    .S(_06064_),
    .X(_06100_));
 sky130_fd_sc_hd__clkbuf_1 _10294_ (.A(_06100_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _10295_ (.A0(net77),
    .A1(\mix1.data_o[53] ),
    .S(_05934_),
    .X(_06101_));
 sky130_fd_sc_hd__mux2_1 _10296_ (.A0(\sub1.data_o[53] ),
    .A1(_06101_),
    .S(_05936_),
    .X(_06102_));
 sky130_fd_sc_hd__a31o_1 _10297_ (.A1(_06090_),
    .A2(_05972_),
    .A3(\sub1.data_o[53] ),
    .B1(_06079_),
    .X(_06103_));
 sky130_fd_sc_hd__a21o_1 _10298_ (.A1(_05949_),
    .A2(_06102_),
    .B1(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__o21a_1 _10299_ (.A1(\mix1.data_o[53] ),
    .A2(_05952_),
    .B1(_06093_),
    .X(_06105_));
 sky130_fd_sc_hd__a221o_1 _10300_ (.A1(\sub1.data_o[53] ),
    .A2(_05971_),
    .B1(_06104_),
    .B2(_06105_),
    .C1(_05941_),
    .X(_06106_));
 sky130_fd_sc_hd__o21ai_1 _10301_ (.A1(_06076_),
    .A2(_06102_),
    .B1(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__mux2_4 _10302_ (.A0(net206),
    .A1(\ks1.key_reg[53] ),
    .S(_06097_),
    .X(_06108_));
 sky130_fd_sc_hd__xnor2_1 _10303_ (.A(_06107_),
    .B(_06108_),
    .Y(_06109_));
 sky130_fd_sc_hd__mux2_1 _10304_ (.A0(\addroundkey_data_o[53] ),
    .A1(_06109_),
    .S(_06064_),
    .X(_06110_));
 sky130_fd_sc_hd__clkbuf_1 _10305_ (.A(_06110_),
    .X(_00206_));
 sky130_fd_sc_hd__buf_4 _10306_ (.A(_05602_),
    .X(_06111_));
 sky130_fd_sc_hd__mux2_1 _10307_ (.A0(net78),
    .A1(\mix1.data_o[54] ),
    .S(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__buf_4 _10308_ (.A(_05608_),
    .X(_06113_));
 sky130_fd_sc_hd__mux2_1 _10309_ (.A0(\sub1.data_o[54] ),
    .A1(_06112_),
    .S(_06113_),
    .X(_06114_));
 sky130_fd_sc_hd__a31o_1 _10310_ (.A1(_06090_),
    .A2(_05972_),
    .A3(\sub1.data_o[54] ),
    .B1(_06079_),
    .X(_06115_));
 sky130_fd_sc_hd__a21o_1 _10311_ (.A1(_05949_),
    .A2(_06114_),
    .B1(_06115_),
    .X(_06116_));
 sky130_fd_sc_hd__o21a_1 _10312_ (.A1(\mix1.data_o[54] ),
    .A2(_05952_),
    .B1(_06093_),
    .X(_06117_));
 sky130_fd_sc_hd__clkbuf_4 _10313_ (.A(_04610_),
    .X(_06118_));
 sky130_fd_sc_hd__a221o_1 _10314_ (.A1(\sub1.data_o[54] ),
    .A2(_05971_),
    .B1(_06116_),
    .B2(_06117_),
    .C1(_06118_),
    .X(_06119_));
 sky130_fd_sc_hd__o21ai_4 _10315_ (.A1(_06076_),
    .A2(_06114_),
    .B1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__mux2_1 _10316_ (.A0(net207),
    .A1(\ks1.key_reg[54] ),
    .S(_06097_),
    .X(_06121_));
 sky130_fd_sc_hd__xnor2_1 _10317_ (.A(_06120_),
    .B(_06121_),
    .Y(_06122_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(\addroundkey_data_o[54] ),
    .A1(_06122_),
    .S(_06064_),
    .X(_06123_));
 sky130_fd_sc_hd__clkbuf_1 _10319_ (.A(_06123_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _10320_ (.A0(net79),
    .A1(\mix1.data_o[55] ),
    .S(_06111_),
    .X(_06124_));
 sky130_fd_sc_hd__mux2_1 _10321_ (.A0(\sub1.data_o[55] ),
    .A1(_06124_),
    .S(_06113_),
    .X(_06125_));
 sky130_fd_sc_hd__clkbuf_4 _10322_ (.A(_05574_),
    .X(_06126_));
 sky130_fd_sc_hd__a31o_1 _10323_ (.A1(_06090_),
    .A2(_05972_),
    .A3(\sub1.data_o[55] ),
    .B1(_06079_),
    .X(_06127_));
 sky130_fd_sc_hd__a21o_1 _10324_ (.A1(_06126_),
    .A2(_06125_),
    .B1(_06127_),
    .X(_06128_));
 sky130_fd_sc_hd__clkbuf_4 _10325_ (.A(_04626_),
    .X(_06129_));
 sky130_fd_sc_hd__o21a_1 _10326_ (.A1(\mix1.data_o[55] ),
    .A2(_06129_),
    .B1(_06093_),
    .X(_06130_));
 sky130_fd_sc_hd__a221o_1 _10327_ (.A1(\sub1.data_o[55] ),
    .A2(_05971_),
    .B1(_06128_),
    .B2(_06130_),
    .C1(_06118_),
    .X(_06131_));
 sky130_fd_sc_hd__o21ai_2 _10328_ (.A1(_06076_),
    .A2(_06125_),
    .B1(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__mux2_4 _10329_ (.A0(net208),
    .A1(\ks1.key_reg[55] ),
    .S(_06097_),
    .X(_06133_));
 sky130_fd_sc_hd__xnor2_1 _10330_ (.A(_06132_),
    .B(_06133_),
    .Y(_06134_));
 sky130_fd_sc_hd__mux2_1 _10331_ (.A0(\addroundkey_data_o[55] ),
    .A1(_06134_),
    .S(_06064_),
    .X(_06135_));
 sky130_fd_sc_hd__clkbuf_1 _10332_ (.A(_06135_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _10333_ (.A0(net80),
    .A1(\mix1.data_o[56] ),
    .S(_05989_),
    .X(_06136_));
 sky130_fd_sc_hd__mux2_1 _10334_ (.A0(\sub1.data_o[56] ),
    .A1(_06136_),
    .S(_05991_),
    .X(_06137_));
 sky130_fd_sc_hd__clkbuf_4 _10335_ (.A(_05585_),
    .X(_06138_));
 sky130_fd_sc_hd__a32o_1 _10336_ (.A1(\mix1.data_o[56] ),
    .A2(_06138_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[56] ),
    .X(_06139_));
 sky130_fd_sc_hd__a22o_1 _10337_ (.A1(_06001_),
    .A2(_06137_),
    .B1(_06139_),
    .B2(_06005_),
    .X(_06140_));
 sky130_fd_sc_hd__mux2_1 _10338_ (.A0(net209),
    .A1(\ks1.key_reg[56] ),
    .S(_05997_),
    .X(_06141_));
 sky130_fd_sc_hd__xor2_1 _10339_ (.A(_06140_),
    .B(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__mux2_1 _10340_ (.A0(\addroundkey_data_o[56] ),
    .A1(_06142_),
    .S(_06064_),
    .X(_06143_));
 sky130_fd_sc_hd__clkbuf_1 _10341_ (.A(_06143_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _10342_ (.A0(net81),
    .A1(\mix1.data_o[57] ),
    .S(_05989_),
    .X(_06144_));
 sky130_fd_sc_hd__mux2_1 _10343_ (.A0(\sub1.data_o[57] ),
    .A1(_06144_),
    .S(_05991_),
    .X(_06145_));
 sky130_fd_sc_hd__a32o_1 _10344_ (.A1(\mix1.data_o[57] ),
    .A2(_06138_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[57] ),
    .X(_06146_));
 sky130_fd_sc_hd__a22o_1 _10345_ (.A1(_06001_),
    .A2(_06145_),
    .B1(_06146_),
    .B2(_06005_),
    .X(_06147_));
 sky130_fd_sc_hd__mux2_1 _10346_ (.A0(net210),
    .A1(\ks1.key_reg[57] ),
    .S(_05997_),
    .X(_06148_));
 sky130_fd_sc_hd__xor2_1 _10347_ (.A(_06147_),
    .B(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__mux2_1 _10348_ (.A0(\addroundkey_data_o[57] ),
    .A1(_06149_),
    .S(_06064_),
    .X(_06150_));
 sky130_fd_sc_hd__clkbuf_1 _10349_ (.A(_06150_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _10350_ (.A0(net82),
    .A1(\mix1.data_o[58] ),
    .S(_05989_),
    .X(_06151_));
 sky130_fd_sc_hd__mux2_1 _10351_ (.A0(\sub1.data_o[58] ),
    .A1(_06151_),
    .S(_05991_),
    .X(_06152_));
 sky130_fd_sc_hd__a32o_1 _10352_ (.A1(\mix1.data_o[58] ),
    .A2(_06138_),
    .A3(_05993_),
    .B1(_05994_),
    .B2(\sub1.data_o[58] ),
    .X(_06153_));
 sky130_fd_sc_hd__a22o_1 _10353_ (.A1(_06001_),
    .A2(_06152_),
    .B1(_06153_),
    .B2(_06005_),
    .X(_06154_));
 sky130_fd_sc_hd__mux2_1 _10354_ (.A0(net211),
    .A1(\ks1.key_reg[58] ),
    .S(_05997_),
    .X(_06155_));
 sky130_fd_sc_hd__xor2_1 _10355_ (.A(_06154_),
    .B(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__mux2_1 _10356_ (.A0(\addroundkey_data_o[58] ),
    .A1(_06156_),
    .S(_06064_),
    .X(_06157_));
 sky130_fd_sc_hd__clkbuf_1 _10357_ (.A(_06157_),
    .X(_00211_));
 sky130_fd_sc_hd__clkbuf_4 _10358_ (.A(_05603_),
    .X(_06158_));
 sky130_fd_sc_hd__mux2_1 _10359_ (.A0(net83),
    .A1(\mix1.data_o[59] ),
    .S(_06158_),
    .X(_06159_));
 sky130_fd_sc_hd__clkbuf_4 _10360_ (.A(_05609_),
    .X(_06160_));
 sky130_fd_sc_hd__mux2_1 _10361_ (.A0(\sub1.data_o[59] ),
    .A1(_06159_),
    .S(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__clkbuf_4 _10362_ (.A(_05757_),
    .X(_06162_));
 sky130_fd_sc_hd__clkbuf_4 _10363_ (.A(_05620_),
    .X(_06163_));
 sky130_fd_sc_hd__a32o_1 _10364_ (.A1(\mix1.data_o[59] ),
    .A2(_06138_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[59] ),
    .X(_06164_));
 sky130_fd_sc_hd__a22o_1 _10365_ (.A1(_06001_),
    .A2(_06161_),
    .B1(_06164_),
    .B2(_06005_),
    .X(_06165_));
 sky130_fd_sc_hd__clkbuf_4 _10366_ (.A(_05707_),
    .X(_06166_));
 sky130_fd_sc_hd__mux2_1 _10367_ (.A0(net212),
    .A1(\ks1.key_reg[59] ),
    .S(_06166_),
    .X(_06167_));
 sky130_fd_sc_hd__xor2_1 _10368_ (.A(_06165_),
    .B(_06167_),
    .X(_06168_));
 sky130_fd_sc_hd__buf_4 _10369_ (.A(_05792_),
    .X(_06169_));
 sky130_fd_sc_hd__mux2_1 _10370_ (.A0(\addroundkey_data_o[59] ),
    .A1(_06168_),
    .S(_06169_),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_1 _10371_ (.A(_06170_),
    .X(_00212_));
 sky130_fd_sc_hd__clkbuf_4 _10372_ (.A(_05615_),
    .X(_06171_));
 sky130_fd_sc_hd__mux2_1 _10373_ (.A0(net85),
    .A1(\mix1.data_o[60] ),
    .S(_06158_),
    .X(_06172_));
 sky130_fd_sc_hd__mux2_1 _10374_ (.A0(\sub1.data_o[60] ),
    .A1(_06172_),
    .S(_06160_),
    .X(_06173_));
 sky130_fd_sc_hd__a32o_1 _10375_ (.A1(\mix1.data_o[60] ),
    .A2(_06138_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[60] ),
    .X(_06174_));
 sky130_fd_sc_hd__clkbuf_4 _10376_ (.A(_04609_),
    .X(_06175_));
 sky130_fd_sc_hd__a22o_1 _10377_ (.A1(_06171_),
    .A2(_06173_),
    .B1(_06174_),
    .B2(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__mux2_1 _10378_ (.A0(net214),
    .A1(\ks1.key_reg[60] ),
    .S(_06166_),
    .X(_06177_));
 sky130_fd_sc_hd__xor2_1 _10379_ (.A(_06176_),
    .B(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__mux2_1 _10380_ (.A0(\addroundkey_data_o[60] ),
    .A1(_06178_),
    .S(_06169_),
    .X(_06179_));
 sky130_fd_sc_hd__clkbuf_1 _10381_ (.A(_06179_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _10382_ (.A0(net86),
    .A1(\mix1.data_o[61] ),
    .S(_06158_),
    .X(_06180_));
 sky130_fd_sc_hd__mux2_1 _10383_ (.A0(\sub1.data_o[61] ),
    .A1(_06180_),
    .S(_06160_),
    .X(_06181_));
 sky130_fd_sc_hd__a32o_1 _10384_ (.A1(\mix1.data_o[61] ),
    .A2(_06138_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[61] ),
    .X(_06182_));
 sky130_fd_sc_hd__a22o_1 _10385_ (.A1(_06171_),
    .A2(_06181_),
    .B1(_06182_),
    .B2(_06175_),
    .X(_06183_));
 sky130_fd_sc_hd__mux2_1 _10386_ (.A0(net215),
    .A1(\ks1.key_reg[61] ),
    .S(_06166_),
    .X(_06184_));
 sky130_fd_sc_hd__xor2_1 _10387_ (.A(_06183_),
    .B(_06184_),
    .X(_06185_));
 sky130_fd_sc_hd__mux2_1 _10388_ (.A0(\addroundkey_data_o[61] ),
    .A1(_06185_),
    .S(_06169_),
    .X(_06186_));
 sky130_fd_sc_hd__clkbuf_1 _10389_ (.A(_06186_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _10390_ (.A0(net87),
    .A1(\mix1.data_o[62] ),
    .S(_06158_),
    .X(_06187_));
 sky130_fd_sc_hd__mux2_1 _10391_ (.A0(\sub1.data_o[62] ),
    .A1(_06187_),
    .S(_06160_),
    .X(_06188_));
 sky130_fd_sc_hd__a32o_1 _10392_ (.A1(\mix1.data_o[62] ),
    .A2(_06138_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[62] ),
    .X(_06189_));
 sky130_fd_sc_hd__a22o_1 _10393_ (.A1(_06171_),
    .A2(_06188_),
    .B1(_06189_),
    .B2(_06175_),
    .X(_06190_));
 sky130_fd_sc_hd__mux2_1 _10394_ (.A0(net216),
    .A1(\ks1.key_reg[62] ),
    .S(_06166_),
    .X(_06191_));
 sky130_fd_sc_hd__xor2_1 _10395_ (.A(_06190_),
    .B(_06191_),
    .X(_06192_));
 sky130_fd_sc_hd__mux2_1 _10396_ (.A0(\addroundkey_data_o[62] ),
    .A1(_06192_),
    .S(_06169_),
    .X(_06193_));
 sky130_fd_sc_hd__clkbuf_1 _10397_ (.A(_06193_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _10398_ (.A0(net88),
    .A1(\mix1.data_o[63] ),
    .S(_06158_),
    .X(_06194_));
 sky130_fd_sc_hd__mux2_1 _10399_ (.A0(\sub1.data_o[63] ),
    .A1(_06194_),
    .S(_06160_),
    .X(_06195_));
 sky130_fd_sc_hd__a32o_1 _10400_ (.A1(\mix1.data_o[63] ),
    .A2(_06138_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[63] ),
    .X(_06196_));
 sky130_fd_sc_hd__a22o_1 _10401_ (.A1(_06171_),
    .A2(_06195_),
    .B1(_06196_),
    .B2(_06175_),
    .X(_06197_));
 sky130_fd_sc_hd__mux2_2 _10402_ (.A0(net217),
    .A1(\ks1.key_reg[63] ),
    .S(_06166_),
    .X(_06198_));
 sky130_fd_sc_hd__xor2_1 _10403_ (.A(_06197_),
    .B(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__mux2_1 _10404_ (.A0(\addroundkey_data_o[63] ),
    .A1(_06199_),
    .S(_06169_),
    .X(_06200_));
 sky130_fd_sc_hd__clkbuf_1 _10405_ (.A(_06200_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _10406_ (.A0(net89),
    .A1(\mix1.data_o[64] ),
    .S(_06158_),
    .X(_06201_));
 sky130_fd_sc_hd__mux2_1 _10407_ (.A0(\sub1.data_o[64] ),
    .A1(_06201_),
    .S(_06160_),
    .X(_06202_));
 sky130_fd_sc_hd__a32o_1 _10408_ (.A1(\mix1.data_o[64] ),
    .A2(_06138_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[64] ),
    .X(_06203_));
 sky130_fd_sc_hd__a22o_1 _10409_ (.A1(_06171_),
    .A2(_06202_),
    .B1(_06203_),
    .B2(_06175_),
    .X(_06204_));
 sky130_fd_sc_hd__mux2_1 _10410_ (.A0(net218),
    .A1(\ks1.key_reg[64] ),
    .S(_06166_),
    .X(_06205_));
 sky130_fd_sc_hd__xor2_1 _10411_ (.A(_06204_),
    .B(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__mux2_1 _10412_ (.A0(\addroundkey_data_o[64] ),
    .A1(_06206_),
    .S(_06169_),
    .X(_06207_));
 sky130_fd_sc_hd__clkbuf_1 _10413_ (.A(_06207_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _10414_ (.A0(net90),
    .A1(\mix1.data_o[65] ),
    .S(_06158_),
    .X(_06208_));
 sky130_fd_sc_hd__mux2_1 _10415_ (.A0(\sub1.data_o[65] ),
    .A1(_06208_),
    .S(_06160_),
    .X(_06209_));
 sky130_fd_sc_hd__a32o_1 _10416_ (.A1(\mix1.data_o[65] ),
    .A2(_06138_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[65] ),
    .X(_06210_));
 sky130_fd_sc_hd__a22o_1 _10417_ (.A1(_06171_),
    .A2(_06209_),
    .B1(_06210_),
    .B2(_06175_),
    .X(_06211_));
 sky130_fd_sc_hd__mux2_1 _10418_ (.A0(net219),
    .A1(\ks1.key_reg[65] ),
    .S(_06166_),
    .X(_06212_));
 sky130_fd_sc_hd__xor2_1 _10419_ (.A(_06211_),
    .B(_06212_),
    .X(_06213_));
 sky130_fd_sc_hd__mux2_1 _10420_ (.A0(\addroundkey_data_o[65] ),
    .A1(_06213_),
    .S(_06169_),
    .X(_06214_));
 sky130_fd_sc_hd__clkbuf_1 _10421_ (.A(_06214_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _10422_ (.A0(net91),
    .A1(\mix1.data_o[66] ),
    .S(_06158_),
    .X(_06215_));
 sky130_fd_sc_hd__mux2_1 _10423_ (.A0(\sub1.data_o[66] ),
    .A1(_06215_),
    .S(_06160_),
    .X(_06216_));
 sky130_fd_sc_hd__clkbuf_4 _10424_ (.A(_05585_),
    .X(_06217_));
 sky130_fd_sc_hd__a32o_1 _10425_ (.A1(\mix1.data_o[66] ),
    .A2(_06217_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[66] ),
    .X(_06218_));
 sky130_fd_sc_hd__a22o_1 _10426_ (.A1(_06171_),
    .A2(_06216_),
    .B1(_06218_),
    .B2(_06175_),
    .X(_06219_));
 sky130_fd_sc_hd__mux2_1 _10427_ (.A0(net220),
    .A1(\ks1.key_reg[66] ),
    .S(_06166_),
    .X(_06220_));
 sky130_fd_sc_hd__xor2_1 _10428_ (.A(_06219_),
    .B(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__mux2_1 _10429_ (.A0(\addroundkey_data_o[66] ),
    .A1(_06221_),
    .S(_06169_),
    .X(_06222_));
 sky130_fd_sc_hd__clkbuf_1 _10430_ (.A(_06222_),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _10431_ (.A0(net92),
    .A1(\mix1.data_o[67] ),
    .S(_06158_),
    .X(_06223_));
 sky130_fd_sc_hd__mux2_1 _10432_ (.A0(\sub1.data_o[67] ),
    .A1(_06223_),
    .S(_06160_),
    .X(_06224_));
 sky130_fd_sc_hd__a32o_1 _10433_ (.A1(\mix1.data_o[67] ),
    .A2(_06217_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[67] ),
    .X(_06225_));
 sky130_fd_sc_hd__a22o_1 _10434_ (.A1(_06171_),
    .A2(_06224_),
    .B1(_06225_),
    .B2(_06175_),
    .X(_06226_));
 sky130_fd_sc_hd__mux2_1 _10435_ (.A0(net221),
    .A1(\ks1.key_reg[67] ),
    .S(_06166_),
    .X(_06227_));
 sky130_fd_sc_hd__xor2_1 _10436_ (.A(_06226_),
    .B(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(\addroundkey_data_o[67] ),
    .A1(_06228_),
    .S(_06169_),
    .X(_06229_));
 sky130_fd_sc_hd__clkbuf_1 _10438_ (.A(_06229_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _10439_ (.A0(net93),
    .A1(\mix1.data_o[68] ),
    .S(_06158_),
    .X(_06230_));
 sky130_fd_sc_hd__mux2_1 _10440_ (.A0(\sub1.data_o[68] ),
    .A1(_06230_),
    .S(_06160_),
    .X(_06231_));
 sky130_fd_sc_hd__a32o_1 _10441_ (.A1(\mix1.data_o[68] ),
    .A2(_06217_),
    .A3(_06162_),
    .B1(_06163_),
    .B2(\sub1.data_o[68] ),
    .X(_06232_));
 sky130_fd_sc_hd__a22o_1 _10442_ (.A1(_06171_),
    .A2(_06231_),
    .B1(_06232_),
    .B2(_06175_),
    .X(_06233_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(net222),
    .A1(\ks1.key_reg[68] ),
    .S(_06166_),
    .X(_06234_));
 sky130_fd_sc_hd__xor2_1 _10444_ (.A(_06233_),
    .B(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__mux2_1 _10445_ (.A0(\addroundkey_data_o[68] ),
    .A1(_06235_),
    .S(_06169_),
    .X(_06236_));
 sky130_fd_sc_hd__clkbuf_1 _10446_ (.A(_06236_),
    .X(_00221_));
 sky130_fd_sc_hd__buf_4 _10447_ (.A(_05749_),
    .X(_06237_));
 sky130_fd_sc_hd__mux2_1 _10448_ (.A0(net94),
    .A1(\mix1.data_o[69] ),
    .S(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__buf_4 _10449_ (.A(_05751_),
    .X(_06239_));
 sky130_fd_sc_hd__mux2_1 _10450_ (.A0(\sub1.data_o[69] ),
    .A1(_06238_),
    .S(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__clkbuf_4 _10451_ (.A(_05757_),
    .X(_06241_));
 sky130_fd_sc_hd__clkbuf_4 _10452_ (.A(_05619_),
    .X(_06242_));
 sky130_fd_sc_hd__a32o_1 _10453_ (.A1(\mix1.data_o[69] ),
    .A2(_06217_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[69] ),
    .X(_06243_));
 sky130_fd_sc_hd__a22o_2 _10454_ (.A1(_06171_),
    .A2(_06240_),
    .B1(_06243_),
    .B2(_06175_),
    .X(_06244_));
 sky130_fd_sc_hd__clkbuf_4 _10455_ (.A(_05707_),
    .X(_06245_));
 sky130_fd_sc_hd__mux2_1 _10456_ (.A0(net223),
    .A1(\ks1.key_reg[69] ),
    .S(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__xor2_1 _10457_ (.A(_06244_),
    .B(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__buf_4 _10458_ (.A(_05792_),
    .X(_06248_));
 sky130_fd_sc_hd__mux2_1 _10459_ (.A0(\addroundkey_data_o[69] ),
    .A1(_06247_),
    .S(_06248_),
    .X(_06249_));
 sky130_fd_sc_hd__clkbuf_1 _10460_ (.A(_06249_),
    .X(_00222_));
 sky130_fd_sc_hd__clkbuf_4 _10461_ (.A(_05614_),
    .X(_06250_));
 sky130_fd_sc_hd__mux2_1 _10462_ (.A0(net96),
    .A1(\mix1.data_o[70] ),
    .S(_06237_),
    .X(_06251_));
 sky130_fd_sc_hd__mux2_1 _10463_ (.A0(\sub1.data_o[70] ),
    .A1(_06251_),
    .S(_06239_),
    .X(_06252_));
 sky130_fd_sc_hd__a32o_1 _10464_ (.A1(\mix1.data_o[70] ),
    .A2(_06217_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[70] ),
    .X(_06253_));
 sky130_fd_sc_hd__clkbuf_4 _10465_ (.A(_04609_),
    .X(_06254_));
 sky130_fd_sc_hd__a22o_1 _10466_ (.A1(_06250_),
    .A2(_06252_),
    .B1(_06253_),
    .B2(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__mux2_1 _10467_ (.A0(net225),
    .A1(\ks1.key_reg[70] ),
    .S(_06245_),
    .X(_06256_));
 sky130_fd_sc_hd__xor2_1 _10468_ (.A(_06255_),
    .B(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__mux2_1 _10469_ (.A0(\addroundkey_data_o[70] ),
    .A1(_06257_),
    .S(_06248_),
    .X(_06258_));
 sky130_fd_sc_hd__clkbuf_1 _10470_ (.A(_06258_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _10471_ (.A0(net97),
    .A1(\mix1.data_o[71] ),
    .S(_06237_),
    .X(_06259_));
 sky130_fd_sc_hd__mux2_1 _10472_ (.A0(\sub1.data_o[71] ),
    .A1(_06259_),
    .S(_06239_),
    .X(_06260_));
 sky130_fd_sc_hd__a32o_1 _10473_ (.A1(\mix1.data_o[71] ),
    .A2(_06217_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[71] ),
    .X(_06261_));
 sky130_fd_sc_hd__a22o_1 _10474_ (.A1(_06250_),
    .A2(_06260_),
    .B1(_06261_),
    .B2(_06254_),
    .X(_06262_));
 sky130_fd_sc_hd__mux2_1 _10475_ (.A0(net226),
    .A1(\ks1.key_reg[71] ),
    .S(_06245_),
    .X(_06263_));
 sky130_fd_sc_hd__xor2_1 _10476_ (.A(_06262_),
    .B(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(\addroundkey_data_o[71] ),
    .A1(_06264_),
    .S(_06248_),
    .X(_06265_));
 sky130_fd_sc_hd__clkbuf_1 _10478_ (.A(_06265_),
    .X(_00224_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(net98),
    .A1(\mix1.data_o[72] ),
    .S(_06237_),
    .X(_06266_));
 sky130_fd_sc_hd__mux2_1 _10480_ (.A0(\sub1.data_o[72] ),
    .A1(_06266_),
    .S(_06239_),
    .X(_06267_));
 sky130_fd_sc_hd__a32o_1 _10481_ (.A1(\mix1.data_o[72] ),
    .A2(_06217_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[72] ),
    .X(_06268_));
 sky130_fd_sc_hd__a22o_1 _10482_ (.A1(_06250_),
    .A2(_06267_),
    .B1(_06268_),
    .B2(_06254_),
    .X(_06269_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(net227),
    .A1(\ks1.key_reg[72] ),
    .S(_06245_),
    .X(_06270_));
 sky130_fd_sc_hd__xor2_1 _10484_ (.A(_06269_),
    .B(_06270_),
    .X(_06271_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(\addroundkey_data_o[72] ),
    .A1(_06271_),
    .S(_06248_),
    .X(_06272_));
 sky130_fd_sc_hd__clkbuf_1 _10486_ (.A(_06272_),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(net99),
    .A1(\mix1.data_o[73] ),
    .S(_06237_),
    .X(_06273_));
 sky130_fd_sc_hd__mux2_1 _10488_ (.A0(\sub1.data_o[73] ),
    .A1(_06273_),
    .S(_06239_),
    .X(_06274_));
 sky130_fd_sc_hd__a32o_1 _10489_ (.A1(\mix1.data_o[73] ),
    .A2(_06217_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[73] ),
    .X(_06275_));
 sky130_fd_sc_hd__a22o_1 _10490_ (.A1(_06250_),
    .A2(_06274_),
    .B1(_06275_),
    .B2(_06254_),
    .X(_06276_));
 sky130_fd_sc_hd__mux2_2 _10491_ (.A0(net228),
    .A1(\ks1.key_reg[73] ),
    .S(_06245_),
    .X(_06277_));
 sky130_fd_sc_hd__xor2_1 _10492_ (.A(_06276_),
    .B(_06277_),
    .X(_06278_));
 sky130_fd_sc_hd__mux2_1 _10493_ (.A0(\addroundkey_data_o[73] ),
    .A1(_06278_),
    .S(_06248_),
    .X(_06279_));
 sky130_fd_sc_hd__clkbuf_1 _10494_ (.A(_06279_),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _10495_ (.A0(net100),
    .A1(\mix1.data_o[74] ),
    .S(_06237_),
    .X(_06280_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(\sub1.data_o[74] ),
    .A1(_06280_),
    .S(_06239_),
    .X(_06281_));
 sky130_fd_sc_hd__a32o_1 _10497_ (.A1(\mix1.data_o[74] ),
    .A2(_06217_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[74] ),
    .X(_06282_));
 sky130_fd_sc_hd__a22o_1 _10498_ (.A1(_06250_),
    .A2(_06281_),
    .B1(_06282_),
    .B2(_06254_),
    .X(_06283_));
 sky130_fd_sc_hd__mux2_1 _10499_ (.A0(net229),
    .A1(\ks1.key_reg[74] ),
    .S(_06245_),
    .X(_06284_));
 sky130_fd_sc_hd__xor2_1 _10500_ (.A(_06283_),
    .B(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(\addroundkey_data_o[74] ),
    .A1(_06285_),
    .S(_06248_),
    .X(_06286_));
 sky130_fd_sc_hd__clkbuf_1 _10502_ (.A(_06286_),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _10503_ (.A0(net101),
    .A1(\mix1.data_o[75] ),
    .S(_06237_),
    .X(_06287_));
 sky130_fd_sc_hd__mux2_1 _10504_ (.A0(\sub1.data_o[75] ),
    .A1(_06287_),
    .S(_06239_),
    .X(_06288_));
 sky130_fd_sc_hd__a32o_1 _10505_ (.A1(\mix1.data_o[75] ),
    .A2(_06217_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[75] ),
    .X(_06289_));
 sky130_fd_sc_hd__a22o_1 _10506_ (.A1(_06250_),
    .A2(_06288_),
    .B1(_06289_),
    .B2(_06254_),
    .X(_06290_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(net230),
    .A1(\ks1.key_reg[75] ),
    .S(_06245_),
    .X(_06291_));
 sky130_fd_sc_hd__xor2_1 _10508_ (.A(_06290_),
    .B(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__mux2_1 _10509_ (.A0(\addroundkey_data_o[75] ),
    .A1(_06292_),
    .S(_06248_),
    .X(_06293_));
 sky130_fd_sc_hd__clkbuf_1 _10510_ (.A(_06293_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(net102),
    .A1(\mix1.data_o[76] ),
    .S(_06237_),
    .X(_06294_));
 sky130_fd_sc_hd__mux2_1 _10512_ (.A0(\sub1.data_o[76] ),
    .A1(_06294_),
    .S(_06239_),
    .X(_06295_));
 sky130_fd_sc_hd__clkbuf_4 _10513_ (.A(_05585_),
    .X(_06296_));
 sky130_fd_sc_hd__a32o_1 _10514_ (.A1(\mix1.data_o[76] ),
    .A2(_06296_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[76] ),
    .X(_06297_));
 sky130_fd_sc_hd__a22o_2 _10515_ (.A1(_06250_),
    .A2(_06295_),
    .B1(_06297_),
    .B2(_06254_),
    .X(_06298_));
 sky130_fd_sc_hd__mux2_1 _10516_ (.A0(net231),
    .A1(\ks1.key_reg[76] ),
    .S(_06245_),
    .X(_06299_));
 sky130_fd_sc_hd__xor2_1 _10517_ (.A(_06298_),
    .B(_06299_),
    .X(_06300_));
 sky130_fd_sc_hd__mux2_1 _10518_ (.A0(\addroundkey_data_o[76] ),
    .A1(_06300_),
    .S(_06248_),
    .X(_06301_));
 sky130_fd_sc_hd__clkbuf_1 _10519_ (.A(_06301_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _10520_ (.A0(net103),
    .A1(\mix1.data_o[77] ),
    .S(_06237_),
    .X(_06302_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(\sub1.data_o[77] ),
    .A1(_06302_),
    .S(_06239_),
    .X(_06303_));
 sky130_fd_sc_hd__a32o_1 _10522_ (.A1(\mix1.data_o[77] ),
    .A2(_06296_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[77] ),
    .X(_06304_));
 sky130_fd_sc_hd__a22o_1 _10523_ (.A1(_06250_),
    .A2(_06303_),
    .B1(_06304_),
    .B2(_06254_),
    .X(_06305_));
 sky130_fd_sc_hd__mux2_1 _10524_ (.A0(net232),
    .A1(\ks1.key_reg[77] ),
    .S(_06245_),
    .X(_06306_));
 sky130_fd_sc_hd__xor2_1 _10525_ (.A(_06305_),
    .B(_06306_),
    .X(_06307_));
 sky130_fd_sc_hd__mux2_1 _10526_ (.A0(\addroundkey_data_o[77] ),
    .A1(_06307_),
    .S(_06248_),
    .X(_06308_));
 sky130_fd_sc_hd__clkbuf_1 _10527_ (.A(_06308_),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _10528_ (.A0(net104),
    .A1(\mix1.data_o[78] ),
    .S(_06237_),
    .X(_06309_));
 sky130_fd_sc_hd__mux2_1 _10529_ (.A0(\sub1.data_o[78] ),
    .A1(_06309_),
    .S(_06239_),
    .X(_06310_));
 sky130_fd_sc_hd__a32o_1 _10530_ (.A1(\mix1.data_o[78] ),
    .A2(_06296_),
    .A3(_06241_),
    .B1(_06242_),
    .B2(\sub1.data_o[78] ),
    .X(_06311_));
 sky130_fd_sc_hd__a22o_2 _10531_ (.A1(_06250_),
    .A2(_06310_),
    .B1(_06311_),
    .B2(_06254_),
    .X(_06312_));
 sky130_fd_sc_hd__mux2_1 _10532_ (.A0(net233),
    .A1(\ks1.key_reg[78] ),
    .S(_06245_),
    .X(_06313_));
 sky130_fd_sc_hd__xor2_1 _10533_ (.A(_06312_),
    .B(_06313_),
    .X(_06314_));
 sky130_fd_sc_hd__mux2_1 _10534_ (.A0(\addroundkey_data_o[78] ),
    .A1(_06314_),
    .S(_06248_),
    .X(_06315_));
 sky130_fd_sc_hd__clkbuf_1 _10535_ (.A(_06315_),
    .X(_00231_));
 sky130_fd_sc_hd__buf_4 _10536_ (.A(_05749_),
    .X(_06316_));
 sky130_fd_sc_hd__mux2_1 _10537_ (.A0(net105),
    .A1(\mix1.data_o[79] ),
    .S(_06316_),
    .X(_06317_));
 sky130_fd_sc_hd__clkbuf_4 _10538_ (.A(_05751_),
    .X(_06318_));
 sky130_fd_sc_hd__mux2_1 _10539_ (.A0(\sub1.data_o[79] ),
    .A1(_06317_),
    .S(_06318_),
    .X(_06319_));
 sky130_fd_sc_hd__clkbuf_4 _10540_ (.A(_05757_),
    .X(_06320_));
 sky130_fd_sc_hd__clkbuf_4 _10541_ (.A(_05619_),
    .X(_06321_));
 sky130_fd_sc_hd__a32o_1 _10542_ (.A1(\mix1.data_o[79] ),
    .A2(_06296_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[79] ),
    .X(_06322_));
 sky130_fd_sc_hd__a22o_1 _10543_ (.A1(_06250_),
    .A2(_06319_),
    .B1(_06322_),
    .B2(_06254_),
    .X(_06323_));
 sky130_fd_sc_hd__buf_4 _10544_ (.A(_05707_),
    .X(_06324_));
 sky130_fd_sc_hd__mux2_2 _10545_ (.A0(net234),
    .A1(\ks1.key_reg[79] ),
    .S(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__xor2_1 _10546_ (.A(_06323_),
    .B(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__buf_6 _10547_ (.A(_05792_),
    .X(_06327_));
 sky130_fd_sc_hd__mux2_1 _10548_ (.A0(\addroundkey_data_o[79] ),
    .A1(_06326_),
    .S(_06327_),
    .X(_06328_));
 sky130_fd_sc_hd__clkbuf_1 _10549_ (.A(_06328_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _10550_ (.A0(net107),
    .A1(\mix1.data_o[80] ),
    .S(_06111_),
    .X(_06329_));
 sky130_fd_sc_hd__mux2_1 _10551_ (.A0(\sub1.data_o[80] ),
    .A1(_06329_),
    .S(_06113_),
    .X(_06330_));
 sky130_fd_sc_hd__a31o_1 _10552_ (.A1(_06090_),
    .A2(_05972_),
    .A3(\sub1.data_o[80] ),
    .B1(_06079_),
    .X(_06331_));
 sky130_fd_sc_hd__a21o_1 _10553_ (.A1(_06126_),
    .A2(_06330_),
    .B1(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__o21a_1 _10554_ (.A1(\mix1.data_o[80] ),
    .A2(_06129_),
    .B1(_06093_),
    .X(_06333_));
 sky130_fd_sc_hd__a221o_1 _10555_ (.A1(\sub1.data_o[80] ),
    .A2(_05971_),
    .B1(_06332_),
    .B2(_06333_),
    .C1(_06118_),
    .X(_06334_));
 sky130_fd_sc_hd__o21ai_1 _10556_ (.A1(_06076_),
    .A2(_06330_),
    .B1(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__mux2_8 _10557_ (.A0(net236),
    .A1(\ks1.key_reg[80] ),
    .S(_06097_),
    .X(_06336_));
 sky130_fd_sc_hd__xnor2_1 _10558_ (.A(_06335_),
    .B(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__mux2_1 _10559_ (.A0(\addroundkey_data_o[80] ),
    .A1(_06337_),
    .S(_06327_),
    .X(_06338_));
 sky130_fd_sc_hd__clkbuf_1 _10560_ (.A(_06338_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _10561_ (.A0(net108),
    .A1(\mix1.data_o[81] ),
    .S(_06111_),
    .X(_06339_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(\sub1.data_o[81] ),
    .A1(_06339_),
    .S(_06113_),
    .X(_06340_));
 sky130_fd_sc_hd__clkbuf_4 _10563_ (.A(_05613_),
    .X(_06341_));
 sky130_fd_sc_hd__clkbuf_4 _10564_ (.A(\sub1.ready_o ),
    .X(_06342_));
 sky130_fd_sc_hd__a31o_1 _10565_ (.A1(_06090_),
    .A2(_06342_),
    .A3(\sub1.data_o[81] ),
    .B1(_06079_),
    .X(_06343_));
 sky130_fd_sc_hd__a21o_1 _10566_ (.A1(_06126_),
    .A2(_06340_),
    .B1(_06343_),
    .X(_06344_));
 sky130_fd_sc_hd__o21a_1 _10567_ (.A1(\mix1.data_o[81] ),
    .A2(_06129_),
    .B1(_06093_),
    .X(_06345_));
 sky130_fd_sc_hd__a221o_1 _10568_ (.A1(\sub1.data_o[81] ),
    .A2(_06341_),
    .B1(_06344_),
    .B2(_06345_),
    .C1(_06118_),
    .X(_06346_));
 sky130_fd_sc_hd__o21ai_1 _10569_ (.A1(_06076_),
    .A2(_06340_),
    .B1(_06346_),
    .Y(_06347_));
 sky130_fd_sc_hd__mux2_4 _10570_ (.A0(net237),
    .A1(\ks1.key_reg[81] ),
    .S(_06097_),
    .X(_06348_));
 sky130_fd_sc_hd__xnor2_1 _10571_ (.A(_06347_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__mux2_1 _10572_ (.A0(\addroundkey_data_o[81] ),
    .A1(_06349_),
    .S(_06327_),
    .X(_06350_));
 sky130_fd_sc_hd__clkbuf_1 _10573_ (.A(_06350_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _10574_ (.A0(net109),
    .A1(\mix1.data_o[82] ),
    .S(_06111_),
    .X(_06351_));
 sky130_fd_sc_hd__mux2_1 _10575_ (.A0(\sub1.data_o[82] ),
    .A1(_06351_),
    .S(_06113_),
    .X(_06352_));
 sky130_fd_sc_hd__a31o_1 _10576_ (.A1(_06090_),
    .A2(_06342_),
    .A3(\sub1.data_o[82] ),
    .B1(_06079_),
    .X(_06353_));
 sky130_fd_sc_hd__a21o_1 _10577_ (.A1(_06126_),
    .A2(_06352_),
    .B1(_06353_),
    .X(_06354_));
 sky130_fd_sc_hd__o21a_1 _10578_ (.A1(\mix1.data_o[82] ),
    .A2(_06129_),
    .B1(_06093_),
    .X(_06355_));
 sky130_fd_sc_hd__a221o_1 _10579_ (.A1(\sub1.data_o[82] ),
    .A2(_06341_),
    .B1(_06354_),
    .B2(_06355_),
    .C1(_06118_),
    .X(_06356_));
 sky130_fd_sc_hd__o21ai_1 _10580_ (.A1(_06076_),
    .A2(_06352_),
    .B1(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__mux2_4 _10581_ (.A0(net238),
    .A1(\ks1.key_reg[82] ),
    .S(_06097_),
    .X(_06358_));
 sky130_fd_sc_hd__xnor2_1 _10582_ (.A(_06357_),
    .B(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(\addroundkey_data_o[82] ),
    .A1(_06359_),
    .S(_06327_),
    .X(_06360_));
 sky130_fd_sc_hd__clkbuf_1 _10584_ (.A(_06360_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(net110),
    .A1(\mix1.data_o[83] ),
    .S(_06111_),
    .X(_06361_));
 sky130_fd_sc_hd__mux2_1 _10586_ (.A0(\sub1.data_o[83] ),
    .A1(_06361_),
    .S(_06113_),
    .X(_06362_));
 sky130_fd_sc_hd__a31o_1 _10587_ (.A1(_06090_),
    .A2(_06342_),
    .A3(\sub1.data_o[83] ),
    .B1(_06079_),
    .X(_06363_));
 sky130_fd_sc_hd__a21o_1 _10588_ (.A1(_06126_),
    .A2(_06362_),
    .B1(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__o21a_1 _10589_ (.A1(\mix1.data_o[83] ),
    .A2(_06129_),
    .B1(_06093_),
    .X(_06365_));
 sky130_fd_sc_hd__a221o_1 _10590_ (.A1(\sub1.data_o[83] ),
    .A2(_06341_),
    .B1(_06364_),
    .B2(_06365_),
    .C1(_06118_),
    .X(_06366_));
 sky130_fd_sc_hd__o21ai_1 _10591_ (.A1(_06076_),
    .A2(_06362_),
    .B1(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__mux2_4 _10592_ (.A0(net239),
    .A1(\ks1.key_reg[83] ),
    .S(_06097_),
    .X(_06368_));
 sky130_fd_sc_hd__xnor2_1 _10593_ (.A(_06367_),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(\addroundkey_data_o[83] ),
    .A1(_06369_),
    .S(_06327_),
    .X(_06370_));
 sky130_fd_sc_hd__clkbuf_1 _10595_ (.A(_06370_),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _10596_ (.A0(net111),
    .A1(\mix1.data_o[84] ),
    .S(_06111_),
    .X(_06371_));
 sky130_fd_sc_hd__mux2_1 _10597_ (.A0(\sub1.data_o[84] ),
    .A1(_06371_),
    .S(_06113_),
    .X(_06372_));
 sky130_fd_sc_hd__a31o_1 _10598_ (.A1(_06090_),
    .A2(_06342_),
    .A3(\sub1.data_o[84] ),
    .B1(_06079_),
    .X(_06373_));
 sky130_fd_sc_hd__a21o_1 _10599_ (.A1(_06126_),
    .A2(_06372_),
    .B1(_06373_),
    .X(_06374_));
 sky130_fd_sc_hd__o21a_1 _10600_ (.A1(\mix1.data_o[84] ),
    .A2(_06129_),
    .B1(_06093_),
    .X(_06375_));
 sky130_fd_sc_hd__a221o_1 _10601_ (.A1(\sub1.data_o[84] ),
    .A2(_06341_),
    .B1(_06374_),
    .B2(_06375_),
    .C1(_06118_),
    .X(_06376_));
 sky130_fd_sc_hd__o21ai_4 _10602_ (.A1(_06076_),
    .A2(_06372_),
    .B1(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(net240),
    .A1(\ks1.key_reg[84] ),
    .S(_06097_),
    .X(_06378_));
 sky130_fd_sc_hd__xnor2_1 _10604_ (.A(_06377_),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__mux2_1 _10605_ (.A0(\addroundkey_data_o[84] ),
    .A1(_06379_),
    .S(_06327_),
    .X(_06380_));
 sky130_fd_sc_hd__clkbuf_1 _10606_ (.A(_06380_),
    .X(_00237_));
 sky130_fd_sc_hd__buf_8 _10607_ (.A(_05567_),
    .X(_06381_));
 sky130_fd_sc_hd__mux2_1 _10608_ (.A0(net112),
    .A1(\mix1.data_o[85] ),
    .S(_06111_),
    .X(_06382_));
 sky130_fd_sc_hd__mux2_1 _10609_ (.A0(\sub1.data_o[85] ),
    .A1(_06382_),
    .S(_06113_),
    .X(_06383_));
 sky130_fd_sc_hd__clkbuf_4 _10610_ (.A(_05584_),
    .X(_06384_));
 sky130_fd_sc_hd__a31o_1 _10611_ (.A1(_06090_),
    .A2(_06342_),
    .A3(\sub1.data_o[85] ),
    .B1(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__a21o_1 _10612_ (.A1(_06126_),
    .A2(_06383_),
    .B1(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__o21a_1 _10613_ (.A1(\mix1.data_o[85] ),
    .A2(_06129_),
    .B1(_06093_),
    .X(_06387_));
 sky130_fd_sc_hd__a221o_1 _10614_ (.A1(\sub1.data_o[85] ),
    .A2(_06341_),
    .B1(_06386_),
    .B2(_06387_),
    .C1(_06118_),
    .X(_06388_));
 sky130_fd_sc_hd__o21ai_1 _10615_ (.A1(_06381_),
    .A2(_06383_),
    .B1(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__mux2_4 _10616_ (.A0(net241),
    .A1(\ks1.key_reg[85] ),
    .S(_06097_),
    .X(_06390_));
 sky130_fd_sc_hd__xnor2_1 _10617_ (.A(_06389_),
    .B(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__mux2_1 _10618_ (.A0(\addroundkey_data_o[85] ),
    .A1(_06391_),
    .S(_06327_),
    .X(_06392_));
 sky130_fd_sc_hd__clkbuf_1 _10619_ (.A(_06392_),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(net113),
    .A1(\mix1.data_o[86] ),
    .S(_06111_),
    .X(_06393_));
 sky130_fd_sc_hd__mux2_1 _10621_ (.A0(\sub1.data_o[86] ),
    .A1(_06393_),
    .S(_06113_),
    .X(_06394_));
 sky130_fd_sc_hd__clkbuf_4 _10622_ (.A(_04624_),
    .X(_06395_));
 sky130_fd_sc_hd__a31o_1 _10623_ (.A1(_06395_),
    .A2(_06342_),
    .A3(\sub1.data_o[86] ),
    .B1(_06384_),
    .X(_06396_));
 sky130_fd_sc_hd__a21o_1 _10624_ (.A1(_06126_),
    .A2(_06394_),
    .B1(_06396_),
    .X(_06397_));
 sky130_fd_sc_hd__clkbuf_4 _10625_ (.A(_05757_),
    .X(_06398_));
 sky130_fd_sc_hd__o21a_1 _10626_ (.A1(\mix1.data_o[86] ),
    .A2(_06129_),
    .B1(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__a221o_1 _10627_ (.A1(\sub1.data_o[86] ),
    .A2(_06341_),
    .B1(_06397_),
    .B2(_06399_),
    .C1(_06118_),
    .X(_06400_));
 sky130_fd_sc_hd__o21ai_4 _10628_ (.A1(_06381_),
    .A2(_06394_),
    .B1(_06400_),
    .Y(_06401_));
 sky130_fd_sc_hd__clkbuf_8 _10629_ (.A(_04638_),
    .X(_06402_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(net242),
    .A1(\ks1.key_reg[86] ),
    .S(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__xnor2_1 _10631_ (.A(_06401_),
    .B(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(\addroundkey_data_o[86] ),
    .A1(_06404_),
    .S(_06327_),
    .X(_06405_));
 sky130_fd_sc_hd__clkbuf_1 _10633_ (.A(_06405_),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(net114),
    .A1(\mix1.data_o[87] ),
    .S(_06111_),
    .X(_06406_));
 sky130_fd_sc_hd__mux2_1 _10635_ (.A0(\sub1.data_o[87] ),
    .A1(_06406_),
    .S(_06113_),
    .X(_06407_));
 sky130_fd_sc_hd__a31o_1 _10636_ (.A1(_06395_),
    .A2(_06342_),
    .A3(\sub1.data_o[87] ),
    .B1(_06384_),
    .X(_06408_));
 sky130_fd_sc_hd__a21o_1 _10637_ (.A1(_06126_),
    .A2(_06407_),
    .B1(_06408_),
    .X(_06409_));
 sky130_fd_sc_hd__o21a_1 _10638_ (.A1(\mix1.data_o[87] ),
    .A2(_06129_),
    .B1(_06398_),
    .X(_06410_));
 sky130_fd_sc_hd__a221o_1 _10639_ (.A1(\sub1.data_o[87] ),
    .A2(_06341_),
    .B1(_06409_),
    .B2(_06410_),
    .C1(_06118_),
    .X(_06411_));
 sky130_fd_sc_hd__o21ai_1 _10640_ (.A1(_06381_),
    .A2(_06407_),
    .B1(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__mux2_8 _10641_ (.A0(net243),
    .A1(\ks1.key_reg[87] ),
    .S(_06402_),
    .X(_06413_));
 sky130_fd_sc_hd__xnor2_1 _10642_ (.A(_06412_),
    .B(_06413_),
    .Y(_06414_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(\addroundkey_data_o[87] ),
    .A1(_06414_),
    .S(_06327_),
    .X(_06415_));
 sky130_fd_sc_hd__clkbuf_1 _10644_ (.A(_06415_),
    .X(_00240_));
 sky130_fd_sc_hd__clkbuf_4 _10645_ (.A(_05614_),
    .X(_06416_));
 sky130_fd_sc_hd__mux2_1 _10646_ (.A0(net115),
    .A1(\mix1.data_o[88] ),
    .S(_06316_),
    .X(_06417_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(\sub1.data_o[88] ),
    .A1(_06417_),
    .S(_06318_),
    .X(_06418_));
 sky130_fd_sc_hd__a32o_1 _10648_ (.A1(\mix1.data_o[88] ),
    .A2(_06296_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[88] ),
    .X(_06419_));
 sky130_fd_sc_hd__clkbuf_4 _10649_ (.A(_04609_),
    .X(_06420_));
 sky130_fd_sc_hd__a22o_1 _10650_ (.A1(_06416_),
    .A2(_06418_),
    .B1(_06419_),
    .B2(_06420_),
    .X(_06421_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(net244),
    .A1(\ks1.key_reg[88] ),
    .S(_06324_),
    .X(_06422_));
 sky130_fd_sc_hd__xor2_1 _10652_ (.A(_06421_),
    .B(_06422_),
    .X(_06423_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(\addroundkey_data_o[88] ),
    .A1(_06423_),
    .S(_06327_),
    .X(_06424_));
 sky130_fd_sc_hd__clkbuf_1 _10654_ (.A(_06424_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(net116),
    .A1(\mix1.data_o[89] ),
    .S(_06316_),
    .X(_06425_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(\sub1.data_o[89] ),
    .A1(_06425_),
    .S(_06318_),
    .X(_06426_));
 sky130_fd_sc_hd__a32o_1 _10657_ (.A1(\mix1.data_o[89] ),
    .A2(_06296_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[89] ),
    .X(_06427_));
 sky130_fd_sc_hd__a22o_2 _10658_ (.A1(_06416_),
    .A2(_06426_),
    .B1(_06427_),
    .B2(_06420_),
    .X(_06428_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(net245),
    .A1(\ks1.key_reg[89] ),
    .S(_06324_),
    .X(_06429_));
 sky130_fd_sc_hd__xor2_1 _10660_ (.A(_06428_),
    .B(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__buf_4 _10661_ (.A(_05792_),
    .X(_06431_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(\addroundkey_data_o[89] ),
    .A1(_06430_),
    .S(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__clkbuf_1 _10663_ (.A(_06432_),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(net118),
    .A1(\mix1.data_o[90] ),
    .S(_06316_),
    .X(_06433_));
 sky130_fd_sc_hd__mux2_1 _10665_ (.A0(\sub1.data_o[90] ),
    .A1(_06433_),
    .S(_06318_),
    .X(_06434_));
 sky130_fd_sc_hd__a32o_1 _10666_ (.A1(\mix1.data_o[90] ),
    .A2(_06296_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[90] ),
    .X(_06435_));
 sky130_fd_sc_hd__a22o_1 _10667_ (.A1(_06416_),
    .A2(_06434_),
    .B1(_06435_),
    .B2(_06420_),
    .X(_06436_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(net247),
    .A1(\ks1.key_reg[90] ),
    .S(_06324_),
    .X(_06437_));
 sky130_fd_sc_hd__xor2_1 _10669_ (.A(_06436_),
    .B(_06437_),
    .X(_06438_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\addroundkey_data_o[90] ),
    .A1(_06438_),
    .S(_06431_),
    .X(_06439_));
 sky130_fd_sc_hd__clkbuf_1 _10671_ (.A(_06439_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(net119),
    .A1(\mix1.data_o[91] ),
    .S(_06316_),
    .X(_06440_));
 sky130_fd_sc_hd__mux2_1 _10673_ (.A0(\sub1.data_o[91] ),
    .A1(_06440_),
    .S(_06318_),
    .X(_06441_));
 sky130_fd_sc_hd__a32o_1 _10674_ (.A1(\mix1.data_o[91] ),
    .A2(_06296_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[91] ),
    .X(_06442_));
 sky130_fd_sc_hd__a22o_1 _10675_ (.A1(_06416_),
    .A2(_06441_),
    .B1(_06442_),
    .B2(_06420_),
    .X(_06443_));
 sky130_fd_sc_hd__mux2_1 _10676_ (.A0(net248),
    .A1(\ks1.key_reg[91] ),
    .S(_06324_),
    .X(_06444_));
 sky130_fd_sc_hd__xor2_1 _10677_ (.A(_06443_),
    .B(_06444_),
    .X(_06445_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(\addroundkey_data_o[91] ),
    .A1(_06445_),
    .S(_06431_),
    .X(_06446_));
 sky130_fd_sc_hd__clkbuf_1 _10679_ (.A(_06446_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(net120),
    .A1(\mix1.data_o[92] ),
    .S(_06316_),
    .X(_06447_));
 sky130_fd_sc_hd__mux2_1 _10681_ (.A0(\sub1.data_o[92] ),
    .A1(_06447_),
    .S(_06318_),
    .X(_06448_));
 sky130_fd_sc_hd__a32o_1 _10682_ (.A1(\mix1.data_o[92] ),
    .A2(_06296_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[92] ),
    .X(_06449_));
 sky130_fd_sc_hd__a22o_1 _10683_ (.A1(_06416_),
    .A2(_06448_),
    .B1(_06449_),
    .B2(_06420_),
    .X(_06450_));
 sky130_fd_sc_hd__mux2_1 _10684_ (.A0(net249),
    .A1(\ks1.key_reg[92] ),
    .S(_06324_),
    .X(_06451_));
 sky130_fd_sc_hd__xor2_1 _10685_ (.A(_06450_),
    .B(_06451_),
    .X(_06452_));
 sky130_fd_sc_hd__mux2_1 _10686_ (.A0(\addroundkey_data_o[92] ),
    .A1(_06452_),
    .S(_06431_),
    .X(_06453_));
 sky130_fd_sc_hd__clkbuf_1 _10687_ (.A(_06453_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _10688_ (.A0(net121),
    .A1(\mix1.data_o[93] ),
    .S(_06316_),
    .X(_06454_));
 sky130_fd_sc_hd__mux2_1 _10689_ (.A0(\sub1.data_o[93] ),
    .A1(_06454_),
    .S(_06318_),
    .X(_06455_));
 sky130_fd_sc_hd__a32o_1 _10690_ (.A1(\mix1.data_o[93] ),
    .A2(_06296_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[93] ),
    .X(_06456_));
 sky130_fd_sc_hd__a22o_1 _10691_ (.A1(_06416_),
    .A2(_06455_),
    .B1(_06456_),
    .B2(_06420_),
    .X(_06457_));
 sky130_fd_sc_hd__mux2_1 _10692_ (.A0(net250),
    .A1(\ks1.key_reg[93] ),
    .S(_06324_),
    .X(_06458_));
 sky130_fd_sc_hd__xor2_1 _10693_ (.A(_06457_),
    .B(_06458_),
    .X(_06459_));
 sky130_fd_sc_hd__mux2_1 _10694_ (.A0(\addroundkey_data_o[93] ),
    .A1(_06459_),
    .S(_06431_),
    .X(_06460_));
 sky130_fd_sc_hd__clkbuf_1 _10695_ (.A(_06460_),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _10696_ (.A0(net122),
    .A1(\mix1.data_o[94] ),
    .S(_06316_),
    .X(_06461_));
 sky130_fd_sc_hd__mux2_1 _10697_ (.A0(\sub1.data_o[94] ),
    .A1(_06461_),
    .S(_06318_),
    .X(_06462_));
 sky130_fd_sc_hd__clkbuf_4 _10698_ (.A(_05585_),
    .X(_06463_));
 sky130_fd_sc_hd__a32o_1 _10699_ (.A1(\mix1.data_o[94] ),
    .A2(_06463_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[94] ),
    .X(_06464_));
 sky130_fd_sc_hd__a22o_1 _10700_ (.A1(_06416_),
    .A2(_06462_),
    .B1(_06464_),
    .B2(_06420_),
    .X(_06465_));
 sky130_fd_sc_hd__mux2_1 _10701_ (.A0(net251),
    .A1(\ks1.key_reg[94] ),
    .S(_06324_),
    .X(_06466_));
 sky130_fd_sc_hd__xor2_1 _10702_ (.A(_06465_),
    .B(_06466_),
    .X(_06467_));
 sky130_fd_sc_hd__mux2_1 _10703_ (.A0(\addroundkey_data_o[94] ),
    .A1(_06467_),
    .S(_06431_),
    .X(_06468_));
 sky130_fd_sc_hd__clkbuf_1 _10704_ (.A(_06468_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _10705_ (.A0(net123),
    .A1(\mix1.data_o[95] ),
    .S(_06316_),
    .X(_06469_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(\sub1.data_o[95] ),
    .A1(_06469_),
    .S(_06318_),
    .X(_06470_));
 sky130_fd_sc_hd__a32o_1 _10707_ (.A1(\mix1.data_o[95] ),
    .A2(_06463_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[95] ),
    .X(_06471_));
 sky130_fd_sc_hd__a22o_2 _10708_ (.A1(_06416_),
    .A2(_06470_),
    .B1(_06471_),
    .B2(_06420_),
    .X(_06472_));
 sky130_fd_sc_hd__mux2_1 _10709_ (.A0(net252),
    .A1(\ks1.key_reg[95] ),
    .S(_06324_),
    .X(_06473_));
 sky130_fd_sc_hd__xor2_1 _10710_ (.A(_06472_),
    .B(_06473_),
    .X(_06474_));
 sky130_fd_sc_hd__mux2_1 _10711_ (.A0(\addroundkey_data_o[95] ),
    .A1(_06474_),
    .S(_06431_),
    .X(_06475_));
 sky130_fd_sc_hd__clkbuf_1 _10712_ (.A(_06475_),
    .X(_00248_));
 sky130_fd_sc_hd__buf_4 _10713_ (.A(_05602_),
    .X(_06476_));
 sky130_fd_sc_hd__mux2_1 _10714_ (.A0(net124),
    .A1(\mix1.data_o[96] ),
    .S(_06476_),
    .X(_06477_));
 sky130_fd_sc_hd__buf_4 _10715_ (.A(_05608_),
    .X(_06478_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(\sub1.data_o[96] ),
    .A1(_06477_),
    .S(_06478_),
    .X(_06479_));
 sky130_fd_sc_hd__a31o_1 _10717_ (.A1(_06395_),
    .A2(_06342_),
    .A3(\sub1.data_o[96] ),
    .B1(_06384_),
    .X(_06480_));
 sky130_fd_sc_hd__a21o_1 _10718_ (.A1(_06126_),
    .A2(_06479_),
    .B1(_06480_),
    .X(_06481_));
 sky130_fd_sc_hd__o21a_1 _10719_ (.A1(\mix1.data_o[96] ),
    .A2(_06129_),
    .B1(_06398_),
    .X(_06482_));
 sky130_fd_sc_hd__clkbuf_4 _10720_ (.A(_04610_),
    .X(_06483_));
 sky130_fd_sc_hd__a221o_1 _10721_ (.A1(\sub1.data_o[96] ),
    .A2(_06341_),
    .B1(_06481_),
    .B2(_06482_),
    .C1(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__o21ai_4 _10722_ (.A1(_06381_),
    .A2(_06479_),
    .B1(_06484_),
    .Y(_06485_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(net253),
    .A1(\ks1.key_reg[96] ),
    .S(_06402_),
    .X(_06486_));
 sky130_fd_sc_hd__xnor2_1 _10724_ (.A(_06485_),
    .B(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(\addroundkey_data_o[96] ),
    .A1(_06487_),
    .S(_06431_),
    .X(_06488_));
 sky130_fd_sc_hd__clkbuf_1 _10726_ (.A(_06488_),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(net125),
    .A1(\mix1.data_o[97] ),
    .S(_06476_),
    .X(_06489_));
 sky130_fd_sc_hd__mux2_1 _10728_ (.A0(\sub1.data_o[97] ),
    .A1(_06489_),
    .S(_06478_),
    .X(_06490_));
 sky130_fd_sc_hd__clkbuf_4 _10729_ (.A(_05574_),
    .X(_06491_));
 sky130_fd_sc_hd__a31o_1 _10730_ (.A1(_06395_),
    .A2(_06342_),
    .A3(\sub1.data_o[97] ),
    .B1(_06384_),
    .X(_06492_));
 sky130_fd_sc_hd__a21o_1 _10731_ (.A1(_06491_),
    .A2(_06490_),
    .B1(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__clkbuf_4 _10732_ (.A(_04626_),
    .X(_06494_));
 sky130_fd_sc_hd__o21a_1 _10733_ (.A1(\mix1.data_o[97] ),
    .A2(_06494_),
    .B1(_06398_),
    .X(_06495_));
 sky130_fd_sc_hd__a221o_1 _10734_ (.A1(\sub1.data_o[97] ),
    .A2(_06341_),
    .B1(_06493_),
    .B2(_06495_),
    .C1(_06483_),
    .X(_06496_));
 sky130_fd_sc_hd__o21ai_4 _10735_ (.A1(_06381_),
    .A2(_06490_),
    .B1(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(net254),
    .A1(\ks1.key_reg[97] ),
    .S(_06402_),
    .X(_06498_));
 sky130_fd_sc_hd__xnor2_1 _10737_ (.A(_06497_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(\addroundkey_data_o[97] ),
    .A1(_06499_),
    .S(_06431_),
    .X(_06500_));
 sky130_fd_sc_hd__clkbuf_1 _10739_ (.A(_06500_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _10740_ (.A0(net126),
    .A1(\mix1.data_o[98] ),
    .S(_06476_),
    .X(_06501_));
 sky130_fd_sc_hd__mux2_1 _10741_ (.A0(\sub1.data_o[98] ),
    .A1(_06501_),
    .S(_06478_),
    .X(_06502_));
 sky130_fd_sc_hd__a31o_1 _10742_ (.A1(_06395_),
    .A2(_06342_),
    .A3(\sub1.data_o[98] ),
    .B1(_06384_),
    .X(_06503_));
 sky130_fd_sc_hd__a21o_1 _10743_ (.A1(_06491_),
    .A2(_06502_),
    .B1(_06503_),
    .X(_06504_));
 sky130_fd_sc_hd__o21a_1 _10744_ (.A1(\mix1.data_o[98] ),
    .A2(_06494_),
    .B1(_06398_),
    .X(_06505_));
 sky130_fd_sc_hd__a221o_1 _10745_ (.A1(\sub1.data_o[98] ),
    .A2(_06341_),
    .B1(_06504_),
    .B2(_06505_),
    .C1(_06483_),
    .X(_06506_));
 sky130_fd_sc_hd__o21ai_4 _10746_ (.A1(_06381_),
    .A2(_06502_),
    .B1(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__mux2_1 _10747_ (.A0(net255),
    .A1(\ks1.key_reg[98] ),
    .S(_06402_),
    .X(_06508_));
 sky130_fd_sc_hd__xnor2_1 _10748_ (.A(_06507_),
    .B(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__mux2_1 _10749_ (.A0(\addroundkey_data_o[98] ),
    .A1(_06509_),
    .S(_06431_),
    .X(_06510_));
 sky130_fd_sc_hd__clkbuf_1 _10750_ (.A(_06510_),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _10751_ (.A0(net127),
    .A1(\mix1.data_o[99] ),
    .S(_06476_),
    .X(_06511_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(\sub1.data_o[99] ),
    .A1(_06511_),
    .S(_06478_),
    .X(_06512_));
 sky130_fd_sc_hd__clkbuf_4 _10753_ (.A(_05613_),
    .X(_06513_));
 sky130_fd_sc_hd__clkbuf_4 _10754_ (.A(\sub1.ready_o ),
    .X(_06514_));
 sky130_fd_sc_hd__a31o_1 _10755_ (.A1(_06395_),
    .A2(_06514_),
    .A3(\sub1.data_o[99] ),
    .B1(_06384_),
    .X(_06515_));
 sky130_fd_sc_hd__a21o_1 _10756_ (.A1(_06491_),
    .A2(_06512_),
    .B1(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__o21a_1 _10757_ (.A1(\mix1.data_o[99] ),
    .A2(_06494_),
    .B1(_06398_),
    .X(_06517_));
 sky130_fd_sc_hd__a221o_1 _10758_ (.A1(\sub1.data_o[99] ),
    .A2(_06513_),
    .B1(_06516_),
    .B2(_06517_),
    .C1(_06483_),
    .X(_06518_));
 sky130_fd_sc_hd__o21ai_4 _10759_ (.A1(_06381_),
    .A2(_06512_),
    .B1(_06518_),
    .Y(_06519_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(net256),
    .A1(\ks1.key_reg[99] ),
    .S(_06402_),
    .X(_06520_));
 sky130_fd_sc_hd__xnor2_1 _10761_ (.A(_06519_),
    .B(_06520_),
    .Y(_06521_));
 sky130_fd_sc_hd__buf_4 _10762_ (.A(_05792_),
    .X(_06522_));
 sky130_fd_sc_hd__mux2_1 _10763_ (.A0(\addroundkey_data_o[99] ),
    .A1(_06521_),
    .S(_06522_),
    .X(_06523_));
 sky130_fd_sc_hd__clkbuf_1 _10764_ (.A(_06523_),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _10765_ (.A0(net2),
    .A1(\mix1.data_o[100] ),
    .S(_06476_),
    .X(_06524_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(\sub1.data_o[100] ),
    .A1(_06524_),
    .S(_06478_),
    .X(_06525_));
 sky130_fd_sc_hd__a31o_1 _10767_ (.A1(_06395_),
    .A2(_06514_),
    .A3(\sub1.data_o[100] ),
    .B1(_06384_),
    .X(_06526_));
 sky130_fd_sc_hd__a21o_1 _10768_ (.A1(_06491_),
    .A2(_06525_),
    .B1(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__o21a_1 _10769_ (.A1(\mix1.data_o[100] ),
    .A2(_06494_),
    .B1(_06398_),
    .X(_06528_));
 sky130_fd_sc_hd__a221o_1 _10770_ (.A1(\sub1.data_o[100] ),
    .A2(_06513_),
    .B1(_06527_),
    .B2(_06528_),
    .C1(_06483_),
    .X(_06529_));
 sky130_fd_sc_hd__o21ai_4 _10771_ (.A1(_06381_),
    .A2(_06525_),
    .B1(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(net131),
    .A1(\ks1.key_reg[100] ),
    .S(_06402_),
    .X(_06531_));
 sky130_fd_sc_hd__xnor2_1 _10773_ (.A(_06530_),
    .B(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(\addroundkey_data_o[100] ),
    .A1(_06532_),
    .S(_06522_),
    .X(_06533_));
 sky130_fd_sc_hd__clkbuf_1 _10775_ (.A(_06533_),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(net3),
    .A1(\mix1.data_o[101] ),
    .S(_06476_),
    .X(_06534_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(\sub1.data_o[101] ),
    .A1(_06534_),
    .S(_06478_),
    .X(_06535_));
 sky130_fd_sc_hd__a31o_1 _10778_ (.A1(_06395_),
    .A2(_06514_),
    .A3(\sub1.data_o[101] ),
    .B1(_06384_),
    .X(_06536_));
 sky130_fd_sc_hd__a21o_1 _10779_ (.A1(_06491_),
    .A2(_06535_),
    .B1(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__o21a_1 _10780_ (.A1(\mix1.data_o[101] ),
    .A2(_06494_),
    .B1(_06398_),
    .X(_06538_));
 sky130_fd_sc_hd__a221o_1 _10781_ (.A1(\sub1.data_o[101] ),
    .A2(_06513_),
    .B1(_06537_),
    .B2(_06538_),
    .C1(_06483_),
    .X(_06539_));
 sky130_fd_sc_hd__o21ai_2 _10782_ (.A1(_06381_),
    .A2(_06535_),
    .B1(_06539_),
    .Y(_06540_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(net132),
    .A1(\ks1.key_reg[101] ),
    .S(_06402_),
    .X(_06541_));
 sky130_fd_sc_hd__xnor2_1 _10784_ (.A(_06540_),
    .B(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(\addroundkey_data_o[101] ),
    .A1(_06542_),
    .S(_06522_),
    .X(_06543_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(_06543_),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(net4),
    .A1(\mix1.data_o[102] ),
    .S(_06476_),
    .X(_06544_));
 sky130_fd_sc_hd__mux2_1 _10788_ (.A0(\sub1.data_o[102] ),
    .A1(_06544_),
    .S(_06478_),
    .X(_06545_));
 sky130_fd_sc_hd__a31o_1 _10789_ (.A1(_06395_),
    .A2(_06514_),
    .A3(\sub1.data_o[102] ),
    .B1(_06384_),
    .X(_06546_));
 sky130_fd_sc_hd__a21o_1 _10790_ (.A1(_06491_),
    .A2(_06545_),
    .B1(_06546_),
    .X(_06547_));
 sky130_fd_sc_hd__o21a_1 _10791_ (.A1(\mix1.data_o[102] ),
    .A2(_06494_),
    .B1(_06398_),
    .X(_06548_));
 sky130_fd_sc_hd__a221o_1 _10792_ (.A1(\sub1.data_o[102] ),
    .A2(_06513_),
    .B1(_06547_),
    .B2(_06548_),
    .C1(_06483_),
    .X(_06549_));
 sky130_fd_sc_hd__o21ai_2 _10793_ (.A1(_06381_),
    .A2(_06545_),
    .B1(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__mux2_1 _10794_ (.A0(net133),
    .A1(\ks1.key_reg[102] ),
    .S(_06402_),
    .X(_06551_));
 sky130_fd_sc_hd__xnor2_1 _10795_ (.A(_06550_),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__mux2_1 _10796_ (.A0(\addroundkey_data_o[102] ),
    .A1(_06552_),
    .S(_06522_),
    .X(_06553_));
 sky130_fd_sc_hd__clkbuf_1 _10797_ (.A(_06553_),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _10798_ (.A0(net5),
    .A1(\mix1.data_o[103] ),
    .S(_06476_),
    .X(_06554_));
 sky130_fd_sc_hd__mux2_1 _10799_ (.A0(\sub1.data_o[103] ),
    .A1(_06554_),
    .S(_06478_),
    .X(_06555_));
 sky130_fd_sc_hd__a31o_1 _10800_ (.A1(_06395_),
    .A2(_06514_),
    .A3(\sub1.data_o[103] ),
    .B1(_05675_),
    .X(_06556_));
 sky130_fd_sc_hd__a21o_1 _10801_ (.A1(_06491_),
    .A2(_06555_),
    .B1(_06556_),
    .X(_06557_));
 sky130_fd_sc_hd__o21a_1 _10802_ (.A1(\mix1.data_o[103] ),
    .A2(_06494_),
    .B1(_06398_),
    .X(_06558_));
 sky130_fd_sc_hd__a221o_1 _10803_ (.A1(\sub1.data_o[103] ),
    .A2(_06513_),
    .B1(_06557_),
    .B2(_06558_),
    .C1(_06483_),
    .X(_06559_));
 sky130_fd_sc_hd__o21ai_4 _10804_ (.A1(_05623_),
    .A2(_06555_),
    .B1(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__mux2_1 _10805_ (.A0(net134),
    .A1(\ks1.key_reg[103] ),
    .S(_06402_),
    .X(_06561_));
 sky130_fd_sc_hd__xnor2_1 _10806_ (.A(_06560_),
    .B(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(\addroundkey_data_o[103] ),
    .A1(_06562_),
    .S(_06522_),
    .X(_06563_));
 sky130_fd_sc_hd__clkbuf_1 _10808_ (.A(_06563_),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _10809_ (.A0(net6),
    .A1(\mix1.data_o[104] ),
    .S(_06316_),
    .X(_06564_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(\sub1.data_o[104] ),
    .A1(_06564_),
    .S(_06318_),
    .X(_06565_));
 sky130_fd_sc_hd__a32o_1 _10811_ (.A1(\mix1.data_o[104] ),
    .A2(_06463_),
    .A3(_06320_),
    .B1(_06321_),
    .B2(\sub1.data_o[104] ),
    .X(_06566_));
 sky130_fd_sc_hd__a22o_1 _10812_ (.A1(_06416_),
    .A2(_06565_),
    .B1(_06566_),
    .B2(_06420_),
    .X(_06567_));
 sky130_fd_sc_hd__mux2_1 _10813_ (.A0(net135),
    .A1(\ks1.key_reg[104] ),
    .S(_06324_),
    .X(_06568_));
 sky130_fd_sc_hd__xor2_1 _10814_ (.A(_06567_),
    .B(_06568_),
    .X(_06569_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(\addroundkey_data_o[104] ),
    .A1(_06569_),
    .S(_06522_),
    .X(_06570_));
 sky130_fd_sc_hd__clkbuf_1 _10816_ (.A(_06570_),
    .X(_00257_));
 sky130_fd_sc_hd__buf_4 _10817_ (.A(_05749_),
    .X(_06571_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(net7),
    .A1(\mix1.data_o[105] ),
    .S(_06571_),
    .X(_06572_));
 sky130_fd_sc_hd__buf_4 _10819_ (.A(_05751_),
    .X(_06573_));
 sky130_fd_sc_hd__mux2_1 _10820_ (.A0(\sub1.data_o[105] ),
    .A1(_06572_),
    .S(_06573_),
    .X(_06574_));
 sky130_fd_sc_hd__clkbuf_4 _10821_ (.A(_05757_),
    .X(_06575_));
 sky130_fd_sc_hd__clkbuf_4 _10822_ (.A(_05619_),
    .X(_06576_));
 sky130_fd_sc_hd__a32o_1 _10823_ (.A1(\mix1.data_o[105] ),
    .A2(_06463_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[105] ),
    .X(_06577_));
 sky130_fd_sc_hd__a22o_1 _10824_ (.A1(_06416_),
    .A2(_06574_),
    .B1(_06577_),
    .B2(_06420_),
    .X(_06578_));
 sky130_fd_sc_hd__buf_4 _10825_ (.A(_05707_),
    .X(_06579_));
 sky130_fd_sc_hd__mux2_1 _10826_ (.A0(net136),
    .A1(\ks1.key_reg[105] ),
    .S(_06579_),
    .X(_06580_));
 sky130_fd_sc_hd__xor2_1 _10827_ (.A(_06578_),
    .B(_06580_),
    .X(_06581_));
 sky130_fd_sc_hd__mux2_1 _10828_ (.A0(\addroundkey_data_o[105] ),
    .A1(_06581_),
    .S(_06522_),
    .X(_06582_));
 sky130_fd_sc_hd__clkbuf_1 _10829_ (.A(_06582_),
    .X(_00258_));
 sky130_fd_sc_hd__clkbuf_4 _10830_ (.A(_05614_),
    .X(_06583_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(net8),
    .A1(\mix1.data_o[106] ),
    .S(_06571_),
    .X(_06584_));
 sky130_fd_sc_hd__mux2_1 _10832_ (.A0(\sub1.data_o[106] ),
    .A1(_06584_),
    .S(_06573_),
    .X(_06585_));
 sky130_fd_sc_hd__a32o_1 _10833_ (.A1(\mix1.data_o[106] ),
    .A2(_06463_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[106] ),
    .X(_06586_));
 sky130_fd_sc_hd__clkbuf_4 _10834_ (.A(_04609_),
    .X(_06587_));
 sky130_fd_sc_hd__a22o_1 _10835_ (.A1(_06583_),
    .A2(_06585_),
    .B1(_06586_),
    .B2(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__mux2_1 _10836_ (.A0(net137),
    .A1(\ks1.key_reg[106] ),
    .S(_06579_),
    .X(_06589_));
 sky130_fd_sc_hd__xor2_1 _10837_ (.A(_06588_),
    .B(_06589_),
    .X(_06590_));
 sky130_fd_sc_hd__mux2_1 _10838_ (.A0(\addroundkey_data_o[106] ),
    .A1(_06590_),
    .S(_06522_),
    .X(_06591_));
 sky130_fd_sc_hd__clkbuf_1 _10839_ (.A(_06591_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _10840_ (.A0(net9),
    .A1(\mix1.data_o[107] ),
    .S(_06571_),
    .X(_06592_));
 sky130_fd_sc_hd__mux2_1 _10841_ (.A0(\sub1.data_o[107] ),
    .A1(_06592_),
    .S(_06573_),
    .X(_06593_));
 sky130_fd_sc_hd__a32o_1 _10842_ (.A1(\mix1.data_o[107] ),
    .A2(_06463_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[107] ),
    .X(_06594_));
 sky130_fd_sc_hd__a22o_1 _10843_ (.A1(_06583_),
    .A2(_06593_),
    .B1(_06594_),
    .B2(_06587_),
    .X(_06595_));
 sky130_fd_sc_hd__mux2_1 _10844_ (.A0(net138),
    .A1(\ks1.key_reg[107] ),
    .S(_06579_),
    .X(_06596_));
 sky130_fd_sc_hd__xor2_1 _10845_ (.A(_06595_),
    .B(_06596_),
    .X(_06597_));
 sky130_fd_sc_hd__mux2_1 _10846_ (.A0(\addroundkey_data_o[107] ),
    .A1(_06597_),
    .S(_06522_),
    .X(_06598_));
 sky130_fd_sc_hd__clkbuf_1 _10847_ (.A(_06598_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _10848_ (.A0(net10),
    .A1(\mix1.data_o[108] ),
    .S(_06571_),
    .X(_06599_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(\sub1.data_o[108] ),
    .A1(_06599_),
    .S(_06573_),
    .X(_06600_));
 sky130_fd_sc_hd__a32o_1 _10850_ (.A1(\mix1.data_o[108] ),
    .A2(_06463_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[108] ),
    .X(_06601_));
 sky130_fd_sc_hd__a22o_1 _10851_ (.A1(_06583_),
    .A2(_06600_),
    .B1(_06601_),
    .B2(_06587_),
    .X(_06602_));
 sky130_fd_sc_hd__mux2_1 _10852_ (.A0(net139),
    .A1(\ks1.key_reg[108] ),
    .S(_06579_),
    .X(_06603_));
 sky130_fd_sc_hd__xor2_1 _10853_ (.A(_06602_),
    .B(_06603_),
    .X(_06604_));
 sky130_fd_sc_hd__mux2_1 _10854_ (.A0(\addroundkey_data_o[108] ),
    .A1(_06604_),
    .S(_06522_),
    .X(_06605_));
 sky130_fd_sc_hd__clkbuf_1 _10855_ (.A(_06605_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _10856_ (.A0(net11),
    .A1(\mix1.data_o[109] ),
    .S(_06571_),
    .X(_06606_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(\sub1.data_o[109] ),
    .A1(_06606_),
    .S(_06573_),
    .X(_06607_));
 sky130_fd_sc_hd__a32o_1 _10858_ (.A1(\mix1.data_o[109] ),
    .A2(_06463_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[109] ),
    .X(_06608_));
 sky130_fd_sc_hd__a22o_1 _10859_ (.A1(_06583_),
    .A2(_06607_),
    .B1(_06608_),
    .B2(_06587_),
    .X(_06609_));
 sky130_fd_sc_hd__mux2_1 _10860_ (.A0(net140),
    .A1(\ks1.key_reg[109] ),
    .S(_06579_),
    .X(_06610_));
 sky130_fd_sc_hd__xor2_1 _10861_ (.A(_06609_),
    .B(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__buf_4 _10862_ (.A(_05792_),
    .X(_06612_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(\addroundkey_data_o[109] ),
    .A1(_06611_),
    .S(_06612_),
    .X(_06613_));
 sky130_fd_sc_hd__clkbuf_1 _10864_ (.A(_06613_),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _10865_ (.A0(net13),
    .A1(\mix1.data_o[110] ),
    .S(_06571_),
    .X(_06614_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(\sub1.data_o[110] ),
    .A1(_06614_),
    .S(_06573_),
    .X(_06615_));
 sky130_fd_sc_hd__a32o_1 _10867_ (.A1(\mix1.data_o[110] ),
    .A2(_06463_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[110] ),
    .X(_06616_));
 sky130_fd_sc_hd__a22o_1 _10868_ (.A1(_06583_),
    .A2(_06615_),
    .B1(_06616_),
    .B2(_06587_),
    .X(_06617_));
 sky130_fd_sc_hd__mux2_1 _10869_ (.A0(net142),
    .A1(\ks1.key_reg[110] ),
    .S(_06579_),
    .X(_06618_));
 sky130_fd_sc_hd__xor2_1 _10870_ (.A(_06617_),
    .B(_06618_),
    .X(_06619_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(\addroundkey_data_o[110] ),
    .A1(_06619_),
    .S(_06612_),
    .X(_06620_));
 sky130_fd_sc_hd__clkbuf_1 _10872_ (.A(_06620_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _10873_ (.A0(net14),
    .A1(\mix1.data_o[111] ),
    .S(_06571_),
    .X(_06621_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(\sub1.data_o[111] ),
    .A1(_06621_),
    .S(_06573_),
    .X(_06622_));
 sky130_fd_sc_hd__a32o_1 _10875_ (.A1(\mix1.data_o[111] ),
    .A2(_06463_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[111] ),
    .X(_06623_));
 sky130_fd_sc_hd__a22o_1 _10876_ (.A1(_06583_),
    .A2(_06622_),
    .B1(_06623_),
    .B2(_06587_),
    .X(_06624_));
 sky130_fd_sc_hd__mux2_1 _10877_ (.A0(net143),
    .A1(\ks1.key_reg[111] ),
    .S(_06579_),
    .X(_06625_));
 sky130_fd_sc_hd__xor2_1 _10878_ (.A(_06624_),
    .B(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__mux2_1 _10879_ (.A0(\addroundkey_data_o[111] ),
    .A1(_06626_),
    .S(_06612_),
    .X(_06627_));
 sky130_fd_sc_hd__clkbuf_1 _10880_ (.A(_06627_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _10881_ (.A0(net15),
    .A1(\mix1.data_o[112] ),
    .S(_06476_),
    .X(_06628_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(\sub1.data_o[112] ),
    .A1(_06628_),
    .S(_06478_),
    .X(_06629_));
 sky130_fd_sc_hd__clkbuf_4 _10883_ (.A(_04624_),
    .X(_06630_));
 sky130_fd_sc_hd__a31o_1 _10884_ (.A1(_06630_),
    .A2(_06514_),
    .A3(\sub1.data_o[112] ),
    .B1(_05675_),
    .X(_06631_));
 sky130_fd_sc_hd__a21o_1 _10885_ (.A1(_06491_),
    .A2(_06629_),
    .B1(_06631_),
    .X(_06632_));
 sky130_fd_sc_hd__o21a_1 _10886_ (.A1(\mix1.data_o[112] ),
    .A2(_06494_),
    .B1(_05617_),
    .X(_06633_));
 sky130_fd_sc_hd__a221o_1 _10887_ (.A1(\sub1.data_o[112] ),
    .A2(_06513_),
    .B1(_06632_),
    .B2(_06633_),
    .C1(_06483_),
    .X(_06634_));
 sky130_fd_sc_hd__o21ai_4 _10888_ (.A1(_05623_),
    .A2(_06629_),
    .B1(_06634_),
    .Y(_06635_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(net144),
    .A1(\ks1.key_reg[112] ),
    .S(_04639_),
    .X(_06636_));
 sky130_fd_sc_hd__xnor2_1 _10890_ (.A(_06635_),
    .B(_06636_),
    .Y(_06637_));
 sky130_fd_sc_hd__mux2_1 _10891_ (.A0(\addroundkey_data_o[112] ),
    .A1(_06637_),
    .S(_06612_),
    .X(_06638_));
 sky130_fd_sc_hd__clkbuf_1 _10892_ (.A(_06638_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(net16),
    .A1(\mix1.data_o[113] ),
    .S(_06476_),
    .X(_06639_));
 sky130_fd_sc_hd__mux2_1 _10894_ (.A0(\sub1.data_o[113] ),
    .A1(_06639_),
    .S(_06478_),
    .X(_06640_));
 sky130_fd_sc_hd__a31o_1 _10895_ (.A1(_06630_),
    .A2(_06514_),
    .A3(\sub1.data_o[113] ),
    .B1(_05675_),
    .X(_06641_));
 sky130_fd_sc_hd__a21o_1 _10896_ (.A1(_06491_),
    .A2(_06640_),
    .B1(_06641_),
    .X(_06642_));
 sky130_fd_sc_hd__o21a_1 _10897_ (.A1(\mix1.data_o[113] ),
    .A2(_06494_),
    .B1(_05617_),
    .X(_06643_));
 sky130_fd_sc_hd__a221o_1 _10898_ (.A1(\sub1.data_o[113] ),
    .A2(_06513_),
    .B1(_06642_),
    .B2(_06643_),
    .C1(_06483_),
    .X(_06644_));
 sky130_fd_sc_hd__o21ai_4 _10899_ (.A1(_05623_),
    .A2(_06640_),
    .B1(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__mux2_1 _10900_ (.A0(net145),
    .A1(\ks1.key_reg[113] ),
    .S(_04639_),
    .X(_06646_));
 sky130_fd_sc_hd__xnor2_1 _10901_ (.A(_06645_),
    .B(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__mux2_1 _10902_ (.A0(\addroundkey_data_o[113] ),
    .A1(_06647_),
    .S(_06612_),
    .X(_06648_));
 sky130_fd_sc_hd__clkbuf_1 _10903_ (.A(_06648_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _10904_ (.A0(net17),
    .A1(\mix1.data_o[114] ),
    .S(_05602_),
    .X(_06649_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(\sub1.data_o[114] ),
    .A1(_06649_),
    .S(_05608_),
    .X(_06650_));
 sky130_fd_sc_hd__a31o_1 _10906_ (.A1(_06630_),
    .A2(_06514_),
    .A3(\sub1.data_o[114] ),
    .B1(_05675_),
    .X(_06651_));
 sky130_fd_sc_hd__a21o_1 _10907_ (.A1(_06491_),
    .A2(_06650_),
    .B1(_06651_),
    .X(_06652_));
 sky130_fd_sc_hd__o21a_1 _10908_ (.A1(\mix1.data_o[114] ),
    .A2(_06494_),
    .B1(_05617_),
    .X(_06653_));
 sky130_fd_sc_hd__a221o_1 _10909_ (.A1(\sub1.data_o[114] ),
    .A2(_06513_),
    .B1(_06652_),
    .B2(_06653_),
    .C1(_04610_),
    .X(_06654_));
 sky130_fd_sc_hd__o21ai_1 _10910_ (.A1(_05623_),
    .A2(_06650_),
    .B1(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__mux2_4 _10911_ (.A0(net146),
    .A1(\ks1.key_reg[114] ),
    .S(_04639_),
    .X(_06656_));
 sky130_fd_sc_hd__xnor2_1 _10912_ (.A(_06655_),
    .B(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(\addroundkey_data_o[114] ),
    .A1(_06657_),
    .S(_06612_),
    .X(_06658_));
 sky130_fd_sc_hd__clkbuf_1 _10914_ (.A(_06658_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _10915_ (.A0(net18),
    .A1(\mix1.data_o[115] ),
    .S(_05602_),
    .X(_06659_));
 sky130_fd_sc_hd__mux2_1 _10916_ (.A0(\sub1.data_o[115] ),
    .A1(_06659_),
    .S(_05608_),
    .X(_06660_));
 sky130_fd_sc_hd__a31o_1 _10917_ (.A1(_06630_),
    .A2(_06514_),
    .A3(\sub1.data_o[115] ),
    .B1(_05675_),
    .X(_06661_));
 sky130_fd_sc_hd__a21o_1 _10918_ (.A1(_05574_),
    .A2(_06660_),
    .B1(_06661_),
    .X(_06662_));
 sky130_fd_sc_hd__o21a_1 _10919_ (.A1(\mix1.data_o[115] ),
    .A2(_04626_),
    .B1(_05617_),
    .X(_06663_));
 sky130_fd_sc_hd__a221o_1 _10920_ (.A1(\sub1.data_o[115] ),
    .A2(_06513_),
    .B1(_06662_),
    .B2(_06663_),
    .C1(_04610_),
    .X(_06664_));
 sky130_fd_sc_hd__o21ai_1 _10921_ (.A1(_05623_),
    .A2(_06660_),
    .B1(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__mux2_2 _10922_ (.A0(net147),
    .A1(\ks1.key_reg[115] ),
    .S(_04639_),
    .X(_06666_));
 sky130_fd_sc_hd__xnor2_1 _10923_ (.A(_06665_),
    .B(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(\addroundkey_data_o[115] ),
    .A1(_06667_),
    .S(_06612_),
    .X(_06668_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(_06668_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(net19),
    .A1(\mix1.data_o[116] ),
    .S(_05602_),
    .X(_06669_));
 sky130_fd_sc_hd__mux2_1 _10927_ (.A0(\sub1.data_o[116] ),
    .A1(_06669_),
    .S(_05608_),
    .X(_06670_));
 sky130_fd_sc_hd__a31o_1 _10928_ (.A1(_06630_),
    .A2(_06514_),
    .A3(\sub1.data_o[116] ),
    .B1(_05675_),
    .X(_06671_));
 sky130_fd_sc_hd__a21o_1 _10929_ (.A1(_05574_),
    .A2(_06670_),
    .B1(_06671_),
    .X(_06672_));
 sky130_fd_sc_hd__o21a_1 _10930_ (.A1(\mix1.data_o[116] ),
    .A2(_04626_),
    .B1(_05617_),
    .X(_06673_));
 sky130_fd_sc_hd__a221o_1 _10931_ (.A1(\sub1.data_o[116] ),
    .A2(_06513_),
    .B1(_06672_),
    .B2(_06673_),
    .C1(_04610_),
    .X(_06674_));
 sky130_fd_sc_hd__o21ai_1 _10932_ (.A1(_05623_),
    .A2(_06670_),
    .B1(_06674_),
    .Y(_06675_));
 sky130_fd_sc_hd__mux2_2 _10933_ (.A0(net148),
    .A1(\ks1.key_reg[116] ),
    .S(_04639_),
    .X(_06676_));
 sky130_fd_sc_hd__xnor2_1 _10934_ (.A(_06675_),
    .B(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(\addroundkey_data_o[116] ),
    .A1(_06677_),
    .S(_06612_),
    .X(_06678_));
 sky130_fd_sc_hd__clkbuf_1 _10936_ (.A(_06678_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(net20),
    .A1(\mix1.data_o[117] ),
    .S(_05602_),
    .X(_06679_));
 sky130_fd_sc_hd__mux2_1 _10938_ (.A0(\sub1.data_o[117] ),
    .A1(_06679_),
    .S(_05608_),
    .X(_06680_));
 sky130_fd_sc_hd__a31o_1 _10939_ (.A1(_06630_),
    .A2(\sub1.ready_o ),
    .A3(\sub1.data_o[117] ),
    .B1(_05675_),
    .X(_06681_));
 sky130_fd_sc_hd__a21o_1 _10940_ (.A1(_05574_),
    .A2(_06680_),
    .B1(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__o21a_1 _10941_ (.A1(\mix1.data_o[117] ),
    .A2(_04626_),
    .B1(_05617_),
    .X(_06683_));
 sky130_fd_sc_hd__a221o_1 _10942_ (.A1(\sub1.data_o[117] ),
    .A2(_05613_),
    .B1(_06682_),
    .B2(_06683_),
    .C1(_04610_),
    .X(_06684_));
 sky130_fd_sc_hd__o21ai_4 _10943_ (.A1(_05623_),
    .A2(_06680_),
    .B1(_06684_),
    .Y(_06685_));
 sky130_fd_sc_hd__mux2_1 _10944_ (.A0(net149),
    .A1(\ks1.key_reg[117] ),
    .S(_04639_),
    .X(_06686_));
 sky130_fd_sc_hd__xnor2_1 _10945_ (.A(_06685_),
    .B(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__mux2_1 _10946_ (.A0(\addroundkey_data_o[117] ),
    .A1(_06687_),
    .S(_06612_),
    .X(_06688_));
 sky130_fd_sc_hd__clkbuf_1 _10947_ (.A(_06688_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _10948_ (.A0(net21),
    .A1(\mix1.data_o[118] ),
    .S(_05602_),
    .X(_06689_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(\sub1.data_o[118] ),
    .A1(_06689_),
    .S(_05608_),
    .X(_06690_));
 sky130_fd_sc_hd__a31o_1 _10950_ (.A1(_06630_),
    .A2(\sub1.ready_o ),
    .A3(\sub1.data_o[118] ),
    .B1(_05675_),
    .X(_06691_));
 sky130_fd_sc_hd__a21o_1 _10951_ (.A1(_05574_),
    .A2(_06690_),
    .B1(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__o21a_1 _10952_ (.A1(\mix1.data_o[118] ),
    .A2(_04626_),
    .B1(_05617_),
    .X(_06693_));
 sky130_fd_sc_hd__a221o_1 _10953_ (.A1(\sub1.data_o[118] ),
    .A2(_05613_),
    .B1(_06692_),
    .B2(_06693_),
    .C1(_04610_),
    .X(_06694_));
 sky130_fd_sc_hd__o21ai_1 _10954_ (.A1(_05623_),
    .A2(_06690_),
    .B1(_06694_),
    .Y(_06695_));
 sky130_fd_sc_hd__mux2_2 _10955_ (.A0(net150),
    .A1(\ks1.key_reg[118] ),
    .S(_04639_),
    .X(_06696_));
 sky130_fd_sc_hd__xnor2_1 _10956_ (.A(_06695_),
    .B(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__mux2_1 _10957_ (.A0(\addroundkey_data_o[118] ),
    .A1(_06697_),
    .S(_06612_),
    .X(_06698_));
 sky130_fd_sc_hd__clkbuf_1 _10958_ (.A(_06698_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _10959_ (.A0(net22),
    .A1(\mix1.data_o[119] ),
    .S(_05602_),
    .X(_06699_));
 sky130_fd_sc_hd__mux2_1 _10960_ (.A0(\sub1.data_o[119] ),
    .A1(_06699_),
    .S(_05608_),
    .X(_06700_));
 sky130_fd_sc_hd__a31o_1 _10961_ (.A1(_06630_),
    .A2(\sub1.ready_o ),
    .A3(\sub1.data_o[119] ),
    .B1(_05675_),
    .X(_06701_));
 sky130_fd_sc_hd__a21o_1 _10962_ (.A1(_05574_),
    .A2(_06700_),
    .B1(_06701_),
    .X(_06702_));
 sky130_fd_sc_hd__o21a_1 _10963_ (.A1(\mix1.data_o[119] ),
    .A2(_04626_),
    .B1(_05617_),
    .X(_06703_));
 sky130_fd_sc_hd__a221o_1 _10964_ (.A1(\sub1.data_o[119] ),
    .A2(_05613_),
    .B1(_06702_),
    .B2(_06703_),
    .C1(_04610_),
    .X(_06704_));
 sky130_fd_sc_hd__o21ai_4 _10965_ (.A1(_05623_),
    .A2(_06700_),
    .B1(_06704_),
    .Y(_06705_));
 sky130_fd_sc_hd__mux2_1 _10966_ (.A0(net151),
    .A1(\ks1.key_reg[119] ),
    .S(_04639_),
    .X(_06706_));
 sky130_fd_sc_hd__xnor2_1 _10967_ (.A(_06705_),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(\addroundkey_data_o[119] ),
    .A1(_06707_),
    .S(_05696_),
    .X(_06708_));
 sky130_fd_sc_hd__clkbuf_1 _10969_ (.A(_06708_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(net24),
    .A1(\mix1.data_o[120] ),
    .S(_06571_),
    .X(_06709_));
 sky130_fd_sc_hd__mux2_1 _10971_ (.A0(\sub1.data_o[120] ),
    .A1(_06709_),
    .S(_06573_),
    .X(_06710_));
 sky130_fd_sc_hd__a32o_1 _10972_ (.A1(\mix1.data_o[120] ),
    .A2(_05676_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[120] ),
    .X(_06711_));
 sky130_fd_sc_hd__a22o_1 _10973_ (.A1(_06583_),
    .A2(_06710_),
    .B1(_06711_),
    .B2(_06587_),
    .X(_06712_));
 sky130_fd_sc_hd__mux2_1 _10974_ (.A0(net153),
    .A1(\ks1.key_reg[120] ),
    .S(_06579_),
    .X(_06713_));
 sky130_fd_sc_hd__xor2_1 _10975_ (.A(_06712_),
    .B(_06713_),
    .X(_06714_));
 sky130_fd_sc_hd__mux2_1 _10976_ (.A0(\addroundkey_data_o[120] ),
    .A1(_06714_),
    .S(_05696_),
    .X(_06715_));
 sky130_fd_sc_hd__clkbuf_1 _10977_ (.A(_06715_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _10978_ (.A0(net25),
    .A1(\mix1.data_o[121] ),
    .S(_06571_),
    .X(_06716_));
 sky130_fd_sc_hd__mux2_1 _10979_ (.A0(\sub1.data_o[121] ),
    .A1(_06716_),
    .S(_06573_),
    .X(_06717_));
 sky130_fd_sc_hd__a32o_1 _10980_ (.A1(\mix1.data_o[121] ),
    .A2(_05676_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[121] ),
    .X(_06718_));
 sky130_fd_sc_hd__a22o_1 _10981_ (.A1(_06583_),
    .A2(_06717_),
    .B1(_06718_),
    .B2(_06587_),
    .X(_06719_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(net154),
    .A1(\ks1.key_reg[121] ),
    .S(_06579_),
    .X(_06720_));
 sky130_fd_sc_hd__xor2_1 _10983_ (.A(_06719_),
    .B(_06720_),
    .X(_06721_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(\addroundkey_data_o[121] ),
    .A1(_06721_),
    .S(_05696_),
    .X(_06722_));
 sky130_fd_sc_hd__clkbuf_1 _10985_ (.A(_06722_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _10986_ (.A0(net26),
    .A1(\mix1.data_o[122] ),
    .S(_06571_),
    .X(_06723_));
 sky130_fd_sc_hd__mux2_1 _10987_ (.A0(\sub1.data_o[122] ),
    .A1(_06723_),
    .S(_06573_),
    .X(_06724_));
 sky130_fd_sc_hd__a32o_1 _10988_ (.A1(\mix1.data_o[122] ),
    .A2(_05676_),
    .A3(_06575_),
    .B1(_06576_),
    .B2(\sub1.data_o[122] ),
    .X(_06725_));
 sky130_fd_sc_hd__a22o_1 _10989_ (.A1(_06583_),
    .A2(_06724_),
    .B1(_06725_),
    .B2(_06587_),
    .X(_06726_));
 sky130_fd_sc_hd__mux2_1 _10990_ (.A0(net155),
    .A1(\ks1.key_reg[122] ),
    .S(_06579_),
    .X(_06727_));
 sky130_fd_sc_hd__xor2_1 _10991_ (.A(_06726_),
    .B(_06727_),
    .X(_06728_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(\addroundkey_data_o[122] ),
    .A1(_06728_),
    .S(_05696_),
    .X(_06729_));
 sky130_fd_sc_hd__clkbuf_1 _10993_ (.A(_06729_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _10994_ (.A0(net27),
    .A1(\mix1.data_o[123] ),
    .S(_05603_),
    .X(_06730_));
 sky130_fd_sc_hd__mux2_1 _10995_ (.A0(\sub1.data_o[123] ),
    .A1(_06730_),
    .S(_05609_),
    .X(_06731_));
 sky130_fd_sc_hd__a32o_1 _10996_ (.A1(\mix1.data_o[123] ),
    .A2(_05676_),
    .A3(_05758_),
    .B1(_05620_),
    .B2(\sub1.data_o[123] ),
    .X(_06732_));
 sky130_fd_sc_hd__a22o_1 _10997_ (.A1(_06583_),
    .A2(_06731_),
    .B1(_06732_),
    .B2(_06587_),
    .X(_06733_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(net156),
    .A1(\ks1.key_reg[123] ),
    .S(_05762_),
    .X(_06734_));
 sky130_fd_sc_hd__xor2_1 _10999_ (.A(_06733_),
    .B(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(\addroundkey_data_o[123] ),
    .A1(_06735_),
    .S(_05696_),
    .X(_06736_));
 sky130_fd_sc_hd__clkbuf_1 _11001_ (.A(_06736_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _11002_ (.A0(net28),
    .A1(\mix1.data_o[124] ),
    .S(_05603_),
    .X(_06737_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(\sub1.data_o[124] ),
    .A1(_06737_),
    .S(_05609_),
    .X(_06738_));
 sky130_fd_sc_hd__a32o_1 _11004_ (.A1(\mix1.data_o[124] ),
    .A2(_05676_),
    .A3(_05758_),
    .B1(_05620_),
    .B2(\sub1.data_o[124] ),
    .X(_06739_));
 sky130_fd_sc_hd__a22o_1 _11005_ (.A1(_05615_),
    .A2(_06738_),
    .B1(_06739_),
    .B2(_05567_),
    .X(_06740_));
 sky130_fd_sc_hd__mux2_1 _11006_ (.A0(net157),
    .A1(\ks1.key_reg[124] ),
    .S(_05762_),
    .X(_06741_));
 sky130_fd_sc_hd__xor2_1 _11007_ (.A(_06740_),
    .B(_06741_),
    .X(_06742_));
 sky130_fd_sc_hd__mux2_1 _11008_ (.A0(\addroundkey_data_o[124] ),
    .A1(_06742_),
    .S(_05696_),
    .X(_06743_));
 sky130_fd_sc_hd__clkbuf_1 _11009_ (.A(_06743_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _11010_ (.A0(net29),
    .A1(\mix1.data_o[125] ),
    .S(_05603_),
    .X(_06744_));
 sky130_fd_sc_hd__mux2_1 _11011_ (.A0(\sub1.data_o[125] ),
    .A1(_06744_),
    .S(_05609_),
    .X(_06745_));
 sky130_fd_sc_hd__a32o_1 _11012_ (.A1(\mix1.data_o[125] ),
    .A2(_05676_),
    .A3(_05758_),
    .B1(_05620_),
    .B2(\sub1.data_o[125] ),
    .X(_06746_));
 sky130_fd_sc_hd__a22o_1 _11013_ (.A1(_05615_),
    .A2(_06745_),
    .B1(_06746_),
    .B2(_05567_),
    .X(_06747_));
 sky130_fd_sc_hd__mux2_1 _11014_ (.A0(net158),
    .A1(\ks1.key_reg[125] ),
    .S(_05762_),
    .X(_06748_));
 sky130_fd_sc_hd__xor2_1 _11015_ (.A(_06747_),
    .B(_06748_),
    .X(_06749_));
 sky130_fd_sc_hd__mux2_1 _11016_ (.A0(\addroundkey_data_o[125] ),
    .A1(_06749_),
    .S(_05696_),
    .X(_06750_));
 sky130_fd_sc_hd__clkbuf_1 _11017_ (.A(_06750_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _11018_ (.A0(net30),
    .A1(\mix1.data_o[126] ),
    .S(_05603_),
    .X(_06751_));
 sky130_fd_sc_hd__mux2_1 _11019_ (.A0(\sub1.data_o[126] ),
    .A1(_06751_),
    .S(_05609_),
    .X(_06752_));
 sky130_fd_sc_hd__a32o_1 _11020_ (.A1(\mix1.data_o[126] ),
    .A2(_05676_),
    .A3(_05758_),
    .B1(_05620_),
    .B2(\sub1.data_o[126] ),
    .X(_06753_));
 sky130_fd_sc_hd__a22o_1 _11021_ (.A1(_05615_),
    .A2(_06752_),
    .B1(_06753_),
    .B2(_05567_),
    .X(_06754_));
 sky130_fd_sc_hd__mux2_1 _11022_ (.A0(net159),
    .A1(\ks1.key_reg[126] ),
    .S(_05762_),
    .X(_06755_));
 sky130_fd_sc_hd__xor2_1 _11023_ (.A(_06754_),
    .B(_06755_),
    .X(_06756_));
 sky130_fd_sc_hd__mux2_1 _11024_ (.A0(\addroundkey_data_o[126] ),
    .A1(_06756_),
    .S(_05696_),
    .X(_06757_));
 sky130_fd_sc_hd__clkbuf_1 _11025_ (.A(_06757_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _11026_ (.A0(net31),
    .A1(\mix1.data_o[127] ),
    .S(_05603_),
    .X(_06758_));
 sky130_fd_sc_hd__mux2_1 _11027_ (.A0(\sub1.data_o[127] ),
    .A1(_06758_),
    .S(_05609_),
    .X(_06759_));
 sky130_fd_sc_hd__a32o_1 _11028_ (.A1(\mix1.data_o[127] ),
    .A2(_05676_),
    .A3(_05758_),
    .B1(_05620_),
    .B2(\sub1.data_o[127] ),
    .X(_06760_));
 sky130_fd_sc_hd__a22o_1 _11029_ (.A1(_05615_),
    .A2(_06759_),
    .B1(_06760_),
    .B2(_05567_),
    .X(_06761_));
 sky130_fd_sc_hd__mux2_1 _11030_ (.A0(net160),
    .A1(\ks1.key_reg[127] ),
    .S(_05762_),
    .X(_06762_));
 sky130_fd_sc_hd__xor2_1 _11031_ (.A(_06761_),
    .B(_06762_),
    .X(_06763_));
 sky130_fd_sc_hd__mux2_1 _11032_ (.A0(\addroundkey_data_o[127] ),
    .A1(_06763_),
    .S(_05696_),
    .X(_06764_));
 sky130_fd_sc_hd__clkbuf_1 _11033_ (.A(_06764_),
    .X(_00280_));
 sky130_fd_sc_hd__inv_2 _11034_ (.A(_05266_),
    .Y(_06765_));
 sky130_fd_sc_hd__or3b_1 _11035_ (.A(_05249_),
    .B(_05250_),
    .C_N(net597),
    .X(_06766_));
 sky130_fd_sc_hd__or4_2 _11036_ (.A(\fifo_bank_register.write_ptr[2] ),
    .B(_05254_),
    .C(_06765_),
    .D(_06766_),
    .X(_06767_));
 sky130_fd_sc_hd__buf_4 _11037_ (.A(_06767_),
    .X(_06768_));
 sky130_fd_sc_hd__clkbuf_4 _11038_ (.A(_06768_),
    .X(_06769_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(_05248_),
    .A1(\fifo_bank_register.bank[8][0] ),
    .S(_06769_),
    .X(_06770_));
 sky130_fd_sc_hd__clkbuf_1 _11040_ (.A(_06770_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _11041_ (.A0(_05272_),
    .A1(\fifo_bank_register.bank[8][1] ),
    .S(_06769_),
    .X(_06771_));
 sky130_fd_sc_hd__clkbuf_1 _11042_ (.A(_06771_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _11043_ (.A0(_05274_),
    .A1(\fifo_bank_register.bank[8][2] ),
    .S(_06769_),
    .X(_06772_));
 sky130_fd_sc_hd__clkbuf_1 _11044_ (.A(_06772_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(_05276_),
    .A1(\fifo_bank_register.bank[8][3] ),
    .S(_06769_),
    .X(_06773_));
 sky130_fd_sc_hd__clkbuf_1 _11046_ (.A(_06773_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _11047_ (.A0(_05278_),
    .A1(\fifo_bank_register.bank[8][4] ),
    .S(_06769_),
    .X(_06774_));
 sky130_fd_sc_hd__clkbuf_1 _11048_ (.A(_06774_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _11049_ (.A0(_05280_),
    .A1(\fifo_bank_register.bank[8][5] ),
    .S(_06769_),
    .X(_06775_));
 sky130_fd_sc_hd__clkbuf_1 _11050_ (.A(_06775_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _11051_ (.A0(_05282_),
    .A1(\fifo_bank_register.bank[8][6] ),
    .S(_06769_),
    .X(_06776_));
 sky130_fd_sc_hd__clkbuf_1 _11052_ (.A(_06776_),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _11053_ (.A0(_05284_),
    .A1(\fifo_bank_register.bank[8][7] ),
    .S(_06769_),
    .X(_06777_));
 sky130_fd_sc_hd__clkbuf_1 _11054_ (.A(_06777_),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _11055_ (.A0(_05286_),
    .A1(\fifo_bank_register.bank[8][8] ),
    .S(_06769_),
    .X(_06778_));
 sky130_fd_sc_hd__clkbuf_1 _11056_ (.A(_06778_),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _11057_ (.A0(_05288_),
    .A1(\fifo_bank_register.bank[8][9] ),
    .S(_06769_),
    .X(_06779_));
 sky130_fd_sc_hd__clkbuf_1 _11058_ (.A(_06779_),
    .X(_00290_));
 sky130_fd_sc_hd__buf_4 _11059_ (.A(_06768_),
    .X(_06780_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(_05290_),
    .A1(\fifo_bank_register.bank[8][10] ),
    .S(_06780_),
    .X(_06781_));
 sky130_fd_sc_hd__clkbuf_1 _11061_ (.A(_06781_),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(_05293_),
    .A1(\fifo_bank_register.bank[8][11] ),
    .S(_06780_),
    .X(_06782_));
 sky130_fd_sc_hd__clkbuf_1 _11063_ (.A(_06782_),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(_05295_),
    .A1(\fifo_bank_register.bank[8][12] ),
    .S(_06780_),
    .X(_06783_));
 sky130_fd_sc_hd__clkbuf_1 _11065_ (.A(_06783_),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(_05297_),
    .A1(\fifo_bank_register.bank[8][13] ),
    .S(_06780_),
    .X(_06784_));
 sky130_fd_sc_hd__clkbuf_1 _11067_ (.A(_06784_),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(_05299_),
    .A1(\fifo_bank_register.bank[8][14] ),
    .S(_06780_),
    .X(_06785_));
 sky130_fd_sc_hd__clkbuf_1 _11069_ (.A(_06785_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _11070_ (.A0(_05301_),
    .A1(\fifo_bank_register.bank[8][15] ),
    .S(_06780_),
    .X(_06786_));
 sky130_fd_sc_hd__clkbuf_1 _11071_ (.A(_06786_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _11072_ (.A0(_05303_),
    .A1(\fifo_bank_register.bank[8][16] ),
    .S(_06780_),
    .X(_06787_));
 sky130_fd_sc_hd__clkbuf_1 _11073_ (.A(_06787_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _11074_ (.A0(_05305_),
    .A1(\fifo_bank_register.bank[8][17] ),
    .S(_06780_),
    .X(_06788_));
 sky130_fd_sc_hd__clkbuf_1 _11075_ (.A(_06788_),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _11076_ (.A0(_05307_),
    .A1(\fifo_bank_register.bank[8][18] ),
    .S(_06780_),
    .X(_06789_));
 sky130_fd_sc_hd__clkbuf_1 _11077_ (.A(_06789_),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _11078_ (.A0(_05309_),
    .A1(\fifo_bank_register.bank[8][19] ),
    .S(_06780_),
    .X(_06790_));
 sky130_fd_sc_hd__clkbuf_1 _11079_ (.A(_06790_),
    .X(_00300_));
 sky130_fd_sc_hd__buf_8 _11080_ (.A(_06767_),
    .X(_06791_));
 sky130_fd_sc_hd__buf_4 _11081_ (.A(_06791_),
    .X(_06792_));
 sky130_fd_sc_hd__mux2_1 _11082_ (.A0(_05311_),
    .A1(\fifo_bank_register.bank[8][20] ),
    .S(_06792_),
    .X(_06793_));
 sky130_fd_sc_hd__clkbuf_1 _11083_ (.A(_06793_),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(_05315_),
    .A1(\fifo_bank_register.bank[8][21] ),
    .S(_06792_),
    .X(_06794_));
 sky130_fd_sc_hd__clkbuf_1 _11085_ (.A(_06794_),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _11086_ (.A0(_05317_),
    .A1(\fifo_bank_register.bank[8][22] ),
    .S(_06792_),
    .X(_06795_));
 sky130_fd_sc_hd__clkbuf_1 _11087_ (.A(_06795_),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(_05319_),
    .A1(\fifo_bank_register.bank[8][23] ),
    .S(_06792_),
    .X(_06796_));
 sky130_fd_sc_hd__clkbuf_1 _11089_ (.A(_06796_),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _11090_ (.A0(_05321_),
    .A1(\fifo_bank_register.bank[8][24] ),
    .S(_06792_),
    .X(_06797_));
 sky130_fd_sc_hd__clkbuf_1 _11091_ (.A(_06797_),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(_05323_),
    .A1(\fifo_bank_register.bank[8][25] ),
    .S(_06792_),
    .X(_06798_));
 sky130_fd_sc_hd__clkbuf_1 _11093_ (.A(_06798_),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(_05325_),
    .A1(\fifo_bank_register.bank[8][26] ),
    .S(_06792_),
    .X(_06799_));
 sky130_fd_sc_hd__clkbuf_1 _11095_ (.A(_06799_),
    .X(_00307_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(_05327_),
    .A1(\fifo_bank_register.bank[8][27] ),
    .S(_06792_),
    .X(_06800_));
 sky130_fd_sc_hd__clkbuf_1 _11097_ (.A(_06800_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(_05329_),
    .A1(\fifo_bank_register.bank[8][28] ),
    .S(_06792_),
    .X(_06801_));
 sky130_fd_sc_hd__clkbuf_1 _11099_ (.A(_06801_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(_05331_),
    .A1(\fifo_bank_register.bank[8][29] ),
    .S(_06792_),
    .X(_06802_));
 sky130_fd_sc_hd__clkbuf_1 _11101_ (.A(_06802_),
    .X(_00310_));
 sky130_fd_sc_hd__buf_4 _11102_ (.A(_06791_),
    .X(_06803_));
 sky130_fd_sc_hd__mux2_1 _11103_ (.A0(_05333_),
    .A1(\fifo_bank_register.bank[8][30] ),
    .S(_06803_),
    .X(_06804_));
 sky130_fd_sc_hd__clkbuf_1 _11104_ (.A(_06804_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _11105_ (.A0(_05336_),
    .A1(\fifo_bank_register.bank[8][31] ),
    .S(_06803_),
    .X(_06805_));
 sky130_fd_sc_hd__clkbuf_1 _11106_ (.A(_06805_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _11107_ (.A0(_05338_),
    .A1(\fifo_bank_register.bank[8][32] ),
    .S(_06803_),
    .X(_06806_));
 sky130_fd_sc_hd__clkbuf_1 _11108_ (.A(_06806_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _11109_ (.A0(_05340_),
    .A1(\fifo_bank_register.bank[8][33] ),
    .S(_06803_),
    .X(_06807_));
 sky130_fd_sc_hd__clkbuf_1 _11110_ (.A(_06807_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _11111_ (.A0(_05342_),
    .A1(\fifo_bank_register.bank[8][34] ),
    .S(_06803_),
    .X(_06808_));
 sky130_fd_sc_hd__clkbuf_1 _11112_ (.A(_06808_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _11113_ (.A0(_05344_),
    .A1(\fifo_bank_register.bank[8][35] ),
    .S(_06803_),
    .X(_06809_));
 sky130_fd_sc_hd__clkbuf_1 _11114_ (.A(_06809_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(_05346_),
    .A1(\fifo_bank_register.bank[8][36] ),
    .S(_06803_),
    .X(_06810_));
 sky130_fd_sc_hd__clkbuf_1 _11116_ (.A(_06810_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(_05348_),
    .A1(\fifo_bank_register.bank[8][37] ),
    .S(_06803_),
    .X(_06811_));
 sky130_fd_sc_hd__clkbuf_1 _11118_ (.A(_06811_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(_05350_),
    .A1(\fifo_bank_register.bank[8][38] ),
    .S(_06803_),
    .X(_06812_));
 sky130_fd_sc_hd__clkbuf_1 _11120_ (.A(_06812_),
    .X(_00319_));
 sky130_fd_sc_hd__mux2_1 _11121_ (.A0(_05352_),
    .A1(\fifo_bank_register.bank[8][39] ),
    .S(_06803_),
    .X(_06813_));
 sky130_fd_sc_hd__clkbuf_1 _11122_ (.A(_06813_),
    .X(_00320_));
 sky130_fd_sc_hd__buf_4 _11123_ (.A(_06791_),
    .X(_06814_));
 sky130_fd_sc_hd__mux2_1 _11124_ (.A0(_05354_),
    .A1(\fifo_bank_register.bank[8][40] ),
    .S(_06814_),
    .X(_06815_));
 sky130_fd_sc_hd__clkbuf_1 _11125_ (.A(_06815_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _11126_ (.A0(_05357_),
    .A1(\fifo_bank_register.bank[8][41] ),
    .S(_06814_),
    .X(_06816_));
 sky130_fd_sc_hd__clkbuf_1 _11127_ (.A(_06816_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _11128_ (.A0(_05359_),
    .A1(\fifo_bank_register.bank[8][42] ),
    .S(_06814_),
    .X(_06817_));
 sky130_fd_sc_hd__clkbuf_1 _11129_ (.A(_06817_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _11130_ (.A0(_05361_),
    .A1(\fifo_bank_register.bank[8][43] ),
    .S(_06814_),
    .X(_06818_));
 sky130_fd_sc_hd__clkbuf_1 _11131_ (.A(_06818_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _11132_ (.A0(_05363_),
    .A1(\fifo_bank_register.bank[8][44] ),
    .S(_06814_),
    .X(_06819_));
 sky130_fd_sc_hd__clkbuf_1 _11133_ (.A(_06819_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _11134_ (.A0(_05365_),
    .A1(\fifo_bank_register.bank[8][45] ),
    .S(_06814_),
    .X(_06820_));
 sky130_fd_sc_hd__clkbuf_1 _11135_ (.A(_06820_),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _11136_ (.A0(_05367_),
    .A1(\fifo_bank_register.bank[8][46] ),
    .S(_06814_),
    .X(_06821_));
 sky130_fd_sc_hd__clkbuf_1 _11137_ (.A(_06821_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _11138_ (.A0(_05369_),
    .A1(\fifo_bank_register.bank[8][47] ),
    .S(_06814_),
    .X(_06822_));
 sky130_fd_sc_hd__clkbuf_1 _11139_ (.A(_06822_),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _11140_ (.A0(_05371_),
    .A1(\fifo_bank_register.bank[8][48] ),
    .S(_06814_),
    .X(_06823_));
 sky130_fd_sc_hd__clkbuf_1 _11141_ (.A(_06823_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _11142_ (.A0(_05373_),
    .A1(\fifo_bank_register.bank[8][49] ),
    .S(_06814_),
    .X(_06824_));
 sky130_fd_sc_hd__clkbuf_1 _11143_ (.A(_06824_),
    .X(_00330_));
 sky130_fd_sc_hd__buf_4 _11144_ (.A(_06791_),
    .X(_06825_));
 sky130_fd_sc_hd__mux2_1 _11145_ (.A0(_05375_),
    .A1(\fifo_bank_register.bank[8][50] ),
    .S(_06825_),
    .X(_06826_));
 sky130_fd_sc_hd__clkbuf_1 _11146_ (.A(_06826_),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _11147_ (.A0(_05378_),
    .A1(\fifo_bank_register.bank[8][51] ),
    .S(_06825_),
    .X(_06827_));
 sky130_fd_sc_hd__clkbuf_1 _11148_ (.A(_06827_),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _11149_ (.A0(_05380_),
    .A1(\fifo_bank_register.bank[8][52] ),
    .S(_06825_),
    .X(_06828_));
 sky130_fd_sc_hd__clkbuf_1 _11150_ (.A(_06828_),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _11151_ (.A0(_05382_),
    .A1(\fifo_bank_register.bank[8][53] ),
    .S(_06825_),
    .X(_06829_));
 sky130_fd_sc_hd__clkbuf_1 _11152_ (.A(_06829_),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _11153_ (.A0(_05384_),
    .A1(\fifo_bank_register.bank[8][54] ),
    .S(_06825_),
    .X(_06830_));
 sky130_fd_sc_hd__clkbuf_1 _11154_ (.A(_06830_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _11155_ (.A0(_05386_),
    .A1(\fifo_bank_register.bank[8][55] ),
    .S(_06825_),
    .X(_06831_));
 sky130_fd_sc_hd__clkbuf_1 _11156_ (.A(_06831_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _11157_ (.A0(_05388_),
    .A1(\fifo_bank_register.bank[8][56] ),
    .S(_06825_),
    .X(_06832_));
 sky130_fd_sc_hd__clkbuf_1 _11158_ (.A(_06832_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _11159_ (.A0(_05390_),
    .A1(\fifo_bank_register.bank[8][57] ),
    .S(_06825_),
    .X(_06833_));
 sky130_fd_sc_hd__clkbuf_1 _11160_ (.A(_06833_),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _11161_ (.A0(_05392_),
    .A1(\fifo_bank_register.bank[8][58] ),
    .S(_06825_),
    .X(_06834_));
 sky130_fd_sc_hd__clkbuf_1 _11162_ (.A(_06834_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _11163_ (.A0(_05394_),
    .A1(\fifo_bank_register.bank[8][59] ),
    .S(_06825_),
    .X(_06835_));
 sky130_fd_sc_hd__clkbuf_1 _11164_ (.A(_06835_),
    .X(_00340_));
 sky130_fd_sc_hd__buf_4 _11165_ (.A(_06791_),
    .X(_06836_));
 sky130_fd_sc_hd__mux2_1 _11166_ (.A0(_05396_),
    .A1(\fifo_bank_register.bank[8][60] ),
    .S(_06836_),
    .X(_06837_));
 sky130_fd_sc_hd__clkbuf_1 _11167_ (.A(_06837_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _11168_ (.A0(_05399_),
    .A1(\fifo_bank_register.bank[8][61] ),
    .S(_06836_),
    .X(_06838_));
 sky130_fd_sc_hd__clkbuf_1 _11169_ (.A(_06838_),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _11170_ (.A0(_05401_),
    .A1(\fifo_bank_register.bank[8][62] ),
    .S(_06836_),
    .X(_06839_));
 sky130_fd_sc_hd__clkbuf_1 _11171_ (.A(_06839_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _11172_ (.A0(_05403_),
    .A1(\fifo_bank_register.bank[8][63] ),
    .S(_06836_),
    .X(_06840_));
 sky130_fd_sc_hd__clkbuf_1 _11173_ (.A(_06840_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _11174_ (.A0(_05405_),
    .A1(\fifo_bank_register.bank[8][64] ),
    .S(_06836_),
    .X(_06841_));
 sky130_fd_sc_hd__clkbuf_1 _11175_ (.A(_06841_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _11176_ (.A0(_05407_),
    .A1(\fifo_bank_register.bank[8][65] ),
    .S(_06836_),
    .X(_06842_));
 sky130_fd_sc_hd__clkbuf_1 _11177_ (.A(_06842_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _11178_ (.A0(_05409_),
    .A1(\fifo_bank_register.bank[8][66] ),
    .S(_06836_),
    .X(_06843_));
 sky130_fd_sc_hd__clkbuf_1 _11179_ (.A(_06843_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _11180_ (.A0(_05411_),
    .A1(\fifo_bank_register.bank[8][67] ),
    .S(_06836_),
    .X(_06844_));
 sky130_fd_sc_hd__clkbuf_1 _11181_ (.A(_06844_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _11182_ (.A0(_05413_),
    .A1(\fifo_bank_register.bank[8][68] ),
    .S(_06836_),
    .X(_06845_));
 sky130_fd_sc_hd__clkbuf_1 _11183_ (.A(_06845_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _11184_ (.A0(_05415_),
    .A1(\fifo_bank_register.bank[8][69] ),
    .S(_06836_),
    .X(_06846_));
 sky130_fd_sc_hd__clkbuf_1 _11185_ (.A(_06846_),
    .X(_00350_));
 sky130_fd_sc_hd__buf_4 _11186_ (.A(_06791_),
    .X(_06847_));
 sky130_fd_sc_hd__mux2_1 _11187_ (.A0(_05417_),
    .A1(\fifo_bank_register.bank[8][70] ),
    .S(_06847_),
    .X(_06848_));
 sky130_fd_sc_hd__clkbuf_1 _11188_ (.A(_06848_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _11189_ (.A0(_05420_),
    .A1(\fifo_bank_register.bank[8][71] ),
    .S(_06847_),
    .X(_06849_));
 sky130_fd_sc_hd__clkbuf_1 _11190_ (.A(_06849_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _11191_ (.A0(_05422_),
    .A1(\fifo_bank_register.bank[8][72] ),
    .S(_06847_),
    .X(_06850_));
 sky130_fd_sc_hd__clkbuf_1 _11192_ (.A(_06850_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _11193_ (.A0(_05424_),
    .A1(\fifo_bank_register.bank[8][73] ),
    .S(_06847_),
    .X(_06851_));
 sky130_fd_sc_hd__clkbuf_1 _11194_ (.A(_06851_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _11195_ (.A0(_05426_),
    .A1(\fifo_bank_register.bank[8][74] ),
    .S(_06847_),
    .X(_06852_));
 sky130_fd_sc_hd__clkbuf_1 _11196_ (.A(_06852_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _11197_ (.A0(_05428_),
    .A1(\fifo_bank_register.bank[8][75] ),
    .S(_06847_),
    .X(_06853_));
 sky130_fd_sc_hd__clkbuf_1 _11198_ (.A(_06853_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _11199_ (.A0(_05430_),
    .A1(\fifo_bank_register.bank[8][76] ),
    .S(_06847_),
    .X(_06854_));
 sky130_fd_sc_hd__clkbuf_1 _11200_ (.A(_06854_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _11201_ (.A0(_05432_),
    .A1(\fifo_bank_register.bank[8][77] ),
    .S(_06847_),
    .X(_06855_));
 sky130_fd_sc_hd__clkbuf_1 _11202_ (.A(_06855_),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _11203_ (.A0(_05434_),
    .A1(\fifo_bank_register.bank[8][78] ),
    .S(_06847_),
    .X(_06856_));
 sky130_fd_sc_hd__clkbuf_1 _11204_ (.A(_06856_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(_05436_),
    .A1(\fifo_bank_register.bank[8][79] ),
    .S(_06847_),
    .X(_06857_));
 sky130_fd_sc_hd__clkbuf_1 _11206_ (.A(_06857_),
    .X(_00360_));
 sky130_fd_sc_hd__buf_4 _11207_ (.A(_06791_),
    .X(_06858_));
 sky130_fd_sc_hd__mux2_1 _11208_ (.A0(_05438_),
    .A1(\fifo_bank_register.bank[8][80] ),
    .S(_06858_),
    .X(_06859_));
 sky130_fd_sc_hd__clkbuf_1 _11209_ (.A(_06859_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _11210_ (.A0(_05441_),
    .A1(\fifo_bank_register.bank[8][81] ),
    .S(_06858_),
    .X(_06860_));
 sky130_fd_sc_hd__clkbuf_1 _11211_ (.A(_06860_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _11212_ (.A0(_05443_),
    .A1(\fifo_bank_register.bank[8][82] ),
    .S(_06858_),
    .X(_06861_));
 sky130_fd_sc_hd__clkbuf_1 _11213_ (.A(_06861_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _11214_ (.A0(_05445_),
    .A1(\fifo_bank_register.bank[8][83] ),
    .S(_06858_),
    .X(_06862_));
 sky130_fd_sc_hd__clkbuf_1 _11215_ (.A(_06862_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _11216_ (.A0(_05447_),
    .A1(\fifo_bank_register.bank[8][84] ),
    .S(_06858_),
    .X(_06863_));
 sky130_fd_sc_hd__clkbuf_1 _11217_ (.A(_06863_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _11218_ (.A0(_05449_),
    .A1(\fifo_bank_register.bank[8][85] ),
    .S(_06858_),
    .X(_06864_));
 sky130_fd_sc_hd__clkbuf_1 _11219_ (.A(_06864_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _11220_ (.A0(_05451_),
    .A1(\fifo_bank_register.bank[8][86] ),
    .S(_06858_),
    .X(_06865_));
 sky130_fd_sc_hd__clkbuf_1 _11221_ (.A(_06865_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _11222_ (.A0(_05453_),
    .A1(\fifo_bank_register.bank[8][87] ),
    .S(_06858_),
    .X(_06866_));
 sky130_fd_sc_hd__clkbuf_1 _11223_ (.A(_06866_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _11224_ (.A0(_05455_),
    .A1(\fifo_bank_register.bank[8][88] ),
    .S(_06858_),
    .X(_06867_));
 sky130_fd_sc_hd__clkbuf_1 _11225_ (.A(_06867_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _11226_ (.A0(_05457_),
    .A1(\fifo_bank_register.bank[8][89] ),
    .S(_06858_),
    .X(_06868_));
 sky130_fd_sc_hd__clkbuf_1 _11227_ (.A(_06868_),
    .X(_00370_));
 sky130_fd_sc_hd__buf_4 _11228_ (.A(_06791_),
    .X(_06869_));
 sky130_fd_sc_hd__mux2_1 _11229_ (.A0(_05459_),
    .A1(\fifo_bank_register.bank[8][90] ),
    .S(_06869_),
    .X(_06870_));
 sky130_fd_sc_hd__clkbuf_1 _11230_ (.A(_06870_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _11231_ (.A0(_05462_),
    .A1(\fifo_bank_register.bank[8][91] ),
    .S(_06869_),
    .X(_06871_));
 sky130_fd_sc_hd__clkbuf_1 _11232_ (.A(_06871_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _11233_ (.A0(_05464_),
    .A1(\fifo_bank_register.bank[8][92] ),
    .S(_06869_),
    .X(_06872_));
 sky130_fd_sc_hd__clkbuf_1 _11234_ (.A(_06872_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _11235_ (.A0(_05466_),
    .A1(\fifo_bank_register.bank[8][93] ),
    .S(_06869_),
    .X(_06873_));
 sky130_fd_sc_hd__clkbuf_1 _11236_ (.A(_06873_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _11237_ (.A0(_05468_),
    .A1(\fifo_bank_register.bank[8][94] ),
    .S(_06869_),
    .X(_06874_));
 sky130_fd_sc_hd__clkbuf_1 _11238_ (.A(_06874_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _11239_ (.A0(_05470_),
    .A1(\fifo_bank_register.bank[8][95] ),
    .S(_06869_),
    .X(_06875_));
 sky130_fd_sc_hd__clkbuf_1 _11240_ (.A(_06875_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _11241_ (.A0(_05472_),
    .A1(\fifo_bank_register.bank[8][96] ),
    .S(_06869_),
    .X(_06876_));
 sky130_fd_sc_hd__clkbuf_1 _11242_ (.A(_06876_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _11243_ (.A0(_05474_),
    .A1(\fifo_bank_register.bank[8][97] ),
    .S(_06869_),
    .X(_06877_));
 sky130_fd_sc_hd__clkbuf_1 _11244_ (.A(_06877_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _11245_ (.A0(_05476_),
    .A1(\fifo_bank_register.bank[8][98] ),
    .S(_06869_),
    .X(_06878_));
 sky130_fd_sc_hd__clkbuf_1 _11246_ (.A(_06878_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _11247_ (.A0(_05478_),
    .A1(\fifo_bank_register.bank[8][99] ),
    .S(_06869_),
    .X(_06879_));
 sky130_fd_sc_hd__clkbuf_1 _11248_ (.A(_06879_),
    .X(_00380_));
 sky130_fd_sc_hd__buf_4 _11249_ (.A(_06791_),
    .X(_06880_));
 sky130_fd_sc_hd__mux2_1 _11250_ (.A0(_05480_),
    .A1(\fifo_bank_register.bank[8][100] ),
    .S(_06880_),
    .X(_06881_));
 sky130_fd_sc_hd__clkbuf_1 _11251_ (.A(_06881_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _11252_ (.A0(_05483_),
    .A1(\fifo_bank_register.bank[8][101] ),
    .S(_06880_),
    .X(_06882_));
 sky130_fd_sc_hd__clkbuf_1 _11253_ (.A(_06882_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _11254_ (.A0(_05485_),
    .A1(\fifo_bank_register.bank[8][102] ),
    .S(_06880_),
    .X(_06883_));
 sky130_fd_sc_hd__clkbuf_1 _11255_ (.A(_06883_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _11256_ (.A0(_05487_),
    .A1(\fifo_bank_register.bank[8][103] ),
    .S(_06880_),
    .X(_06884_));
 sky130_fd_sc_hd__clkbuf_1 _11257_ (.A(_06884_),
    .X(_00384_));
 sky130_fd_sc_hd__mux2_1 _11258_ (.A0(_05489_),
    .A1(\fifo_bank_register.bank[8][104] ),
    .S(_06880_),
    .X(_06885_));
 sky130_fd_sc_hd__clkbuf_1 _11259_ (.A(_06885_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _11260_ (.A0(_05491_),
    .A1(\fifo_bank_register.bank[8][105] ),
    .S(_06880_),
    .X(_06886_));
 sky130_fd_sc_hd__clkbuf_1 _11261_ (.A(_06886_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _11262_ (.A0(_05493_),
    .A1(\fifo_bank_register.bank[8][106] ),
    .S(_06880_),
    .X(_06887_));
 sky130_fd_sc_hd__clkbuf_1 _11263_ (.A(_06887_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _11264_ (.A0(_05495_),
    .A1(\fifo_bank_register.bank[8][107] ),
    .S(_06880_),
    .X(_06888_));
 sky130_fd_sc_hd__clkbuf_1 _11265_ (.A(_06888_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _11266_ (.A0(_05497_),
    .A1(\fifo_bank_register.bank[8][108] ),
    .S(_06880_),
    .X(_06889_));
 sky130_fd_sc_hd__clkbuf_1 _11267_ (.A(_06889_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _11268_ (.A0(_05499_),
    .A1(\fifo_bank_register.bank[8][109] ),
    .S(_06880_),
    .X(_06890_));
 sky130_fd_sc_hd__clkbuf_1 _11269_ (.A(_06890_),
    .X(_00390_));
 sky130_fd_sc_hd__buf_4 _11270_ (.A(_06791_),
    .X(_06891_));
 sky130_fd_sc_hd__mux2_1 _11271_ (.A0(_05501_),
    .A1(\fifo_bank_register.bank[8][110] ),
    .S(_06891_),
    .X(_06892_));
 sky130_fd_sc_hd__clkbuf_1 _11272_ (.A(_06892_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _11273_ (.A0(_05504_),
    .A1(\fifo_bank_register.bank[8][111] ),
    .S(_06891_),
    .X(_06893_));
 sky130_fd_sc_hd__clkbuf_1 _11274_ (.A(_06893_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _11275_ (.A0(_05506_),
    .A1(\fifo_bank_register.bank[8][112] ),
    .S(_06891_),
    .X(_06894_));
 sky130_fd_sc_hd__clkbuf_1 _11276_ (.A(_06894_),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _11277_ (.A0(_05508_),
    .A1(\fifo_bank_register.bank[8][113] ),
    .S(_06891_),
    .X(_06895_));
 sky130_fd_sc_hd__clkbuf_1 _11278_ (.A(_06895_),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _11279_ (.A0(_05510_),
    .A1(\fifo_bank_register.bank[8][114] ),
    .S(_06891_),
    .X(_06896_));
 sky130_fd_sc_hd__clkbuf_1 _11280_ (.A(_06896_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _11281_ (.A0(_05512_),
    .A1(\fifo_bank_register.bank[8][115] ),
    .S(_06891_),
    .X(_06897_));
 sky130_fd_sc_hd__clkbuf_1 _11282_ (.A(_06897_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _11283_ (.A0(_05514_),
    .A1(\fifo_bank_register.bank[8][116] ),
    .S(_06891_),
    .X(_06898_));
 sky130_fd_sc_hd__clkbuf_1 _11284_ (.A(_06898_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _11285_ (.A0(_05516_),
    .A1(\fifo_bank_register.bank[8][117] ),
    .S(_06891_),
    .X(_06899_));
 sky130_fd_sc_hd__clkbuf_1 _11286_ (.A(_06899_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _11287_ (.A0(_05518_),
    .A1(\fifo_bank_register.bank[8][118] ),
    .S(_06891_),
    .X(_06900_));
 sky130_fd_sc_hd__clkbuf_1 _11288_ (.A(_06900_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(_05520_),
    .A1(\fifo_bank_register.bank[8][119] ),
    .S(_06891_),
    .X(_06901_));
 sky130_fd_sc_hd__clkbuf_1 _11290_ (.A(_06901_),
    .X(_00400_));
 sky130_fd_sc_hd__mux2_1 _11291_ (.A0(_05522_),
    .A1(\fifo_bank_register.bank[8][120] ),
    .S(_06768_),
    .X(_06902_));
 sky130_fd_sc_hd__clkbuf_1 _11292_ (.A(_06902_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _11293_ (.A0(_05524_),
    .A1(\fifo_bank_register.bank[8][121] ),
    .S(_06768_),
    .X(_06903_));
 sky130_fd_sc_hd__clkbuf_1 _11294_ (.A(_06903_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(_05526_),
    .A1(\fifo_bank_register.bank[8][122] ),
    .S(_06768_),
    .X(_06904_));
 sky130_fd_sc_hd__clkbuf_1 _11296_ (.A(_06904_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _11297_ (.A0(_05528_),
    .A1(\fifo_bank_register.bank[8][123] ),
    .S(_06768_),
    .X(_06905_));
 sky130_fd_sc_hd__clkbuf_1 _11298_ (.A(_06905_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _11299_ (.A0(_05530_),
    .A1(\fifo_bank_register.bank[8][124] ),
    .S(_06768_),
    .X(_06906_));
 sky130_fd_sc_hd__clkbuf_1 _11300_ (.A(_06906_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _11301_ (.A0(_05532_),
    .A1(\fifo_bank_register.bank[8][125] ),
    .S(_06768_),
    .X(_06907_));
 sky130_fd_sc_hd__clkbuf_1 _11302_ (.A(_06907_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _11303_ (.A0(_05534_),
    .A1(\fifo_bank_register.bank[8][126] ),
    .S(_06768_),
    .X(_06908_));
 sky130_fd_sc_hd__clkbuf_1 _11304_ (.A(_06908_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _11305_ (.A0(_05536_),
    .A1(\fifo_bank_register.bank[8][127] ),
    .S(_06768_),
    .X(_06909_));
 sky130_fd_sc_hd__clkbuf_1 _11306_ (.A(_06909_),
    .X(_00408_));
 sky130_fd_sc_hd__and3_1 _11307_ (.A(\fifo_bank_register.write_ptr[2] ),
    .B(_05254_),
    .C(_05266_),
    .X(_06910_));
 sky130_fd_sc_hd__and4_1 _11308_ (.A(net597),
    .B(_05249_),
    .C(_05250_),
    .D(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__buf_4 _11309_ (.A(_06911_),
    .X(_06912_));
 sky130_fd_sc_hd__buf_4 _11310_ (.A(_06912_),
    .X(_06913_));
 sky130_fd_sc_hd__mux2_1 _11311_ (.A0(\fifo_bank_register.bank[7][0] ),
    .A1(_05248_),
    .S(_06913_),
    .X(_06914_));
 sky130_fd_sc_hd__clkbuf_1 _11312_ (.A(_06914_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _11313_ (.A0(\fifo_bank_register.bank[7][1] ),
    .A1(_05272_),
    .S(_06913_),
    .X(_06915_));
 sky130_fd_sc_hd__clkbuf_1 _11314_ (.A(_06915_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _11315_ (.A0(\fifo_bank_register.bank[7][2] ),
    .A1(_05274_),
    .S(_06913_),
    .X(_06916_));
 sky130_fd_sc_hd__clkbuf_1 _11316_ (.A(_06916_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _11317_ (.A0(\fifo_bank_register.bank[7][3] ),
    .A1(_05276_),
    .S(_06913_),
    .X(_06917_));
 sky130_fd_sc_hd__clkbuf_1 _11318_ (.A(_06917_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _11319_ (.A0(\fifo_bank_register.bank[7][4] ),
    .A1(_05278_),
    .S(_06913_),
    .X(_06918_));
 sky130_fd_sc_hd__clkbuf_1 _11320_ (.A(_06918_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _11321_ (.A0(\fifo_bank_register.bank[7][5] ),
    .A1(_05280_),
    .S(_06913_),
    .X(_06919_));
 sky130_fd_sc_hd__clkbuf_1 _11322_ (.A(_06919_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _11323_ (.A0(\fifo_bank_register.bank[7][6] ),
    .A1(_05282_),
    .S(_06913_),
    .X(_06920_));
 sky130_fd_sc_hd__clkbuf_1 _11324_ (.A(_06920_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _11325_ (.A0(\fifo_bank_register.bank[7][7] ),
    .A1(_05284_),
    .S(_06913_),
    .X(_06921_));
 sky130_fd_sc_hd__clkbuf_1 _11326_ (.A(_06921_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _11327_ (.A0(\fifo_bank_register.bank[7][8] ),
    .A1(_05286_),
    .S(_06913_),
    .X(_06922_));
 sky130_fd_sc_hd__clkbuf_1 _11328_ (.A(_06922_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _11329_ (.A0(\fifo_bank_register.bank[7][9] ),
    .A1(_05288_),
    .S(_06913_),
    .X(_06923_));
 sky130_fd_sc_hd__clkbuf_1 _11330_ (.A(_06923_),
    .X(_00418_));
 sky130_fd_sc_hd__buf_4 _11331_ (.A(_06912_),
    .X(_06924_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(\fifo_bank_register.bank[7][10] ),
    .A1(_05290_),
    .S(_06924_),
    .X(_06925_));
 sky130_fd_sc_hd__clkbuf_1 _11333_ (.A(_06925_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _11334_ (.A0(\fifo_bank_register.bank[7][11] ),
    .A1(_05293_),
    .S(_06924_),
    .X(_06926_));
 sky130_fd_sc_hd__clkbuf_1 _11335_ (.A(_06926_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _11336_ (.A0(\fifo_bank_register.bank[7][12] ),
    .A1(_05295_),
    .S(_06924_),
    .X(_06927_));
 sky130_fd_sc_hd__clkbuf_1 _11337_ (.A(_06927_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _11338_ (.A0(\fifo_bank_register.bank[7][13] ),
    .A1(_05297_),
    .S(_06924_),
    .X(_06928_));
 sky130_fd_sc_hd__clkbuf_1 _11339_ (.A(_06928_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _11340_ (.A0(\fifo_bank_register.bank[7][14] ),
    .A1(_05299_),
    .S(_06924_),
    .X(_06929_));
 sky130_fd_sc_hd__clkbuf_1 _11341_ (.A(_06929_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _11342_ (.A0(\fifo_bank_register.bank[7][15] ),
    .A1(_05301_),
    .S(_06924_),
    .X(_06930_));
 sky130_fd_sc_hd__clkbuf_1 _11343_ (.A(_06930_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _11344_ (.A0(\fifo_bank_register.bank[7][16] ),
    .A1(_05303_),
    .S(_06924_),
    .X(_06931_));
 sky130_fd_sc_hd__clkbuf_1 _11345_ (.A(_06931_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _11346_ (.A0(\fifo_bank_register.bank[7][17] ),
    .A1(_05305_),
    .S(_06924_),
    .X(_06932_));
 sky130_fd_sc_hd__clkbuf_1 _11347_ (.A(_06932_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _11348_ (.A0(\fifo_bank_register.bank[7][18] ),
    .A1(_05307_),
    .S(_06924_),
    .X(_06933_));
 sky130_fd_sc_hd__clkbuf_1 _11349_ (.A(_06933_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _11350_ (.A0(\fifo_bank_register.bank[7][19] ),
    .A1(_05309_),
    .S(_06924_),
    .X(_06934_));
 sky130_fd_sc_hd__clkbuf_1 _11351_ (.A(_06934_),
    .X(_00428_));
 sky130_fd_sc_hd__buf_6 _11352_ (.A(_06911_),
    .X(_06935_));
 sky130_fd_sc_hd__buf_4 _11353_ (.A(_06935_),
    .X(_06936_));
 sky130_fd_sc_hd__mux2_1 _11354_ (.A0(\fifo_bank_register.bank[7][20] ),
    .A1(_05311_),
    .S(_06936_),
    .X(_06937_));
 sky130_fd_sc_hd__clkbuf_1 _11355_ (.A(_06937_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _11356_ (.A0(\fifo_bank_register.bank[7][21] ),
    .A1(_05315_),
    .S(_06936_),
    .X(_06938_));
 sky130_fd_sc_hd__clkbuf_1 _11357_ (.A(_06938_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _11358_ (.A0(\fifo_bank_register.bank[7][22] ),
    .A1(_05317_),
    .S(_06936_),
    .X(_06939_));
 sky130_fd_sc_hd__clkbuf_1 _11359_ (.A(_06939_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _11360_ (.A0(\fifo_bank_register.bank[7][23] ),
    .A1(_05319_),
    .S(_06936_),
    .X(_06940_));
 sky130_fd_sc_hd__clkbuf_1 _11361_ (.A(_06940_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _11362_ (.A0(\fifo_bank_register.bank[7][24] ),
    .A1(_05321_),
    .S(_06936_),
    .X(_06941_));
 sky130_fd_sc_hd__clkbuf_1 _11363_ (.A(_06941_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _11364_ (.A0(\fifo_bank_register.bank[7][25] ),
    .A1(_05323_),
    .S(_06936_),
    .X(_06942_));
 sky130_fd_sc_hd__clkbuf_1 _11365_ (.A(_06942_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _11366_ (.A0(\fifo_bank_register.bank[7][26] ),
    .A1(_05325_),
    .S(_06936_),
    .X(_06943_));
 sky130_fd_sc_hd__clkbuf_1 _11367_ (.A(_06943_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _11368_ (.A0(\fifo_bank_register.bank[7][27] ),
    .A1(_05327_),
    .S(_06936_),
    .X(_06944_));
 sky130_fd_sc_hd__clkbuf_1 _11369_ (.A(_06944_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _11370_ (.A0(\fifo_bank_register.bank[7][28] ),
    .A1(_05329_),
    .S(_06936_),
    .X(_06945_));
 sky130_fd_sc_hd__clkbuf_1 _11371_ (.A(_06945_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _11372_ (.A0(\fifo_bank_register.bank[7][29] ),
    .A1(_05331_),
    .S(_06936_),
    .X(_06946_));
 sky130_fd_sc_hd__clkbuf_1 _11373_ (.A(_06946_),
    .X(_00438_));
 sky130_fd_sc_hd__buf_4 _11374_ (.A(_06935_),
    .X(_06947_));
 sky130_fd_sc_hd__mux2_1 _11375_ (.A0(\fifo_bank_register.bank[7][30] ),
    .A1(_05333_),
    .S(_06947_),
    .X(_06948_));
 sky130_fd_sc_hd__clkbuf_1 _11376_ (.A(_06948_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _11377_ (.A0(\fifo_bank_register.bank[7][31] ),
    .A1(_05336_),
    .S(_06947_),
    .X(_06949_));
 sky130_fd_sc_hd__clkbuf_1 _11378_ (.A(_06949_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _11379_ (.A0(\fifo_bank_register.bank[7][32] ),
    .A1(_05338_),
    .S(_06947_),
    .X(_06950_));
 sky130_fd_sc_hd__clkbuf_1 _11380_ (.A(_06950_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _11381_ (.A0(\fifo_bank_register.bank[7][33] ),
    .A1(_05340_),
    .S(_06947_),
    .X(_06951_));
 sky130_fd_sc_hd__clkbuf_1 _11382_ (.A(_06951_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _11383_ (.A0(\fifo_bank_register.bank[7][34] ),
    .A1(_05342_),
    .S(_06947_),
    .X(_06952_));
 sky130_fd_sc_hd__clkbuf_1 _11384_ (.A(_06952_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _11385_ (.A0(\fifo_bank_register.bank[7][35] ),
    .A1(_05344_),
    .S(_06947_),
    .X(_06953_));
 sky130_fd_sc_hd__clkbuf_1 _11386_ (.A(_06953_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _11387_ (.A0(\fifo_bank_register.bank[7][36] ),
    .A1(_05346_),
    .S(_06947_),
    .X(_06954_));
 sky130_fd_sc_hd__clkbuf_1 _11388_ (.A(_06954_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _11389_ (.A0(\fifo_bank_register.bank[7][37] ),
    .A1(_05348_),
    .S(_06947_),
    .X(_06955_));
 sky130_fd_sc_hd__clkbuf_1 _11390_ (.A(_06955_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _11391_ (.A0(\fifo_bank_register.bank[7][38] ),
    .A1(_05350_),
    .S(_06947_),
    .X(_06956_));
 sky130_fd_sc_hd__clkbuf_1 _11392_ (.A(_06956_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _11393_ (.A0(\fifo_bank_register.bank[7][39] ),
    .A1(_05352_),
    .S(_06947_),
    .X(_06957_));
 sky130_fd_sc_hd__clkbuf_1 _11394_ (.A(_06957_),
    .X(_00448_));
 sky130_fd_sc_hd__buf_4 _11395_ (.A(_06935_),
    .X(_06958_));
 sky130_fd_sc_hd__mux2_1 _11396_ (.A0(\fifo_bank_register.bank[7][40] ),
    .A1(_05354_),
    .S(_06958_),
    .X(_06959_));
 sky130_fd_sc_hd__clkbuf_1 _11397_ (.A(_06959_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _11398_ (.A0(\fifo_bank_register.bank[7][41] ),
    .A1(_05357_),
    .S(_06958_),
    .X(_06960_));
 sky130_fd_sc_hd__clkbuf_1 _11399_ (.A(_06960_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _11400_ (.A0(\fifo_bank_register.bank[7][42] ),
    .A1(_05359_),
    .S(_06958_),
    .X(_06961_));
 sky130_fd_sc_hd__clkbuf_1 _11401_ (.A(_06961_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _11402_ (.A0(\fifo_bank_register.bank[7][43] ),
    .A1(_05361_),
    .S(_06958_),
    .X(_06962_));
 sky130_fd_sc_hd__clkbuf_1 _11403_ (.A(_06962_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _11404_ (.A0(\fifo_bank_register.bank[7][44] ),
    .A1(_05363_),
    .S(_06958_),
    .X(_06963_));
 sky130_fd_sc_hd__clkbuf_1 _11405_ (.A(_06963_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _11406_ (.A0(\fifo_bank_register.bank[7][45] ),
    .A1(_05365_),
    .S(_06958_),
    .X(_06964_));
 sky130_fd_sc_hd__clkbuf_1 _11407_ (.A(_06964_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _11408_ (.A0(\fifo_bank_register.bank[7][46] ),
    .A1(_05367_),
    .S(_06958_),
    .X(_06965_));
 sky130_fd_sc_hd__clkbuf_1 _11409_ (.A(_06965_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _11410_ (.A0(\fifo_bank_register.bank[7][47] ),
    .A1(_05369_),
    .S(_06958_),
    .X(_06966_));
 sky130_fd_sc_hd__clkbuf_1 _11411_ (.A(_06966_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _11412_ (.A0(\fifo_bank_register.bank[7][48] ),
    .A1(_05371_),
    .S(_06958_),
    .X(_06967_));
 sky130_fd_sc_hd__clkbuf_1 _11413_ (.A(_06967_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _11414_ (.A0(\fifo_bank_register.bank[7][49] ),
    .A1(_05373_),
    .S(_06958_),
    .X(_06968_));
 sky130_fd_sc_hd__clkbuf_1 _11415_ (.A(_06968_),
    .X(_00458_));
 sky130_fd_sc_hd__buf_4 _11416_ (.A(_06935_),
    .X(_06969_));
 sky130_fd_sc_hd__mux2_1 _11417_ (.A0(\fifo_bank_register.bank[7][50] ),
    .A1(_05375_),
    .S(_06969_),
    .X(_06970_));
 sky130_fd_sc_hd__clkbuf_1 _11418_ (.A(_06970_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _11419_ (.A0(\fifo_bank_register.bank[7][51] ),
    .A1(_05378_),
    .S(_06969_),
    .X(_06971_));
 sky130_fd_sc_hd__clkbuf_1 _11420_ (.A(_06971_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _11421_ (.A0(\fifo_bank_register.bank[7][52] ),
    .A1(_05380_),
    .S(_06969_),
    .X(_06972_));
 sky130_fd_sc_hd__clkbuf_1 _11422_ (.A(_06972_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _11423_ (.A0(\fifo_bank_register.bank[7][53] ),
    .A1(_05382_),
    .S(_06969_),
    .X(_06973_));
 sky130_fd_sc_hd__clkbuf_1 _11424_ (.A(_06973_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _11425_ (.A0(\fifo_bank_register.bank[7][54] ),
    .A1(_05384_),
    .S(_06969_),
    .X(_06974_));
 sky130_fd_sc_hd__clkbuf_1 _11426_ (.A(_06974_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _11427_ (.A0(\fifo_bank_register.bank[7][55] ),
    .A1(_05386_),
    .S(_06969_),
    .X(_06975_));
 sky130_fd_sc_hd__clkbuf_1 _11428_ (.A(_06975_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _11429_ (.A0(\fifo_bank_register.bank[7][56] ),
    .A1(_05388_),
    .S(_06969_),
    .X(_06976_));
 sky130_fd_sc_hd__clkbuf_1 _11430_ (.A(_06976_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _11431_ (.A0(\fifo_bank_register.bank[7][57] ),
    .A1(_05390_),
    .S(_06969_),
    .X(_06977_));
 sky130_fd_sc_hd__clkbuf_1 _11432_ (.A(_06977_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _11433_ (.A0(\fifo_bank_register.bank[7][58] ),
    .A1(_05392_),
    .S(_06969_),
    .X(_06978_));
 sky130_fd_sc_hd__clkbuf_1 _11434_ (.A(_06978_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _11435_ (.A0(\fifo_bank_register.bank[7][59] ),
    .A1(_05394_),
    .S(_06969_),
    .X(_06979_));
 sky130_fd_sc_hd__clkbuf_1 _11436_ (.A(_06979_),
    .X(_00468_));
 sky130_fd_sc_hd__buf_4 _11437_ (.A(_06935_),
    .X(_06980_));
 sky130_fd_sc_hd__mux2_1 _11438_ (.A0(\fifo_bank_register.bank[7][60] ),
    .A1(_05396_),
    .S(_06980_),
    .X(_06981_));
 sky130_fd_sc_hd__clkbuf_1 _11439_ (.A(_06981_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _11440_ (.A0(\fifo_bank_register.bank[7][61] ),
    .A1(_05399_),
    .S(_06980_),
    .X(_06982_));
 sky130_fd_sc_hd__clkbuf_1 _11441_ (.A(_06982_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _11442_ (.A0(\fifo_bank_register.bank[7][62] ),
    .A1(_05401_),
    .S(_06980_),
    .X(_06983_));
 sky130_fd_sc_hd__clkbuf_1 _11443_ (.A(_06983_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _11444_ (.A0(\fifo_bank_register.bank[7][63] ),
    .A1(_05403_),
    .S(_06980_),
    .X(_06984_));
 sky130_fd_sc_hd__clkbuf_1 _11445_ (.A(_06984_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _11446_ (.A0(\fifo_bank_register.bank[7][64] ),
    .A1(_05405_),
    .S(_06980_),
    .X(_06985_));
 sky130_fd_sc_hd__clkbuf_1 _11447_ (.A(_06985_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _11448_ (.A0(\fifo_bank_register.bank[7][65] ),
    .A1(_05407_),
    .S(_06980_),
    .X(_06986_));
 sky130_fd_sc_hd__clkbuf_1 _11449_ (.A(_06986_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _11450_ (.A0(\fifo_bank_register.bank[7][66] ),
    .A1(_05409_),
    .S(_06980_),
    .X(_06987_));
 sky130_fd_sc_hd__clkbuf_1 _11451_ (.A(_06987_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _11452_ (.A0(\fifo_bank_register.bank[7][67] ),
    .A1(_05411_),
    .S(_06980_),
    .X(_06988_));
 sky130_fd_sc_hd__clkbuf_1 _11453_ (.A(_06988_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _11454_ (.A0(\fifo_bank_register.bank[7][68] ),
    .A1(_05413_),
    .S(_06980_),
    .X(_06989_));
 sky130_fd_sc_hd__clkbuf_1 _11455_ (.A(_06989_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _11456_ (.A0(\fifo_bank_register.bank[7][69] ),
    .A1(_05415_),
    .S(_06980_),
    .X(_06990_));
 sky130_fd_sc_hd__clkbuf_1 _11457_ (.A(_06990_),
    .X(_00478_));
 sky130_fd_sc_hd__clkbuf_4 _11458_ (.A(_06935_),
    .X(_06991_));
 sky130_fd_sc_hd__mux2_1 _11459_ (.A0(\fifo_bank_register.bank[7][70] ),
    .A1(_05417_),
    .S(_06991_),
    .X(_06992_));
 sky130_fd_sc_hd__clkbuf_1 _11460_ (.A(_06992_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _11461_ (.A0(\fifo_bank_register.bank[7][71] ),
    .A1(_05420_),
    .S(_06991_),
    .X(_06993_));
 sky130_fd_sc_hd__clkbuf_1 _11462_ (.A(_06993_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _11463_ (.A0(\fifo_bank_register.bank[7][72] ),
    .A1(_05422_),
    .S(_06991_),
    .X(_06994_));
 sky130_fd_sc_hd__clkbuf_1 _11464_ (.A(_06994_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _11465_ (.A0(\fifo_bank_register.bank[7][73] ),
    .A1(_05424_),
    .S(_06991_),
    .X(_06995_));
 sky130_fd_sc_hd__clkbuf_1 _11466_ (.A(_06995_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _11467_ (.A0(\fifo_bank_register.bank[7][74] ),
    .A1(_05426_),
    .S(_06991_),
    .X(_06996_));
 sky130_fd_sc_hd__clkbuf_1 _11468_ (.A(_06996_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _11469_ (.A0(\fifo_bank_register.bank[7][75] ),
    .A1(_05428_),
    .S(_06991_),
    .X(_06997_));
 sky130_fd_sc_hd__clkbuf_1 _11470_ (.A(_06997_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _11471_ (.A0(\fifo_bank_register.bank[7][76] ),
    .A1(_05430_),
    .S(_06991_),
    .X(_06998_));
 sky130_fd_sc_hd__clkbuf_1 _11472_ (.A(_06998_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _11473_ (.A0(\fifo_bank_register.bank[7][77] ),
    .A1(_05432_),
    .S(_06991_),
    .X(_06999_));
 sky130_fd_sc_hd__clkbuf_1 _11474_ (.A(_06999_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _11475_ (.A0(\fifo_bank_register.bank[7][78] ),
    .A1(_05434_),
    .S(_06991_),
    .X(_07000_));
 sky130_fd_sc_hd__clkbuf_1 _11476_ (.A(_07000_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _11477_ (.A0(\fifo_bank_register.bank[7][79] ),
    .A1(_05436_),
    .S(_06991_),
    .X(_07001_));
 sky130_fd_sc_hd__clkbuf_1 _11478_ (.A(_07001_),
    .X(_00488_));
 sky130_fd_sc_hd__buf_4 _11479_ (.A(_06935_),
    .X(_07002_));
 sky130_fd_sc_hd__mux2_1 _11480_ (.A0(\fifo_bank_register.bank[7][80] ),
    .A1(_05438_),
    .S(_07002_),
    .X(_07003_));
 sky130_fd_sc_hd__clkbuf_1 _11481_ (.A(_07003_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _11482_ (.A0(\fifo_bank_register.bank[7][81] ),
    .A1(_05441_),
    .S(_07002_),
    .X(_07004_));
 sky130_fd_sc_hd__clkbuf_1 _11483_ (.A(_07004_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _11484_ (.A0(\fifo_bank_register.bank[7][82] ),
    .A1(_05443_),
    .S(_07002_),
    .X(_07005_));
 sky130_fd_sc_hd__clkbuf_1 _11485_ (.A(_07005_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _11486_ (.A0(\fifo_bank_register.bank[7][83] ),
    .A1(_05445_),
    .S(_07002_),
    .X(_07006_));
 sky130_fd_sc_hd__clkbuf_1 _11487_ (.A(_07006_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _11488_ (.A0(\fifo_bank_register.bank[7][84] ),
    .A1(_05447_),
    .S(_07002_),
    .X(_07007_));
 sky130_fd_sc_hd__clkbuf_1 _11489_ (.A(_07007_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _11490_ (.A0(\fifo_bank_register.bank[7][85] ),
    .A1(_05449_),
    .S(_07002_),
    .X(_07008_));
 sky130_fd_sc_hd__clkbuf_1 _11491_ (.A(_07008_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _11492_ (.A0(\fifo_bank_register.bank[7][86] ),
    .A1(_05451_),
    .S(_07002_),
    .X(_07009_));
 sky130_fd_sc_hd__clkbuf_1 _11493_ (.A(_07009_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _11494_ (.A0(\fifo_bank_register.bank[7][87] ),
    .A1(_05453_),
    .S(_07002_),
    .X(_07010_));
 sky130_fd_sc_hd__clkbuf_1 _11495_ (.A(_07010_),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _11496_ (.A0(\fifo_bank_register.bank[7][88] ),
    .A1(_05455_),
    .S(_07002_),
    .X(_07011_));
 sky130_fd_sc_hd__clkbuf_1 _11497_ (.A(_07011_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _11498_ (.A0(\fifo_bank_register.bank[7][89] ),
    .A1(_05457_),
    .S(_07002_),
    .X(_07012_));
 sky130_fd_sc_hd__clkbuf_1 _11499_ (.A(_07012_),
    .X(_00498_));
 sky130_fd_sc_hd__buf_4 _11500_ (.A(_06935_),
    .X(_07013_));
 sky130_fd_sc_hd__mux2_1 _11501_ (.A0(\fifo_bank_register.bank[7][90] ),
    .A1(_05459_),
    .S(_07013_),
    .X(_07014_));
 sky130_fd_sc_hd__clkbuf_1 _11502_ (.A(_07014_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _11503_ (.A0(\fifo_bank_register.bank[7][91] ),
    .A1(_05462_),
    .S(_07013_),
    .X(_07015_));
 sky130_fd_sc_hd__clkbuf_1 _11504_ (.A(_07015_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _11505_ (.A0(\fifo_bank_register.bank[7][92] ),
    .A1(_05464_),
    .S(_07013_),
    .X(_07016_));
 sky130_fd_sc_hd__clkbuf_1 _11506_ (.A(_07016_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _11507_ (.A0(\fifo_bank_register.bank[7][93] ),
    .A1(_05466_),
    .S(_07013_),
    .X(_07017_));
 sky130_fd_sc_hd__clkbuf_1 _11508_ (.A(_07017_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _11509_ (.A0(\fifo_bank_register.bank[7][94] ),
    .A1(_05468_),
    .S(_07013_),
    .X(_07018_));
 sky130_fd_sc_hd__clkbuf_1 _11510_ (.A(_07018_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _11511_ (.A0(\fifo_bank_register.bank[7][95] ),
    .A1(_05470_),
    .S(_07013_),
    .X(_07019_));
 sky130_fd_sc_hd__clkbuf_1 _11512_ (.A(_07019_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _11513_ (.A0(\fifo_bank_register.bank[7][96] ),
    .A1(_05472_),
    .S(_07013_),
    .X(_07020_));
 sky130_fd_sc_hd__clkbuf_1 _11514_ (.A(_07020_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(\fifo_bank_register.bank[7][97] ),
    .A1(_05474_),
    .S(_07013_),
    .X(_07021_));
 sky130_fd_sc_hd__clkbuf_1 _11516_ (.A(_07021_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _11517_ (.A0(\fifo_bank_register.bank[7][98] ),
    .A1(_05476_),
    .S(_07013_),
    .X(_07022_));
 sky130_fd_sc_hd__clkbuf_1 _11518_ (.A(_07022_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _11519_ (.A0(\fifo_bank_register.bank[7][99] ),
    .A1(_05478_),
    .S(_07013_),
    .X(_07023_));
 sky130_fd_sc_hd__clkbuf_1 _11520_ (.A(_07023_),
    .X(_00508_));
 sky130_fd_sc_hd__buf_4 _11521_ (.A(_06935_),
    .X(_07024_));
 sky130_fd_sc_hd__mux2_1 _11522_ (.A0(\fifo_bank_register.bank[7][100] ),
    .A1(_05480_),
    .S(_07024_),
    .X(_07025_));
 sky130_fd_sc_hd__clkbuf_1 _11523_ (.A(_07025_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _11524_ (.A0(\fifo_bank_register.bank[7][101] ),
    .A1(_05483_),
    .S(_07024_),
    .X(_07026_));
 sky130_fd_sc_hd__clkbuf_1 _11525_ (.A(_07026_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _11526_ (.A0(\fifo_bank_register.bank[7][102] ),
    .A1(_05485_),
    .S(_07024_),
    .X(_07027_));
 sky130_fd_sc_hd__clkbuf_1 _11527_ (.A(_07027_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _11528_ (.A0(\fifo_bank_register.bank[7][103] ),
    .A1(_05487_),
    .S(_07024_),
    .X(_07028_));
 sky130_fd_sc_hd__clkbuf_1 _11529_ (.A(_07028_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _11530_ (.A0(\fifo_bank_register.bank[7][104] ),
    .A1(_05489_),
    .S(_07024_),
    .X(_07029_));
 sky130_fd_sc_hd__clkbuf_1 _11531_ (.A(_07029_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _11532_ (.A0(\fifo_bank_register.bank[7][105] ),
    .A1(_05491_),
    .S(_07024_),
    .X(_07030_));
 sky130_fd_sc_hd__clkbuf_1 _11533_ (.A(_07030_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _11534_ (.A0(\fifo_bank_register.bank[7][106] ),
    .A1(_05493_),
    .S(_07024_),
    .X(_07031_));
 sky130_fd_sc_hd__clkbuf_1 _11535_ (.A(_07031_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _11536_ (.A0(\fifo_bank_register.bank[7][107] ),
    .A1(_05495_),
    .S(_07024_),
    .X(_07032_));
 sky130_fd_sc_hd__clkbuf_1 _11537_ (.A(_07032_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _11538_ (.A0(\fifo_bank_register.bank[7][108] ),
    .A1(_05497_),
    .S(_07024_),
    .X(_07033_));
 sky130_fd_sc_hd__clkbuf_1 _11539_ (.A(_07033_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _11540_ (.A0(\fifo_bank_register.bank[7][109] ),
    .A1(_05499_),
    .S(_07024_),
    .X(_07034_));
 sky130_fd_sc_hd__clkbuf_1 _11541_ (.A(_07034_),
    .X(_00518_));
 sky130_fd_sc_hd__buf_4 _11542_ (.A(_06935_),
    .X(_07035_));
 sky130_fd_sc_hd__mux2_1 _11543_ (.A0(\fifo_bank_register.bank[7][110] ),
    .A1(_05501_),
    .S(_07035_),
    .X(_07036_));
 sky130_fd_sc_hd__clkbuf_1 _11544_ (.A(_07036_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _11545_ (.A0(\fifo_bank_register.bank[7][111] ),
    .A1(_05504_),
    .S(_07035_),
    .X(_07037_));
 sky130_fd_sc_hd__clkbuf_1 _11546_ (.A(_07037_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _11547_ (.A0(\fifo_bank_register.bank[7][112] ),
    .A1(_05506_),
    .S(_07035_),
    .X(_07038_));
 sky130_fd_sc_hd__clkbuf_1 _11548_ (.A(_07038_),
    .X(_00521_));
 sky130_fd_sc_hd__mux2_1 _11549_ (.A0(\fifo_bank_register.bank[7][113] ),
    .A1(_05508_),
    .S(_07035_),
    .X(_07039_));
 sky130_fd_sc_hd__clkbuf_1 _11550_ (.A(_07039_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _11551_ (.A0(\fifo_bank_register.bank[7][114] ),
    .A1(_05510_),
    .S(_07035_),
    .X(_07040_));
 sky130_fd_sc_hd__clkbuf_1 _11552_ (.A(_07040_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _11553_ (.A0(\fifo_bank_register.bank[7][115] ),
    .A1(_05512_),
    .S(_07035_),
    .X(_07041_));
 sky130_fd_sc_hd__clkbuf_1 _11554_ (.A(_07041_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _11555_ (.A0(\fifo_bank_register.bank[7][116] ),
    .A1(_05514_),
    .S(_07035_),
    .X(_07042_));
 sky130_fd_sc_hd__clkbuf_1 _11556_ (.A(_07042_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _11557_ (.A0(\fifo_bank_register.bank[7][117] ),
    .A1(_05516_),
    .S(_07035_),
    .X(_07043_));
 sky130_fd_sc_hd__clkbuf_1 _11558_ (.A(_07043_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _11559_ (.A0(\fifo_bank_register.bank[7][118] ),
    .A1(_05518_),
    .S(_07035_),
    .X(_07044_));
 sky130_fd_sc_hd__clkbuf_1 _11560_ (.A(_07044_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _11561_ (.A0(\fifo_bank_register.bank[7][119] ),
    .A1(_05520_),
    .S(_07035_),
    .X(_07045_));
 sky130_fd_sc_hd__clkbuf_1 _11562_ (.A(_07045_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _11563_ (.A0(\fifo_bank_register.bank[7][120] ),
    .A1(_05522_),
    .S(_06912_),
    .X(_07046_));
 sky130_fd_sc_hd__clkbuf_1 _11564_ (.A(_07046_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _11565_ (.A0(\fifo_bank_register.bank[7][121] ),
    .A1(_05524_),
    .S(_06912_),
    .X(_07047_));
 sky130_fd_sc_hd__clkbuf_1 _11566_ (.A(_07047_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _11567_ (.A0(\fifo_bank_register.bank[7][122] ),
    .A1(_05526_),
    .S(_06912_),
    .X(_07048_));
 sky130_fd_sc_hd__clkbuf_1 _11568_ (.A(_07048_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _11569_ (.A0(\fifo_bank_register.bank[7][123] ),
    .A1(_05528_),
    .S(_06912_),
    .X(_07049_));
 sky130_fd_sc_hd__clkbuf_1 _11570_ (.A(_07049_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _11571_ (.A0(\fifo_bank_register.bank[7][124] ),
    .A1(_05530_),
    .S(_06912_),
    .X(_07050_));
 sky130_fd_sc_hd__clkbuf_1 _11572_ (.A(_07050_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _11573_ (.A0(\fifo_bank_register.bank[7][125] ),
    .A1(_05532_),
    .S(_06912_),
    .X(_07051_));
 sky130_fd_sc_hd__clkbuf_1 _11574_ (.A(_07051_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _11575_ (.A0(\fifo_bank_register.bank[7][126] ),
    .A1(_05534_),
    .S(_06912_),
    .X(_07052_));
 sky130_fd_sc_hd__clkbuf_1 _11576_ (.A(_07052_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _11577_ (.A0(\fifo_bank_register.bank[7][127] ),
    .A1(_05536_),
    .S(_06912_),
    .X(_07053_));
 sky130_fd_sc_hd__clkbuf_1 _11578_ (.A(_07053_),
    .X(_00536_));
 sky130_fd_sc_hd__and4b_1 _11579_ (.A_N(_05249_),
    .B(_05250_),
    .C(_06910_),
    .D(net597),
    .X(_07054_));
 sky130_fd_sc_hd__buf_4 _11580_ (.A(_07054_),
    .X(_07055_));
 sky130_fd_sc_hd__clkbuf_4 _11581_ (.A(_07055_),
    .X(_07056_));
 sky130_fd_sc_hd__mux2_1 _11582_ (.A0(\fifo_bank_register.bank[6][0] ),
    .A1(_05248_),
    .S(_07056_),
    .X(_07057_));
 sky130_fd_sc_hd__clkbuf_1 _11583_ (.A(_07057_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _11584_ (.A0(\fifo_bank_register.bank[6][1] ),
    .A1(_05272_),
    .S(_07056_),
    .X(_07058_));
 sky130_fd_sc_hd__clkbuf_1 _11585_ (.A(_07058_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _11586_ (.A0(\fifo_bank_register.bank[6][2] ),
    .A1(_05274_),
    .S(_07056_),
    .X(_07059_));
 sky130_fd_sc_hd__clkbuf_1 _11587_ (.A(_07059_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _11588_ (.A0(\fifo_bank_register.bank[6][3] ),
    .A1(_05276_),
    .S(_07056_),
    .X(_07060_));
 sky130_fd_sc_hd__clkbuf_1 _11589_ (.A(_07060_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _11590_ (.A0(\fifo_bank_register.bank[6][4] ),
    .A1(_05278_),
    .S(_07056_),
    .X(_07061_));
 sky130_fd_sc_hd__clkbuf_1 _11591_ (.A(_07061_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _11592_ (.A0(\fifo_bank_register.bank[6][5] ),
    .A1(_05280_),
    .S(_07056_),
    .X(_07062_));
 sky130_fd_sc_hd__clkbuf_1 _11593_ (.A(_07062_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _11594_ (.A0(\fifo_bank_register.bank[6][6] ),
    .A1(_05282_),
    .S(_07056_),
    .X(_07063_));
 sky130_fd_sc_hd__clkbuf_1 _11595_ (.A(_07063_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _11596_ (.A0(\fifo_bank_register.bank[6][7] ),
    .A1(_05284_),
    .S(_07056_),
    .X(_07064_));
 sky130_fd_sc_hd__clkbuf_1 _11597_ (.A(_07064_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _11598_ (.A0(\fifo_bank_register.bank[6][8] ),
    .A1(_05286_),
    .S(_07056_),
    .X(_07065_));
 sky130_fd_sc_hd__clkbuf_1 _11599_ (.A(_07065_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _11600_ (.A0(\fifo_bank_register.bank[6][9] ),
    .A1(_05288_),
    .S(_07056_),
    .X(_07066_));
 sky130_fd_sc_hd__clkbuf_1 _11601_ (.A(_07066_),
    .X(_00546_));
 sky130_fd_sc_hd__buf_4 _11602_ (.A(_07055_),
    .X(_07067_));
 sky130_fd_sc_hd__mux2_1 _11603_ (.A0(\fifo_bank_register.bank[6][10] ),
    .A1(_05290_),
    .S(_07067_),
    .X(_07068_));
 sky130_fd_sc_hd__clkbuf_1 _11604_ (.A(_07068_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _11605_ (.A0(\fifo_bank_register.bank[6][11] ),
    .A1(_05293_),
    .S(_07067_),
    .X(_07069_));
 sky130_fd_sc_hd__clkbuf_1 _11606_ (.A(_07069_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _11607_ (.A0(\fifo_bank_register.bank[6][12] ),
    .A1(_05295_),
    .S(_07067_),
    .X(_07070_));
 sky130_fd_sc_hd__clkbuf_1 _11608_ (.A(_07070_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _11609_ (.A0(\fifo_bank_register.bank[6][13] ),
    .A1(_05297_),
    .S(_07067_),
    .X(_07071_));
 sky130_fd_sc_hd__clkbuf_1 _11610_ (.A(_07071_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _11611_ (.A0(\fifo_bank_register.bank[6][14] ),
    .A1(_05299_),
    .S(_07067_),
    .X(_07072_));
 sky130_fd_sc_hd__clkbuf_1 _11612_ (.A(_07072_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _11613_ (.A0(\fifo_bank_register.bank[6][15] ),
    .A1(_05301_),
    .S(_07067_),
    .X(_07073_));
 sky130_fd_sc_hd__clkbuf_1 _11614_ (.A(_07073_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _11615_ (.A0(\fifo_bank_register.bank[6][16] ),
    .A1(_05303_),
    .S(_07067_),
    .X(_07074_));
 sky130_fd_sc_hd__clkbuf_1 _11616_ (.A(_07074_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _11617_ (.A0(\fifo_bank_register.bank[6][17] ),
    .A1(_05305_),
    .S(_07067_),
    .X(_07075_));
 sky130_fd_sc_hd__clkbuf_1 _11618_ (.A(_07075_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _11619_ (.A0(\fifo_bank_register.bank[6][18] ),
    .A1(_05307_),
    .S(_07067_),
    .X(_07076_));
 sky130_fd_sc_hd__clkbuf_1 _11620_ (.A(_07076_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _11621_ (.A0(\fifo_bank_register.bank[6][19] ),
    .A1(_05309_),
    .S(_07067_),
    .X(_07077_));
 sky130_fd_sc_hd__clkbuf_1 _11622_ (.A(_07077_),
    .X(_00556_));
 sky130_fd_sc_hd__buf_8 _11623_ (.A(_07054_),
    .X(_07078_));
 sky130_fd_sc_hd__buf_4 _11624_ (.A(_07078_),
    .X(_07079_));
 sky130_fd_sc_hd__mux2_1 _11625_ (.A0(\fifo_bank_register.bank[6][20] ),
    .A1(_05311_),
    .S(_07079_),
    .X(_07080_));
 sky130_fd_sc_hd__clkbuf_1 _11626_ (.A(_07080_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _11627_ (.A0(\fifo_bank_register.bank[6][21] ),
    .A1(_05315_),
    .S(_07079_),
    .X(_07081_));
 sky130_fd_sc_hd__clkbuf_1 _11628_ (.A(_07081_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _11629_ (.A0(\fifo_bank_register.bank[6][22] ),
    .A1(_05317_),
    .S(_07079_),
    .X(_07082_));
 sky130_fd_sc_hd__clkbuf_1 _11630_ (.A(_07082_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _11631_ (.A0(\fifo_bank_register.bank[6][23] ),
    .A1(_05319_),
    .S(_07079_),
    .X(_07083_));
 sky130_fd_sc_hd__clkbuf_1 _11632_ (.A(_07083_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _11633_ (.A0(\fifo_bank_register.bank[6][24] ),
    .A1(_05321_),
    .S(_07079_),
    .X(_07084_));
 sky130_fd_sc_hd__clkbuf_1 _11634_ (.A(_07084_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _11635_ (.A0(\fifo_bank_register.bank[6][25] ),
    .A1(_05323_),
    .S(_07079_),
    .X(_07085_));
 sky130_fd_sc_hd__clkbuf_1 _11636_ (.A(_07085_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _11637_ (.A0(\fifo_bank_register.bank[6][26] ),
    .A1(_05325_),
    .S(_07079_),
    .X(_07086_));
 sky130_fd_sc_hd__clkbuf_1 _11638_ (.A(_07086_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _11639_ (.A0(\fifo_bank_register.bank[6][27] ),
    .A1(_05327_),
    .S(_07079_),
    .X(_07087_));
 sky130_fd_sc_hd__clkbuf_1 _11640_ (.A(_07087_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _11641_ (.A0(\fifo_bank_register.bank[6][28] ),
    .A1(_05329_),
    .S(_07079_),
    .X(_07088_));
 sky130_fd_sc_hd__clkbuf_1 _11642_ (.A(_07088_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _11643_ (.A0(\fifo_bank_register.bank[6][29] ),
    .A1(_05331_),
    .S(_07079_),
    .X(_07089_));
 sky130_fd_sc_hd__clkbuf_1 _11644_ (.A(_07089_),
    .X(_00566_));
 sky130_fd_sc_hd__buf_4 _11645_ (.A(_07078_),
    .X(_07090_));
 sky130_fd_sc_hd__mux2_1 _11646_ (.A0(\fifo_bank_register.bank[6][30] ),
    .A1(_05333_),
    .S(_07090_),
    .X(_07091_));
 sky130_fd_sc_hd__clkbuf_1 _11647_ (.A(_07091_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _11648_ (.A0(\fifo_bank_register.bank[6][31] ),
    .A1(_05336_),
    .S(_07090_),
    .X(_07092_));
 sky130_fd_sc_hd__clkbuf_1 _11649_ (.A(_07092_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _11650_ (.A0(\fifo_bank_register.bank[6][32] ),
    .A1(_05338_),
    .S(_07090_),
    .X(_07093_));
 sky130_fd_sc_hd__clkbuf_1 _11651_ (.A(_07093_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _11652_ (.A0(\fifo_bank_register.bank[6][33] ),
    .A1(_05340_),
    .S(_07090_),
    .X(_07094_));
 sky130_fd_sc_hd__clkbuf_1 _11653_ (.A(_07094_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _11654_ (.A0(\fifo_bank_register.bank[6][34] ),
    .A1(_05342_),
    .S(_07090_),
    .X(_07095_));
 sky130_fd_sc_hd__clkbuf_1 _11655_ (.A(_07095_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _11656_ (.A0(\fifo_bank_register.bank[6][35] ),
    .A1(_05344_),
    .S(_07090_),
    .X(_07096_));
 sky130_fd_sc_hd__clkbuf_1 _11657_ (.A(_07096_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _11658_ (.A0(\fifo_bank_register.bank[6][36] ),
    .A1(_05346_),
    .S(_07090_),
    .X(_07097_));
 sky130_fd_sc_hd__clkbuf_1 _11659_ (.A(_07097_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _11660_ (.A0(\fifo_bank_register.bank[6][37] ),
    .A1(_05348_),
    .S(_07090_),
    .X(_07098_));
 sky130_fd_sc_hd__clkbuf_1 _11661_ (.A(_07098_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _11662_ (.A0(\fifo_bank_register.bank[6][38] ),
    .A1(_05350_),
    .S(_07090_),
    .X(_07099_));
 sky130_fd_sc_hd__clkbuf_1 _11663_ (.A(_07099_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(\fifo_bank_register.bank[6][39] ),
    .A1(_05352_),
    .S(_07090_),
    .X(_07100_));
 sky130_fd_sc_hd__clkbuf_1 _11665_ (.A(_07100_),
    .X(_00576_));
 sky130_fd_sc_hd__buf_4 _11666_ (.A(_07078_),
    .X(_07101_));
 sky130_fd_sc_hd__mux2_1 _11667_ (.A0(\fifo_bank_register.bank[6][40] ),
    .A1(_05354_),
    .S(_07101_),
    .X(_07102_));
 sky130_fd_sc_hd__clkbuf_1 _11668_ (.A(_07102_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _11669_ (.A0(\fifo_bank_register.bank[6][41] ),
    .A1(_05357_),
    .S(_07101_),
    .X(_07103_));
 sky130_fd_sc_hd__clkbuf_1 _11670_ (.A(_07103_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _11671_ (.A0(\fifo_bank_register.bank[6][42] ),
    .A1(_05359_),
    .S(_07101_),
    .X(_07104_));
 sky130_fd_sc_hd__clkbuf_1 _11672_ (.A(_07104_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _11673_ (.A0(\fifo_bank_register.bank[6][43] ),
    .A1(_05361_),
    .S(_07101_),
    .X(_07105_));
 sky130_fd_sc_hd__clkbuf_1 _11674_ (.A(_07105_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _11675_ (.A0(\fifo_bank_register.bank[6][44] ),
    .A1(_05363_),
    .S(_07101_),
    .X(_07106_));
 sky130_fd_sc_hd__clkbuf_1 _11676_ (.A(_07106_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _11677_ (.A0(\fifo_bank_register.bank[6][45] ),
    .A1(_05365_),
    .S(_07101_),
    .X(_07107_));
 sky130_fd_sc_hd__clkbuf_1 _11678_ (.A(_07107_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _11679_ (.A0(\fifo_bank_register.bank[6][46] ),
    .A1(_05367_),
    .S(_07101_),
    .X(_07108_));
 sky130_fd_sc_hd__clkbuf_1 _11680_ (.A(_07108_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _11681_ (.A0(\fifo_bank_register.bank[6][47] ),
    .A1(_05369_),
    .S(_07101_),
    .X(_07109_));
 sky130_fd_sc_hd__clkbuf_1 _11682_ (.A(_07109_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _11683_ (.A0(\fifo_bank_register.bank[6][48] ),
    .A1(_05371_),
    .S(_07101_),
    .X(_07110_));
 sky130_fd_sc_hd__clkbuf_1 _11684_ (.A(_07110_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _11685_ (.A0(\fifo_bank_register.bank[6][49] ),
    .A1(_05373_),
    .S(_07101_),
    .X(_07111_));
 sky130_fd_sc_hd__clkbuf_1 _11686_ (.A(_07111_),
    .X(_00586_));
 sky130_fd_sc_hd__buf_4 _11687_ (.A(_07078_),
    .X(_07112_));
 sky130_fd_sc_hd__mux2_1 _11688_ (.A0(\fifo_bank_register.bank[6][50] ),
    .A1(_05375_),
    .S(_07112_),
    .X(_07113_));
 sky130_fd_sc_hd__clkbuf_1 _11689_ (.A(_07113_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _11690_ (.A0(\fifo_bank_register.bank[6][51] ),
    .A1(_05378_),
    .S(_07112_),
    .X(_07114_));
 sky130_fd_sc_hd__clkbuf_1 _11691_ (.A(_07114_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _11692_ (.A0(\fifo_bank_register.bank[6][52] ),
    .A1(_05380_),
    .S(_07112_),
    .X(_07115_));
 sky130_fd_sc_hd__clkbuf_1 _11693_ (.A(_07115_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(\fifo_bank_register.bank[6][53] ),
    .A1(_05382_),
    .S(_07112_),
    .X(_07116_));
 sky130_fd_sc_hd__clkbuf_1 _11695_ (.A(_07116_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _11696_ (.A0(\fifo_bank_register.bank[6][54] ),
    .A1(_05384_),
    .S(_07112_),
    .X(_07117_));
 sky130_fd_sc_hd__clkbuf_1 _11697_ (.A(_07117_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _11698_ (.A0(\fifo_bank_register.bank[6][55] ),
    .A1(_05386_),
    .S(_07112_),
    .X(_07118_));
 sky130_fd_sc_hd__clkbuf_1 _11699_ (.A(_07118_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(\fifo_bank_register.bank[6][56] ),
    .A1(_05388_),
    .S(_07112_),
    .X(_07119_));
 sky130_fd_sc_hd__clkbuf_1 _11701_ (.A(_07119_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(\fifo_bank_register.bank[6][57] ),
    .A1(_05390_),
    .S(_07112_),
    .X(_07120_));
 sky130_fd_sc_hd__clkbuf_1 _11703_ (.A(_07120_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(\fifo_bank_register.bank[6][58] ),
    .A1(_05392_),
    .S(_07112_),
    .X(_07121_));
 sky130_fd_sc_hd__clkbuf_1 _11705_ (.A(_07121_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(\fifo_bank_register.bank[6][59] ),
    .A1(_05394_),
    .S(_07112_),
    .X(_07122_));
 sky130_fd_sc_hd__clkbuf_1 _11707_ (.A(_07122_),
    .X(_00596_));
 sky130_fd_sc_hd__buf_4 _11708_ (.A(_07078_),
    .X(_07123_));
 sky130_fd_sc_hd__mux2_1 _11709_ (.A0(\fifo_bank_register.bank[6][60] ),
    .A1(_05396_),
    .S(_07123_),
    .X(_07124_));
 sky130_fd_sc_hd__clkbuf_1 _11710_ (.A(_07124_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _11711_ (.A0(\fifo_bank_register.bank[6][61] ),
    .A1(_05399_),
    .S(_07123_),
    .X(_07125_));
 sky130_fd_sc_hd__clkbuf_1 _11712_ (.A(_07125_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _11713_ (.A0(\fifo_bank_register.bank[6][62] ),
    .A1(_05401_),
    .S(_07123_),
    .X(_07126_));
 sky130_fd_sc_hd__clkbuf_1 _11714_ (.A(_07126_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _11715_ (.A0(\fifo_bank_register.bank[6][63] ),
    .A1(_05403_),
    .S(_07123_),
    .X(_07127_));
 sky130_fd_sc_hd__clkbuf_1 _11716_ (.A(_07127_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _11717_ (.A0(\fifo_bank_register.bank[6][64] ),
    .A1(_05405_),
    .S(_07123_),
    .X(_07128_));
 sky130_fd_sc_hd__clkbuf_1 _11718_ (.A(_07128_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _11719_ (.A0(\fifo_bank_register.bank[6][65] ),
    .A1(_05407_),
    .S(_07123_),
    .X(_07129_));
 sky130_fd_sc_hd__clkbuf_1 _11720_ (.A(_07129_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _11721_ (.A0(\fifo_bank_register.bank[6][66] ),
    .A1(_05409_),
    .S(_07123_),
    .X(_07130_));
 sky130_fd_sc_hd__clkbuf_1 _11722_ (.A(_07130_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _11723_ (.A0(\fifo_bank_register.bank[6][67] ),
    .A1(_05411_),
    .S(_07123_),
    .X(_07131_));
 sky130_fd_sc_hd__clkbuf_1 _11724_ (.A(_07131_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _11725_ (.A0(\fifo_bank_register.bank[6][68] ),
    .A1(_05413_),
    .S(_07123_),
    .X(_07132_));
 sky130_fd_sc_hd__clkbuf_1 _11726_ (.A(_07132_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _11727_ (.A0(\fifo_bank_register.bank[6][69] ),
    .A1(_05415_),
    .S(_07123_),
    .X(_07133_));
 sky130_fd_sc_hd__clkbuf_1 _11728_ (.A(_07133_),
    .X(_00606_));
 sky130_fd_sc_hd__buf_4 _11729_ (.A(_07078_),
    .X(_07134_));
 sky130_fd_sc_hd__mux2_1 _11730_ (.A0(\fifo_bank_register.bank[6][70] ),
    .A1(_05417_),
    .S(_07134_),
    .X(_07135_));
 sky130_fd_sc_hd__clkbuf_1 _11731_ (.A(_07135_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _11732_ (.A0(\fifo_bank_register.bank[6][71] ),
    .A1(_05420_),
    .S(_07134_),
    .X(_07136_));
 sky130_fd_sc_hd__clkbuf_1 _11733_ (.A(_07136_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _11734_ (.A0(\fifo_bank_register.bank[6][72] ),
    .A1(_05422_),
    .S(_07134_),
    .X(_07137_));
 sky130_fd_sc_hd__clkbuf_1 _11735_ (.A(_07137_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(\fifo_bank_register.bank[6][73] ),
    .A1(_05424_),
    .S(_07134_),
    .X(_07138_));
 sky130_fd_sc_hd__clkbuf_1 _11737_ (.A(_07138_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _11738_ (.A0(\fifo_bank_register.bank[6][74] ),
    .A1(_05426_),
    .S(_07134_),
    .X(_07139_));
 sky130_fd_sc_hd__clkbuf_1 _11739_ (.A(_07139_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _11740_ (.A0(\fifo_bank_register.bank[6][75] ),
    .A1(_05428_),
    .S(_07134_),
    .X(_07140_));
 sky130_fd_sc_hd__clkbuf_1 _11741_ (.A(_07140_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _11742_ (.A0(\fifo_bank_register.bank[6][76] ),
    .A1(_05430_),
    .S(_07134_),
    .X(_07141_));
 sky130_fd_sc_hd__clkbuf_1 _11743_ (.A(_07141_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _11744_ (.A0(\fifo_bank_register.bank[6][77] ),
    .A1(_05432_),
    .S(_07134_),
    .X(_07142_));
 sky130_fd_sc_hd__clkbuf_1 _11745_ (.A(_07142_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _11746_ (.A0(\fifo_bank_register.bank[6][78] ),
    .A1(_05434_),
    .S(_07134_),
    .X(_07143_));
 sky130_fd_sc_hd__clkbuf_1 _11747_ (.A(_07143_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _11748_ (.A0(\fifo_bank_register.bank[6][79] ),
    .A1(_05436_),
    .S(_07134_),
    .X(_07144_));
 sky130_fd_sc_hd__clkbuf_1 _11749_ (.A(_07144_),
    .X(_00616_));
 sky130_fd_sc_hd__buf_4 _11750_ (.A(_07078_),
    .X(_07145_));
 sky130_fd_sc_hd__mux2_1 _11751_ (.A0(\fifo_bank_register.bank[6][80] ),
    .A1(_05438_),
    .S(_07145_),
    .X(_07146_));
 sky130_fd_sc_hd__clkbuf_1 _11752_ (.A(_07146_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _11753_ (.A0(\fifo_bank_register.bank[6][81] ),
    .A1(_05441_),
    .S(_07145_),
    .X(_07147_));
 sky130_fd_sc_hd__clkbuf_1 _11754_ (.A(_07147_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _11755_ (.A0(\fifo_bank_register.bank[6][82] ),
    .A1(_05443_),
    .S(_07145_),
    .X(_07148_));
 sky130_fd_sc_hd__clkbuf_1 _11756_ (.A(_07148_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _11757_ (.A0(\fifo_bank_register.bank[6][83] ),
    .A1(_05445_),
    .S(_07145_),
    .X(_07149_));
 sky130_fd_sc_hd__clkbuf_1 _11758_ (.A(_07149_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _11759_ (.A0(\fifo_bank_register.bank[6][84] ),
    .A1(_05447_),
    .S(_07145_),
    .X(_07150_));
 sky130_fd_sc_hd__clkbuf_1 _11760_ (.A(_07150_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _11761_ (.A0(\fifo_bank_register.bank[6][85] ),
    .A1(_05449_),
    .S(_07145_),
    .X(_07151_));
 sky130_fd_sc_hd__clkbuf_1 _11762_ (.A(_07151_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _11763_ (.A0(\fifo_bank_register.bank[6][86] ),
    .A1(_05451_),
    .S(_07145_),
    .X(_07152_));
 sky130_fd_sc_hd__clkbuf_1 _11764_ (.A(_07152_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _11765_ (.A0(\fifo_bank_register.bank[6][87] ),
    .A1(_05453_),
    .S(_07145_),
    .X(_07153_));
 sky130_fd_sc_hd__clkbuf_1 _11766_ (.A(_07153_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _11767_ (.A0(\fifo_bank_register.bank[6][88] ),
    .A1(_05455_),
    .S(_07145_),
    .X(_07154_));
 sky130_fd_sc_hd__clkbuf_1 _11768_ (.A(_07154_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _11769_ (.A0(\fifo_bank_register.bank[6][89] ),
    .A1(_05457_),
    .S(_07145_),
    .X(_07155_));
 sky130_fd_sc_hd__clkbuf_1 _11770_ (.A(_07155_),
    .X(_00626_));
 sky130_fd_sc_hd__buf_4 _11771_ (.A(_07078_),
    .X(_07156_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(\fifo_bank_register.bank[6][90] ),
    .A1(_05459_),
    .S(_07156_),
    .X(_07157_));
 sky130_fd_sc_hd__clkbuf_1 _11773_ (.A(_07157_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _11774_ (.A0(\fifo_bank_register.bank[6][91] ),
    .A1(_05462_),
    .S(_07156_),
    .X(_07158_));
 sky130_fd_sc_hd__clkbuf_1 _11775_ (.A(_07158_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _11776_ (.A0(\fifo_bank_register.bank[6][92] ),
    .A1(_05464_),
    .S(_07156_),
    .X(_07159_));
 sky130_fd_sc_hd__clkbuf_1 _11777_ (.A(_07159_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _11778_ (.A0(\fifo_bank_register.bank[6][93] ),
    .A1(_05466_),
    .S(_07156_),
    .X(_07160_));
 sky130_fd_sc_hd__clkbuf_1 _11779_ (.A(_07160_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _11780_ (.A0(\fifo_bank_register.bank[6][94] ),
    .A1(_05468_),
    .S(_07156_),
    .X(_07161_));
 sky130_fd_sc_hd__clkbuf_1 _11781_ (.A(_07161_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _11782_ (.A0(\fifo_bank_register.bank[6][95] ),
    .A1(_05470_),
    .S(_07156_),
    .X(_07162_));
 sky130_fd_sc_hd__clkbuf_1 _11783_ (.A(_07162_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _11784_ (.A0(\fifo_bank_register.bank[6][96] ),
    .A1(_05472_),
    .S(_07156_),
    .X(_07163_));
 sky130_fd_sc_hd__clkbuf_1 _11785_ (.A(_07163_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _11786_ (.A0(\fifo_bank_register.bank[6][97] ),
    .A1(_05474_),
    .S(_07156_),
    .X(_07164_));
 sky130_fd_sc_hd__clkbuf_1 _11787_ (.A(_07164_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _11788_ (.A0(\fifo_bank_register.bank[6][98] ),
    .A1(_05476_),
    .S(_07156_),
    .X(_07165_));
 sky130_fd_sc_hd__clkbuf_1 _11789_ (.A(_07165_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _11790_ (.A0(\fifo_bank_register.bank[6][99] ),
    .A1(_05478_),
    .S(_07156_),
    .X(_07166_));
 sky130_fd_sc_hd__clkbuf_1 _11791_ (.A(_07166_),
    .X(_00636_));
 sky130_fd_sc_hd__buf_4 _11792_ (.A(_07078_),
    .X(_07167_));
 sky130_fd_sc_hd__mux2_1 _11793_ (.A0(\fifo_bank_register.bank[6][100] ),
    .A1(_05480_),
    .S(_07167_),
    .X(_07168_));
 sky130_fd_sc_hd__clkbuf_1 _11794_ (.A(_07168_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _11795_ (.A0(\fifo_bank_register.bank[6][101] ),
    .A1(_05483_),
    .S(_07167_),
    .X(_07169_));
 sky130_fd_sc_hd__clkbuf_1 _11796_ (.A(_07169_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _11797_ (.A0(\fifo_bank_register.bank[6][102] ),
    .A1(_05485_),
    .S(_07167_),
    .X(_07170_));
 sky130_fd_sc_hd__clkbuf_1 _11798_ (.A(_07170_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _11799_ (.A0(\fifo_bank_register.bank[6][103] ),
    .A1(_05487_),
    .S(_07167_),
    .X(_07171_));
 sky130_fd_sc_hd__clkbuf_1 _11800_ (.A(_07171_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _11801_ (.A0(\fifo_bank_register.bank[6][104] ),
    .A1(_05489_),
    .S(_07167_),
    .X(_07172_));
 sky130_fd_sc_hd__clkbuf_1 _11802_ (.A(_07172_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _11803_ (.A0(\fifo_bank_register.bank[6][105] ),
    .A1(_05491_),
    .S(_07167_),
    .X(_07173_));
 sky130_fd_sc_hd__clkbuf_1 _11804_ (.A(_07173_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _11805_ (.A0(\fifo_bank_register.bank[6][106] ),
    .A1(_05493_),
    .S(_07167_),
    .X(_07174_));
 sky130_fd_sc_hd__clkbuf_1 _11806_ (.A(_07174_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _11807_ (.A0(\fifo_bank_register.bank[6][107] ),
    .A1(_05495_),
    .S(_07167_),
    .X(_07175_));
 sky130_fd_sc_hd__clkbuf_1 _11808_ (.A(_07175_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _11809_ (.A0(\fifo_bank_register.bank[6][108] ),
    .A1(_05497_),
    .S(_07167_),
    .X(_07176_));
 sky130_fd_sc_hd__clkbuf_1 _11810_ (.A(_07176_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _11811_ (.A0(\fifo_bank_register.bank[6][109] ),
    .A1(_05499_),
    .S(_07167_),
    .X(_07177_));
 sky130_fd_sc_hd__clkbuf_1 _11812_ (.A(_07177_),
    .X(_00646_));
 sky130_fd_sc_hd__buf_4 _11813_ (.A(_07078_),
    .X(_07178_));
 sky130_fd_sc_hd__mux2_1 _11814_ (.A0(\fifo_bank_register.bank[6][110] ),
    .A1(_05501_),
    .S(_07178_),
    .X(_07179_));
 sky130_fd_sc_hd__clkbuf_1 _11815_ (.A(_07179_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _11816_ (.A0(\fifo_bank_register.bank[6][111] ),
    .A1(_05504_),
    .S(_07178_),
    .X(_07180_));
 sky130_fd_sc_hd__clkbuf_1 _11817_ (.A(_07180_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _11818_ (.A0(\fifo_bank_register.bank[6][112] ),
    .A1(_05506_),
    .S(_07178_),
    .X(_07181_));
 sky130_fd_sc_hd__clkbuf_1 _11819_ (.A(_07181_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _11820_ (.A0(\fifo_bank_register.bank[6][113] ),
    .A1(_05508_),
    .S(_07178_),
    .X(_07182_));
 sky130_fd_sc_hd__clkbuf_1 _11821_ (.A(_07182_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _11822_ (.A0(\fifo_bank_register.bank[6][114] ),
    .A1(_05510_),
    .S(_07178_),
    .X(_07183_));
 sky130_fd_sc_hd__clkbuf_1 _11823_ (.A(_07183_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _11824_ (.A0(\fifo_bank_register.bank[6][115] ),
    .A1(_05512_),
    .S(_07178_),
    .X(_07184_));
 sky130_fd_sc_hd__clkbuf_1 _11825_ (.A(_07184_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _11826_ (.A0(\fifo_bank_register.bank[6][116] ),
    .A1(_05514_),
    .S(_07178_),
    .X(_07185_));
 sky130_fd_sc_hd__clkbuf_1 _11827_ (.A(_07185_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _11828_ (.A0(\fifo_bank_register.bank[6][117] ),
    .A1(_05516_),
    .S(_07178_),
    .X(_07186_));
 sky130_fd_sc_hd__clkbuf_1 _11829_ (.A(_07186_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _11830_ (.A0(\fifo_bank_register.bank[6][118] ),
    .A1(_05518_),
    .S(_07178_),
    .X(_07187_));
 sky130_fd_sc_hd__clkbuf_1 _11831_ (.A(_07187_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _11832_ (.A0(\fifo_bank_register.bank[6][119] ),
    .A1(_05520_),
    .S(_07178_),
    .X(_07188_));
 sky130_fd_sc_hd__clkbuf_1 _11833_ (.A(_07188_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _11834_ (.A0(\fifo_bank_register.bank[6][120] ),
    .A1(_05522_),
    .S(_07055_),
    .X(_07189_));
 sky130_fd_sc_hd__clkbuf_1 _11835_ (.A(_07189_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _11836_ (.A0(\fifo_bank_register.bank[6][121] ),
    .A1(_05524_),
    .S(_07055_),
    .X(_07190_));
 sky130_fd_sc_hd__clkbuf_1 _11837_ (.A(_07190_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _11838_ (.A0(\fifo_bank_register.bank[6][122] ),
    .A1(_05526_),
    .S(_07055_),
    .X(_07191_));
 sky130_fd_sc_hd__clkbuf_1 _11839_ (.A(_07191_),
    .X(_00659_));
 sky130_fd_sc_hd__mux2_1 _11840_ (.A0(\fifo_bank_register.bank[6][123] ),
    .A1(_05528_),
    .S(_07055_),
    .X(_07192_));
 sky130_fd_sc_hd__clkbuf_1 _11841_ (.A(_07192_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(\fifo_bank_register.bank[6][124] ),
    .A1(_05530_),
    .S(_07055_),
    .X(_07193_));
 sky130_fd_sc_hd__clkbuf_1 _11843_ (.A(_07193_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _11844_ (.A0(\fifo_bank_register.bank[6][125] ),
    .A1(_05532_),
    .S(_07055_),
    .X(_07194_));
 sky130_fd_sc_hd__clkbuf_1 _11845_ (.A(_07194_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(\fifo_bank_register.bank[6][126] ),
    .A1(_05534_),
    .S(_07055_),
    .X(_07195_));
 sky130_fd_sc_hd__clkbuf_1 _11847_ (.A(_07195_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _11848_ (.A0(\fifo_bank_register.bank[6][127] ),
    .A1(_05536_),
    .S(_07055_),
    .X(_07196_));
 sky130_fd_sc_hd__clkbuf_1 _11849_ (.A(_07196_),
    .X(_00664_));
 sky130_fd_sc_hd__and2_1 _11850_ (.A(_05267_),
    .B(_06910_),
    .X(_07197_));
 sky130_fd_sc_hd__clkbuf_4 _11851_ (.A(_07197_),
    .X(_07198_));
 sky130_fd_sc_hd__buf_4 _11852_ (.A(_07198_),
    .X(_07199_));
 sky130_fd_sc_hd__mux2_1 _11853_ (.A0(\fifo_bank_register.bank[5][0] ),
    .A1(_05248_),
    .S(_07199_),
    .X(_07200_));
 sky130_fd_sc_hd__clkbuf_1 _11854_ (.A(_07200_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _11855_ (.A0(\fifo_bank_register.bank[5][1] ),
    .A1(_05272_),
    .S(_07199_),
    .X(_07201_));
 sky130_fd_sc_hd__clkbuf_1 _11856_ (.A(_07201_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _11857_ (.A0(\fifo_bank_register.bank[5][2] ),
    .A1(_05274_),
    .S(_07199_),
    .X(_07202_));
 sky130_fd_sc_hd__clkbuf_1 _11858_ (.A(_07202_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _11859_ (.A0(\fifo_bank_register.bank[5][3] ),
    .A1(_05276_),
    .S(_07199_),
    .X(_07203_));
 sky130_fd_sc_hd__clkbuf_1 _11860_ (.A(_07203_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _11861_ (.A0(\fifo_bank_register.bank[5][4] ),
    .A1(_05278_),
    .S(_07199_),
    .X(_07204_));
 sky130_fd_sc_hd__clkbuf_1 _11862_ (.A(_07204_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _11863_ (.A0(\fifo_bank_register.bank[5][5] ),
    .A1(_05280_),
    .S(_07199_),
    .X(_07205_));
 sky130_fd_sc_hd__clkbuf_1 _11864_ (.A(_07205_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(\fifo_bank_register.bank[5][6] ),
    .A1(_05282_),
    .S(_07199_),
    .X(_07206_));
 sky130_fd_sc_hd__clkbuf_1 _11866_ (.A(_07206_),
    .X(_00671_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(\fifo_bank_register.bank[5][7] ),
    .A1(_05284_),
    .S(_07199_),
    .X(_07207_));
 sky130_fd_sc_hd__clkbuf_1 _11868_ (.A(_07207_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(\fifo_bank_register.bank[5][8] ),
    .A1(_05286_),
    .S(_07199_),
    .X(_07208_));
 sky130_fd_sc_hd__clkbuf_1 _11870_ (.A(_07208_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _11871_ (.A0(\fifo_bank_register.bank[5][9] ),
    .A1(_05288_),
    .S(_07199_),
    .X(_07209_));
 sky130_fd_sc_hd__clkbuf_1 _11872_ (.A(_07209_),
    .X(_00674_));
 sky130_fd_sc_hd__buf_4 _11873_ (.A(_07198_),
    .X(_07210_));
 sky130_fd_sc_hd__mux2_1 _11874_ (.A0(\fifo_bank_register.bank[5][10] ),
    .A1(_05290_),
    .S(_07210_),
    .X(_07211_));
 sky130_fd_sc_hd__clkbuf_1 _11875_ (.A(_07211_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _11876_ (.A0(\fifo_bank_register.bank[5][11] ),
    .A1(_05293_),
    .S(_07210_),
    .X(_07212_));
 sky130_fd_sc_hd__clkbuf_1 _11877_ (.A(_07212_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _11878_ (.A0(\fifo_bank_register.bank[5][12] ),
    .A1(_05295_),
    .S(_07210_),
    .X(_07213_));
 sky130_fd_sc_hd__clkbuf_1 _11879_ (.A(_07213_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _11880_ (.A0(\fifo_bank_register.bank[5][13] ),
    .A1(_05297_),
    .S(_07210_),
    .X(_07214_));
 sky130_fd_sc_hd__clkbuf_1 _11881_ (.A(_07214_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _11882_ (.A0(\fifo_bank_register.bank[5][14] ),
    .A1(_05299_),
    .S(_07210_),
    .X(_07215_));
 sky130_fd_sc_hd__clkbuf_1 _11883_ (.A(_07215_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _11884_ (.A0(\fifo_bank_register.bank[5][15] ),
    .A1(_05301_),
    .S(_07210_),
    .X(_07216_));
 sky130_fd_sc_hd__clkbuf_1 _11885_ (.A(_07216_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _11886_ (.A0(\fifo_bank_register.bank[5][16] ),
    .A1(_05303_),
    .S(_07210_),
    .X(_07217_));
 sky130_fd_sc_hd__clkbuf_1 _11887_ (.A(_07217_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _11888_ (.A0(\fifo_bank_register.bank[5][17] ),
    .A1(_05305_),
    .S(_07210_),
    .X(_07218_));
 sky130_fd_sc_hd__clkbuf_1 _11889_ (.A(_07218_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _11890_ (.A0(\fifo_bank_register.bank[5][18] ),
    .A1(_05307_),
    .S(_07210_),
    .X(_07219_));
 sky130_fd_sc_hd__clkbuf_1 _11891_ (.A(_07219_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _11892_ (.A0(\fifo_bank_register.bank[5][19] ),
    .A1(_05309_),
    .S(_07210_),
    .X(_07220_));
 sky130_fd_sc_hd__clkbuf_1 _11893_ (.A(_07220_),
    .X(_00684_));
 sky130_fd_sc_hd__buf_8 _11894_ (.A(_07197_),
    .X(_07221_));
 sky130_fd_sc_hd__clkbuf_4 _11895_ (.A(_07221_),
    .X(_07222_));
 sky130_fd_sc_hd__mux2_1 _11896_ (.A0(\fifo_bank_register.bank[5][20] ),
    .A1(_05311_),
    .S(_07222_),
    .X(_07223_));
 sky130_fd_sc_hd__clkbuf_1 _11897_ (.A(_07223_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _11898_ (.A0(\fifo_bank_register.bank[5][21] ),
    .A1(_05315_),
    .S(_07222_),
    .X(_07224_));
 sky130_fd_sc_hd__clkbuf_1 _11899_ (.A(_07224_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _11900_ (.A0(\fifo_bank_register.bank[5][22] ),
    .A1(_05317_),
    .S(_07222_),
    .X(_07225_));
 sky130_fd_sc_hd__clkbuf_1 _11901_ (.A(_07225_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _11902_ (.A0(\fifo_bank_register.bank[5][23] ),
    .A1(_05319_),
    .S(_07222_),
    .X(_07226_));
 sky130_fd_sc_hd__clkbuf_1 _11903_ (.A(_07226_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _11904_ (.A0(\fifo_bank_register.bank[5][24] ),
    .A1(_05321_),
    .S(_07222_),
    .X(_07227_));
 sky130_fd_sc_hd__clkbuf_1 _11905_ (.A(_07227_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _11906_ (.A0(\fifo_bank_register.bank[5][25] ),
    .A1(_05323_),
    .S(_07222_),
    .X(_07228_));
 sky130_fd_sc_hd__clkbuf_1 _11907_ (.A(_07228_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _11908_ (.A0(\fifo_bank_register.bank[5][26] ),
    .A1(_05325_),
    .S(_07222_),
    .X(_07229_));
 sky130_fd_sc_hd__clkbuf_1 _11909_ (.A(_07229_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _11910_ (.A0(\fifo_bank_register.bank[5][27] ),
    .A1(_05327_),
    .S(_07222_),
    .X(_07230_));
 sky130_fd_sc_hd__clkbuf_1 _11911_ (.A(_07230_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _11912_ (.A0(\fifo_bank_register.bank[5][28] ),
    .A1(_05329_),
    .S(_07222_),
    .X(_07231_));
 sky130_fd_sc_hd__clkbuf_1 _11913_ (.A(_07231_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _11914_ (.A0(\fifo_bank_register.bank[5][29] ),
    .A1(_05331_),
    .S(_07222_),
    .X(_07232_));
 sky130_fd_sc_hd__clkbuf_1 _11915_ (.A(_07232_),
    .X(_00694_));
 sky130_fd_sc_hd__buf_4 _11916_ (.A(_07221_),
    .X(_07233_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(\fifo_bank_register.bank[5][30] ),
    .A1(_05333_),
    .S(_07233_),
    .X(_07234_));
 sky130_fd_sc_hd__clkbuf_1 _11918_ (.A(_07234_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _11919_ (.A0(\fifo_bank_register.bank[5][31] ),
    .A1(_05336_),
    .S(_07233_),
    .X(_07235_));
 sky130_fd_sc_hd__clkbuf_1 _11920_ (.A(_07235_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _11921_ (.A0(\fifo_bank_register.bank[5][32] ),
    .A1(_05338_),
    .S(_07233_),
    .X(_07236_));
 sky130_fd_sc_hd__clkbuf_1 _11922_ (.A(_07236_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _11923_ (.A0(\fifo_bank_register.bank[5][33] ),
    .A1(_05340_),
    .S(_07233_),
    .X(_07237_));
 sky130_fd_sc_hd__clkbuf_1 _11924_ (.A(_07237_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _11925_ (.A0(\fifo_bank_register.bank[5][34] ),
    .A1(_05342_),
    .S(_07233_),
    .X(_07238_));
 sky130_fd_sc_hd__clkbuf_1 _11926_ (.A(_07238_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _11927_ (.A0(\fifo_bank_register.bank[5][35] ),
    .A1(_05344_),
    .S(_07233_),
    .X(_07239_));
 sky130_fd_sc_hd__clkbuf_1 _11928_ (.A(_07239_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _11929_ (.A0(\fifo_bank_register.bank[5][36] ),
    .A1(_05346_),
    .S(_07233_),
    .X(_07240_));
 sky130_fd_sc_hd__clkbuf_1 _11930_ (.A(_07240_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _11931_ (.A0(\fifo_bank_register.bank[5][37] ),
    .A1(_05348_),
    .S(_07233_),
    .X(_07241_));
 sky130_fd_sc_hd__clkbuf_1 _11932_ (.A(_07241_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _11933_ (.A0(\fifo_bank_register.bank[5][38] ),
    .A1(_05350_),
    .S(_07233_),
    .X(_07242_));
 sky130_fd_sc_hd__clkbuf_1 _11934_ (.A(_07242_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _11935_ (.A0(\fifo_bank_register.bank[5][39] ),
    .A1(_05352_),
    .S(_07233_),
    .X(_07243_));
 sky130_fd_sc_hd__clkbuf_1 _11936_ (.A(_07243_),
    .X(_00704_));
 sky130_fd_sc_hd__buf_4 _11937_ (.A(_07221_),
    .X(_07244_));
 sky130_fd_sc_hd__mux2_1 _11938_ (.A0(\fifo_bank_register.bank[5][40] ),
    .A1(_05354_),
    .S(_07244_),
    .X(_07245_));
 sky130_fd_sc_hd__clkbuf_1 _11939_ (.A(_07245_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _11940_ (.A0(\fifo_bank_register.bank[5][41] ),
    .A1(_05357_),
    .S(_07244_),
    .X(_07246_));
 sky130_fd_sc_hd__clkbuf_1 _11941_ (.A(_07246_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _11942_ (.A0(\fifo_bank_register.bank[5][42] ),
    .A1(_05359_),
    .S(_07244_),
    .X(_07247_));
 sky130_fd_sc_hd__clkbuf_1 _11943_ (.A(_07247_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _11944_ (.A0(\fifo_bank_register.bank[5][43] ),
    .A1(_05361_),
    .S(_07244_),
    .X(_07248_));
 sky130_fd_sc_hd__clkbuf_1 _11945_ (.A(_07248_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _11946_ (.A0(\fifo_bank_register.bank[5][44] ),
    .A1(_05363_),
    .S(_07244_),
    .X(_07249_));
 sky130_fd_sc_hd__clkbuf_1 _11947_ (.A(_07249_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _11948_ (.A0(\fifo_bank_register.bank[5][45] ),
    .A1(_05365_),
    .S(_07244_),
    .X(_07250_));
 sky130_fd_sc_hd__clkbuf_1 _11949_ (.A(_07250_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _11950_ (.A0(\fifo_bank_register.bank[5][46] ),
    .A1(_05367_),
    .S(_07244_),
    .X(_07251_));
 sky130_fd_sc_hd__clkbuf_1 _11951_ (.A(_07251_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _11952_ (.A0(\fifo_bank_register.bank[5][47] ),
    .A1(_05369_),
    .S(_07244_),
    .X(_07252_));
 sky130_fd_sc_hd__clkbuf_1 _11953_ (.A(_07252_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _11954_ (.A0(\fifo_bank_register.bank[5][48] ),
    .A1(_05371_),
    .S(_07244_),
    .X(_07253_));
 sky130_fd_sc_hd__clkbuf_1 _11955_ (.A(_07253_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _11956_ (.A0(\fifo_bank_register.bank[5][49] ),
    .A1(_05373_),
    .S(_07244_),
    .X(_07254_));
 sky130_fd_sc_hd__clkbuf_1 _11957_ (.A(_07254_),
    .X(_00714_));
 sky130_fd_sc_hd__buf_4 _11958_ (.A(_07221_),
    .X(_07255_));
 sky130_fd_sc_hd__mux2_1 _11959_ (.A0(\fifo_bank_register.bank[5][50] ),
    .A1(_05375_),
    .S(_07255_),
    .X(_07256_));
 sky130_fd_sc_hd__clkbuf_1 _11960_ (.A(_07256_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _11961_ (.A0(\fifo_bank_register.bank[5][51] ),
    .A1(_05378_),
    .S(_07255_),
    .X(_07257_));
 sky130_fd_sc_hd__clkbuf_1 _11962_ (.A(_07257_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _11963_ (.A0(\fifo_bank_register.bank[5][52] ),
    .A1(_05380_),
    .S(_07255_),
    .X(_07258_));
 sky130_fd_sc_hd__clkbuf_1 _11964_ (.A(_07258_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _11965_ (.A0(\fifo_bank_register.bank[5][53] ),
    .A1(_05382_),
    .S(_07255_),
    .X(_07259_));
 sky130_fd_sc_hd__clkbuf_1 _11966_ (.A(_07259_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _11967_ (.A0(\fifo_bank_register.bank[5][54] ),
    .A1(_05384_),
    .S(_07255_),
    .X(_07260_));
 sky130_fd_sc_hd__clkbuf_1 _11968_ (.A(_07260_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _11969_ (.A0(\fifo_bank_register.bank[5][55] ),
    .A1(_05386_),
    .S(_07255_),
    .X(_07261_));
 sky130_fd_sc_hd__clkbuf_1 _11970_ (.A(_07261_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _11971_ (.A0(\fifo_bank_register.bank[5][56] ),
    .A1(_05388_),
    .S(_07255_),
    .X(_07262_));
 sky130_fd_sc_hd__clkbuf_1 _11972_ (.A(_07262_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _11973_ (.A0(\fifo_bank_register.bank[5][57] ),
    .A1(_05390_),
    .S(_07255_),
    .X(_07263_));
 sky130_fd_sc_hd__clkbuf_1 _11974_ (.A(_07263_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _11975_ (.A0(\fifo_bank_register.bank[5][58] ),
    .A1(_05392_),
    .S(_07255_),
    .X(_07264_));
 sky130_fd_sc_hd__clkbuf_1 _11976_ (.A(_07264_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _11977_ (.A0(\fifo_bank_register.bank[5][59] ),
    .A1(_05394_),
    .S(_07255_),
    .X(_07265_));
 sky130_fd_sc_hd__clkbuf_1 _11978_ (.A(_07265_),
    .X(_00724_));
 sky130_fd_sc_hd__buf_4 _11979_ (.A(_07221_),
    .X(_07266_));
 sky130_fd_sc_hd__mux2_1 _11980_ (.A0(\fifo_bank_register.bank[5][60] ),
    .A1(_05396_),
    .S(_07266_),
    .X(_07267_));
 sky130_fd_sc_hd__clkbuf_1 _11981_ (.A(_07267_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _11982_ (.A0(\fifo_bank_register.bank[5][61] ),
    .A1(_05399_),
    .S(_07266_),
    .X(_07268_));
 sky130_fd_sc_hd__clkbuf_1 _11983_ (.A(_07268_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _11984_ (.A0(\fifo_bank_register.bank[5][62] ),
    .A1(_05401_),
    .S(_07266_),
    .X(_07269_));
 sky130_fd_sc_hd__clkbuf_1 _11985_ (.A(_07269_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _11986_ (.A0(\fifo_bank_register.bank[5][63] ),
    .A1(_05403_),
    .S(_07266_),
    .X(_07270_));
 sky130_fd_sc_hd__clkbuf_1 _11987_ (.A(_07270_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _11988_ (.A0(\fifo_bank_register.bank[5][64] ),
    .A1(_05405_),
    .S(_07266_),
    .X(_07271_));
 sky130_fd_sc_hd__clkbuf_1 _11989_ (.A(_07271_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _11990_ (.A0(\fifo_bank_register.bank[5][65] ),
    .A1(_05407_),
    .S(_07266_),
    .X(_07272_));
 sky130_fd_sc_hd__clkbuf_1 _11991_ (.A(_07272_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _11992_ (.A0(\fifo_bank_register.bank[5][66] ),
    .A1(_05409_),
    .S(_07266_),
    .X(_07273_));
 sky130_fd_sc_hd__clkbuf_1 _11993_ (.A(_07273_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _11994_ (.A0(\fifo_bank_register.bank[5][67] ),
    .A1(_05411_),
    .S(_07266_),
    .X(_07274_));
 sky130_fd_sc_hd__clkbuf_1 _11995_ (.A(_07274_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _11996_ (.A0(\fifo_bank_register.bank[5][68] ),
    .A1(_05413_),
    .S(_07266_),
    .X(_07275_));
 sky130_fd_sc_hd__clkbuf_1 _11997_ (.A(_07275_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _11998_ (.A0(\fifo_bank_register.bank[5][69] ),
    .A1(_05415_),
    .S(_07266_),
    .X(_07276_));
 sky130_fd_sc_hd__clkbuf_1 _11999_ (.A(_07276_),
    .X(_00734_));
 sky130_fd_sc_hd__clkbuf_4 _12000_ (.A(_07221_),
    .X(_07277_));
 sky130_fd_sc_hd__mux2_1 _12001_ (.A0(\fifo_bank_register.bank[5][70] ),
    .A1(_05417_),
    .S(_07277_),
    .X(_07278_));
 sky130_fd_sc_hd__clkbuf_1 _12002_ (.A(_07278_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _12003_ (.A0(\fifo_bank_register.bank[5][71] ),
    .A1(_05420_),
    .S(_07277_),
    .X(_07279_));
 sky130_fd_sc_hd__clkbuf_1 _12004_ (.A(_07279_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _12005_ (.A0(\fifo_bank_register.bank[5][72] ),
    .A1(_05422_),
    .S(_07277_),
    .X(_07280_));
 sky130_fd_sc_hd__clkbuf_1 _12006_ (.A(_07280_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _12007_ (.A0(\fifo_bank_register.bank[5][73] ),
    .A1(_05424_),
    .S(_07277_),
    .X(_07281_));
 sky130_fd_sc_hd__clkbuf_1 _12008_ (.A(_07281_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _12009_ (.A0(\fifo_bank_register.bank[5][74] ),
    .A1(_05426_),
    .S(_07277_),
    .X(_07282_));
 sky130_fd_sc_hd__clkbuf_1 _12010_ (.A(_07282_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _12011_ (.A0(\fifo_bank_register.bank[5][75] ),
    .A1(_05428_),
    .S(_07277_),
    .X(_07283_));
 sky130_fd_sc_hd__clkbuf_1 _12012_ (.A(_07283_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _12013_ (.A0(\fifo_bank_register.bank[5][76] ),
    .A1(_05430_),
    .S(_07277_),
    .X(_07284_));
 sky130_fd_sc_hd__clkbuf_1 _12014_ (.A(_07284_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _12015_ (.A0(\fifo_bank_register.bank[5][77] ),
    .A1(_05432_),
    .S(_07277_),
    .X(_07285_));
 sky130_fd_sc_hd__clkbuf_1 _12016_ (.A(_07285_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _12017_ (.A0(\fifo_bank_register.bank[5][78] ),
    .A1(_05434_),
    .S(_07277_),
    .X(_07286_));
 sky130_fd_sc_hd__clkbuf_1 _12018_ (.A(_07286_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _12019_ (.A0(\fifo_bank_register.bank[5][79] ),
    .A1(_05436_),
    .S(_07277_),
    .X(_07287_));
 sky130_fd_sc_hd__clkbuf_1 _12020_ (.A(_07287_),
    .X(_00744_));
 sky130_fd_sc_hd__buf_4 _12021_ (.A(_07221_),
    .X(_07288_));
 sky130_fd_sc_hd__mux2_1 _12022_ (.A0(\fifo_bank_register.bank[5][80] ),
    .A1(_05438_),
    .S(_07288_),
    .X(_07289_));
 sky130_fd_sc_hd__clkbuf_1 _12023_ (.A(_07289_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _12024_ (.A0(\fifo_bank_register.bank[5][81] ),
    .A1(_05441_),
    .S(_07288_),
    .X(_07290_));
 sky130_fd_sc_hd__clkbuf_1 _12025_ (.A(_07290_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _12026_ (.A0(\fifo_bank_register.bank[5][82] ),
    .A1(_05443_),
    .S(_07288_),
    .X(_07291_));
 sky130_fd_sc_hd__clkbuf_1 _12027_ (.A(_07291_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _12028_ (.A0(\fifo_bank_register.bank[5][83] ),
    .A1(_05445_),
    .S(_07288_),
    .X(_07292_));
 sky130_fd_sc_hd__clkbuf_1 _12029_ (.A(_07292_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _12030_ (.A0(\fifo_bank_register.bank[5][84] ),
    .A1(_05447_),
    .S(_07288_),
    .X(_07293_));
 sky130_fd_sc_hd__clkbuf_1 _12031_ (.A(_07293_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _12032_ (.A0(\fifo_bank_register.bank[5][85] ),
    .A1(_05449_),
    .S(_07288_),
    .X(_07294_));
 sky130_fd_sc_hd__clkbuf_1 _12033_ (.A(_07294_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _12034_ (.A0(\fifo_bank_register.bank[5][86] ),
    .A1(_05451_),
    .S(_07288_),
    .X(_07295_));
 sky130_fd_sc_hd__clkbuf_1 _12035_ (.A(_07295_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _12036_ (.A0(\fifo_bank_register.bank[5][87] ),
    .A1(_05453_),
    .S(_07288_),
    .X(_07296_));
 sky130_fd_sc_hd__clkbuf_1 _12037_ (.A(_07296_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _12038_ (.A0(\fifo_bank_register.bank[5][88] ),
    .A1(_05455_),
    .S(_07288_),
    .X(_07297_));
 sky130_fd_sc_hd__clkbuf_1 _12039_ (.A(_07297_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _12040_ (.A0(\fifo_bank_register.bank[5][89] ),
    .A1(_05457_),
    .S(_07288_),
    .X(_07298_));
 sky130_fd_sc_hd__clkbuf_1 _12041_ (.A(_07298_),
    .X(_00754_));
 sky130_fd_sc_hd__buf_4 _12042_ (.A(_07221_),
    .X(_07299_));
 sky130_fd_sc_hd__mux2_1 _12043_ (.A0(\fifo_bank_register.bank[5][90] ),
    .A1(_05459_),
    .S(_07299_),
    .X(_07300_));
 sky130_fd_sc_hd__clkbuf_1 _12044_ (.A(_07300_),
    .X(_00755_));
 sky130_fd_sc_hd__mux2_1 _12045_ (.A0(\fifo_bank_register.bank[5][91] ),
    .A1(_05462_),
    .S(_07299_),
    .X(_07301_));
 sky130_fd_sc_hd__clkbuf_1 _12046_ (.A(_07301_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _12047_ (.A0(\fifo_bank_register.bank[5][92] ),
    .A1(_05464_),
    .S(_07299_),
    .X(_07302_));
 sky130_fd_sc_hd__clkbuf_1 _12048_ (.A(_07302_),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _12049_ (.A0(\fifo_bank_register.bank[5][93] ),
    .A1(_05466_),
    .S(_07299_),
    .X(_07303_));
 sky130_fd_sc_hd__clkbuf_1 _12050_ (.A(_07303_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _12051_ (.A0(\fifo_bank_register.bank[5][94] ),
    .A1(_05468_),
    .S(_07299_),
    .X(_07304_));
 sky130_fd_sc_hd__clkbuf_1 _12052_ (.A(_07304_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _12053_ (.A0(\fifo_bank_register.bank[5][95] ),
    .A1(_05470_),
    .S(_07299_),
    .X(_07305_));
 sky130_fd_sc_hd__clkbuf_1 _12054_ (.A(_07305_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _12055_ (.A0(\fifo_bank_register.bank[5][96] ),
    .A1(_05472_),
    .S(_07299_),
    .X(_07306_));
 sky130_fd_sc_hd__clkbuf_1 _12056_ (.A(_07306_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _12057_ (.A0(\fifo_bank_register.bank[5][97] ),
    .A1(_05474_),
    .S(_07299_),
    .X(_07307_));
 sky130_fd_sc_hd__clkbuf_1 _12058_ (.A(_07307_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _12059_ (.A0(\fifo_bank_register.bank[5][98] ),
    .A1(_05476_),
    .S(_07299_),
    .X(_07308_));
 sky130_fd_sc_hd__clkbuf_1 _12060_ (.A(_07308_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _12061_ (.A0(\fifo_bank_register.bank[5][99] ),
    .A1(_05478_),
    .S(_07299_),
    .X(_07309_));
 sky130_fd_sc_hd__clkbuf_1 _12062_ (.A(_07309_),
    .X(_00764_));
 sky130_fd_sc_hd__buf_4 _12063_ (.A(_07221_),
    .X(_07310_));
 sky130_fd_sc_hd__mux2_1 _12064_ (.A0(\fifo_bank_register.bank[5][100] ),
    .A1(_05480_),
    .S(_07310_),
    .X(_07311_));
 sky130_fd_sc_hd__clkbuf_1 _12065_ (.A(_07311_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _12066_ (.A0(\fifo_bank_register.bank[5][101] ),
    .A1(_05483_),
    .S(_07310_),
    .X(_07312_));
 sky130_fd_sc_hd__clkbuf_1 _12067_ (.A(_07312_),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _12068_ (.A0(\fifo_bank_register.bank[5][102] ),
    .A1(_05485_),
    .S(_07310_),
    .X(_07313_));
 sky130_fd_sc_hd__clkbuf_1 _12069_ (.A(_07313_),
    .X(_00767_));
 sky130_fd_sc_hd__mux2_1 _12070_ (.A0(\fifo_bank_register.bank[5][103] ),
    .A1(_05487_),
    .S(_07310_),
    .X(_07314_));
 sky130_fd_sc_hd__clkbuf_1 _12071_ (.A(_07314_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _12072_ (.A0(\fifo_bank_register.bank[5][104] ),
    .A1(_05489_),
    .S(_07310_),
    .X(_07315_));
 sky130_fd_sc_hd__clkbuf_1 _12073_ (.A(_07315_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _12074_ (.A0(\fifo_bank_register.bank[5][105] ),
    .A1(_05491_),
    .S(_07310_),
    .X(_07316_));
 sky130_fd_sc_hd__clkbuf_1 _12075_ (.A(_07316_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _12076_ (.A0(\fifo_bank_register.bank[5][106] ),
    .A1(_05493_),
    .S(_07310_),
    .X(_07317_));
 sky130_fd_sc_hd__clkbuf_1 _12077_ (.A(_07317_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _12078_ (.A0(\fifo_bank_register.bank[5][107] ),
    .A1(_05495_),
    .S(_07310_),
    .X(_07318_));
 sky130_fd_sc_hd__clkbuf_1 _12079_ (.A(_07318_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _12080_ (.A0(\fifo_bank_register.bank[5][108] ),
    .A1(_05497_),
    .S(_07310_),
    .X(_07319_));
 sky130_fd_sc_hd__clkbuf_1 _12081_ (.A(_07319_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _12082_ (.A0(\fifo_bank_register.bank[5][109] ),
    .A1(_05499_),
    .S(_07310_),
    .X(_07320_));
 sky130_fd_sc_hd__clkbuf_1 _12083_ (.A(_07320_),
    .X(_00774_));
 sky130_fd_sc_hd__buf_4 _12084_ (.A(_07221_),
    .X(_07321_));
 sky130_fd_sc_hd__mux2_1 _12085_ (.A0(\fifo_bank_register.bank[5][110] ),
    .A1(_05501_),
    .S(_07321_),
    .X(_07322_));
 sky130_fd_sc_hd__clkbuf_1 _12086_ (.A(_07322_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _12087_ (.A0(\fifo_bank_register.bank[5][111] ),
    .A1(_05504_),
    .S(_07321_),
    .X(_07323_));
 sky130_fd_sc_hd__clkbuf_1 _12088_ (.A(_07323_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _12089_ (.A0(\fifo_bank_register.bank[5][112] ),
    .A1(_05506_),
    .S(_07321_),
    .X(_07324_));
 sky130_fd_sc_hd__clkbuf_1 _12090_ (.A(_07324_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _12091_ (.A0(\fifo_bank_register.bank[5][113] ),
    .A1(_05508_),
    .S(_07321_),
    .X(_07325_));
 sky130_fd_sc_hd__clkbuf_1 _12092_ (.A(_07325_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _12093_ (.A0(\fifo_bank_register.bank[5][114] ),
    .A1(_05510_),
    .S(_07321_),
    .X(_07326_));
 sky130_fd_sc_hd__clkbuf_1 _12094_ (.A(_07326_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _12095_ (.A0(\fifo_bank_register.bank[5][115] ),
    .A1(_05512_),
    .S(_07321_),
    .X(_07327_));
 sky130_fd_sc_hd__clkbuf_1 _12096_ (.A(_07327_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _12097_ (.A0(\fifo_bank_register.bank[5][116] ),
    .A1(_05514_),
    .S(_07321_),
    .X(_07328_));
 sky130_fd_sc_hd__clkbuf_1 _12098_ (.A(_07328_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _12099_ (.A0(\fifo_bank_register.bank[5][117] ),
    .A1(_05516_),
    .S(_07321_),
    .X(_07329_));
 sky130_fd_sc_hd__clkbuf_1 _12100_ (.A(_07329_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _12101_ (.A0(\fifo_bank_register.bank[5][118] ),
    .A1(_05518_),
    .S(_07321_),
    .X(_07330_));
 sky130_fd_sc_hd__clkbuf_1 _12102_ (.A(_07330_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _12103_ (.A0(\fifo_bank_register.bank[5][119] ),
    .A1(_05520_),
    .S(_07321_),
    .X(_07331_));
 sky130_fd_sc_hd__clkbuf_1 _12104_ (.A(_07331_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _12105_ (.A0(\fifo_bank_register.bank[5][120] ),
    .A1(_05522_),
    .S(_07198_),
    .X(_07332_));
 sky130_fd_sc_hd__clkbuf_1 _12106_ (.A(_07332_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _12107_ (.A0(\fifo_bank_register.bank[5][121] ),
    .A1(_05524_),
    .S(_07198_),
    .X(_07333_));
 sky130_fd_sc_hd__clkbuf_1 _12108_ (.A(_07333_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _12109_ (.A0(\fifo_bank_register.bank[5][122] ),
    .A1(_05526_),
    .S(_07198_),
    .X(_07334_));
 sky130_fd_sc_hd__clkbuf_1 _12110_ (.A(_07334_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _12111_ (.A0(\fifo_bank_register.bank[5][123] ),
    .A1(_05528_),
    .S(_07198_),
    .X(_07335_));
 sky130_fd_sc_hd__clkbuf_1 _12112_ (.A(_07335_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _12113_ (.A0(\fifo_bank_register.bank[5][124] ),
    .A1(_05530_),
    .S(_07198_),
    .X(_07336_));
 sky130_fd_sc_hd__clkbuf_1 _12114_ (.A(_07336_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _12115_ (.A0(\fifo_bank_register.bank[5][125] ),
    .A1(_05532_),
    .S(_07198_),
    .X(_07337_));
 sky130_fd_sc_hd__clkbuf_1 _12116_ (.A(_07337_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _12117_ (.A0(\fifo_bank_register.bank[5][126] ),
    .A1(_05534_),
    .S(_07198_),
    .X(_07338_));
 sky130_fd_sc_hd__clkbuf_1 _12118_ (.A(_07338_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _12119_ (.A0(\fifo_bank_register.bank[5][127] ),
    .A1(_05536_),
    .S(_07198_),
    .X(_07339_));
 sky130_fd_sc_hd__clkbuf_1 _12120_ (.A(_07339_),
    .X(_00792_));
 sky130_fd_sc_hd__or2b_1 _12121_ (.A(_06766_),
    .B_N(_06910_),
    .X(_07340_));
 sky130_fd_sc_hd__buf_4 _12122_ (.A(_07340_),
    .X(_07341_));
 sky130_fd_sc_hd__clkbuf_4 _12123_ (.A(_07341_),
    .X(_07342_));
 sky130_fd_sc_hd__mux2_1 _12124_ (.A0(_05248_),
    .A1(\fifo_bank_register.bank[4][0] ),
    .S(_07342_),
    .X(_07343_));
 sky130_fd_sc_hd__clkbuf_1 _12125_ (.A(_07343_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _12126_ (.A0(_05272_),
    .A1(\fifo_bank_register.bank[4][1] ),
    .S(_07342_),
    .X(_07344_));
 sky130_fd_sc_hd__clkbuf_1 _12127_ (.A(_07344_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _12128_ (.A0(_05274_),
    .A1(\fifo_bank_register.bank[4][2] ),
    .S(_07342_),
    .X(_07345_));
 sky130_fd_sc_hd__clkbuf_1 _12129_ (.A(_07345_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _12130_ (.A0(_05276_),
    .A1(\fifo_bank_register.bank[4][3] ),
    .S(_07342_),
    .X(_07346_));
 sky130_fd_sc_hd__clkbuf_1 _12131_ (.A(_07346_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _12132_ (.A0(_05278_),
    .A1(\fifo_bank_register.bank[4][4] ),
    .S(_07342_),
    .X(_07347_));
 sky130_fd_sc_hd__clkbuf_1 _12133_ (.A(_07347_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _12134_ (.A0(_05280_),
    .A1(\fifo_bank_register.bank[4][5] ),
    .S(_07342_),
    .X(_07348_));
 sky130_fd_sc_hd__clkbuf_1 _12135_ (.A(_07348_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _12136_ (.A0(_05282_),
    .A1(\fifo_bank_register.bank[4][6] ),
    .S(_07342_),
    .X(_07349_));
 sky130_fd_sc_hd__clkbuf_1 _12137_ (.A(_07349_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _12138_ (.A0(_05284_),
    .A1(\fifo_bank_register.bank[4][7] ),
    .S(_07342_),
    .X(_07350_));
 sky130_fd_sc_hd__clkbuf_1 _12139_ (.A(_07350_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _12140_ (.A0(_05286_),
    .A1(\fifo_bank_register.bank[4][8] ),
    .S(_07342_),
    .X(_07351_));
 sky130_fd_sc_hd__clkbuf_1 _12141_ (.A(_07351_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _12142_ (.A0(_05288_),
    .A1(\fifo_bank_register.bank[4][9] ),
    .S(_07342_),
    .X(_07352_));
 sky130_fd_sc_hd__clkbuf_1 _12143_ (.A(_07352_),
    .X(_00802_));
 sky130_fd_sc_hd__buf_4 _12144_ (.A(_07341_),
    .X(_07353_));
 sky130_fd_sc_hd__mux2_1 _12145_ (.A0(_05290_),
    .A1(\fifo_bank_register.bank[4][10] ),
    .S(_07353_),
    .X(_07354_));
 sky130_fd_sc_hd__clkbuf_1 _12146_ (.A(_07354_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _12147_ (.A0(_05293_),
    .A1(\fifo_bank_register.bank[4][11] ),
    .S(_07353_),
    .X(_07355_));
 sky130_fd_sc_hd__clkbuf_1 _12148_ (.A(_07355_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _12149_ (.A0(_05295_),
    .A1(\fifo_bank_register.bank[4][12] ),
    .S(_07353_),
    .X(_07356_));
 sky130_fd_sc_hd__clkbuf_1 _12150_ (.A(_07356_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _12151_ (.A0(_05297_),
    .A1(\fifo_bank_register.bank[4][13] ),
    .S(_07353_),
    .X(_07357_));
 sky130_fd_sc_hd__clkbuf_1 _12152_ (.A(_07357_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _12153_ (.A0(_05299_),
    .A1(\fifo_bank_register.bank[4][14] ),
    .S(_07353_),
    .X(_07358_));
 sky130_fd_sc_hd__clkbuf_1 _12154_ (.A(_07358_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _12155_ (.A0(_05301_),
    .A1(\fifo_bank_register.bank[4][15] ),
    .S(_07353_),
    .X(_07359_));
 sky130_fd_sc_hd__clkbuf_1 _12156_ (.A(_07359_),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _12157_ (.A0(_05303_),
    .A1(\fifo_bank_register.bank[4][16] ),
    .S(_07353_),
    .X(_07360_));
 sky130_fd_sc_hd__clkbuf_1 _12158_ (.A(_07360_),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _12159_ (.A0(_05305_),
    .A1(\fifo_bank_register.bank[4][17] ),
    .S(_07353_),
    .X(_07361_));
 sky130_fd_sc_hd__clkbuf_1 _12160_ (.A(_07361_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _12161_ (.A0(_05307_),
    .A1(\fifo_bank_register.bank[4][18] ),
    .S(_07353_),
    .X(_07362_));
 sky130_fd_sc_hd__clkbuf_1 _12162_ (.A(_07362_),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _12163_ (.A0(_05309_),
    .A1(\fifo_bank_register.bank[4][19] ),
    .S(_07353_),
    .X(_07363_));
 sky130_fd_sc_hd__clkbuf_1 _12164_ (.A(_07363_),
    .X(_00812_));
 sky130_fd_sc_hd__buf_6 _12165_ (.A(_07340_),
    .X(_07364_));
 sky130_fd_sc_hd__buf_4 _12166_ (.A(_07364_),
    .X(_07365_));
 sky130_fd_sc_hd__mux2_1 _12167_ (.A0(_05311_),
    .A1(\fifo_bank_register.bank[4][20] ),
    .S(_07365_),
    .X(_07366_));
 sky130_fd_sc_hd__clkbuf_1 _12168_ (.A(_07366_),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _12169_ (.A0(_05315_),
    .A1(\fifo_bank_register.bank[4][21] ),
    .S(_07365_),
    .X(_07367_));
 sky130_fd_sc_hd__clkbuf_1 _12170_ (.A(_07367_),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _12171_ (.A0(_05317_),
    .A1(\fifo_bank_register.bank[4][22] ),
    .S(_07365_),
    .X(_07368_));
 sky130_fd_sc_hd__clkbuf_1 _12172_ (.A(_07368_),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(_05319_),
    .A1(\fifo_bank_register.bank[4][23] ),
    .S(_07365_),
    .X(_07369_));
 sky130_fd_sc_hd__clkbuf_1 _12174_ (.A(_07369_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(_05321_),
    .A1(\fifo_bank_register.bank[4][24] ),
    .S(_07365_),
    .X(_07370_));
 sky130_fd_sc_hd__clkbuf_1 _12176_ (.A(_07370_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _12177_ (.A0(_05323_),
    .A1(\fifo_bank_register.bank[4][25] ),
    .S(_07365_),
    .X(_07371_));
 sky130_fd_sc_hd__clkbuf_1 _12178_ (.A(_07371_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _12179_ (.A0(_05325_),
    .A1(\fifo_bank_register.bank[4][26] ),
    .S(_07365_),
    .X(_07372_));
 sky130_fd_sc_hd__clkbuf_1 _12180_ (.A(_07372_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _12181_ (.A0(_05327_),
    .A1(\fifo_bank_register.bank[4][27] ),
    .S(_07365_),
    .X(_07373_));
 sky130_fd_sc_hd__clkbuf_1 _12182_ (.A(_07373_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _12183_ (.A0(_05329_),
    .A1(\fifo_bank_register.bank[4][28] ),
    .S(_07365_),
    .X(_07374_));
 sky130_fd_sc_hd__clkbuf_1 _12184_ (.A(_07374_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _12185_ (.A0(_05331_),
    .A1(\fifo_bank_register.bank[4][29] ),
    .S(_07365_),
    .X(_07375_));
 sky130_fd_sc_hd__clkbuf_1 _12186_ (.A(_07375_),
    .X(_00822_));
 sky130_fd_sc_hd__buf_4 _12187_ (.A(_07364_),
    .X(_07376_));
 sky130_fd_sc_hd__mux2_1 _12188_ (.A0(_05333_),
    .A1(\fifo_bank_register.bank[4][30] ),
    .S(_07376_),
    .X(_07377_));
 sky130_fd_sc_hd__clkbuf_1 _12189_ (.A(_07377_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _12190_ (.A0(_05336_),
    .A1(\fifo_bank_register.bank[4][31] ),
    .S(_07376_),
    .X(_07378_));
 sky130_fd_sc_hd__clkbuf_1 _12191_ (.A(_07378_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _12192_ (.A0(_05338_),
    .A1(\fifo_bank_register.bank[4][32] ),
    .S(_07376_),
    .X(_07379_));
 sky130_fd_sc_hd__clkbuf_1 _12193_ (.A(_07379_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _12194_ (.A0(_05340_),
    .A1(\fifo_bank_register.bank[4][33] ),
    .S(_07376_),
    .X(_07380_));
 sky130_fd_sc_hd__clkbuf_1 _12195_ (.A(_07380_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _12196_ (.A0(_05342_),
    .A1(\fifo_bank_register.bank[4][34] ),
    .S(_07376_),
    .X(_07381_));
 sky130_fd_sc_hd__clkbuf_1 _12197_ (.A(_07381_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _12198_ (.A0(_05344_),
    .A1(\fifo_bank_register.bank[4][35] ),
    .S(_07376_),
    .X(_07382_));
 sky130_fd_sc_hd__clkbuf_1 _12199_ (.A(_07382_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _12200_ (.A0(_05346_),
    .A1(\fifo_bank_register.bank[4][36] ),
    .S(_07376_),
    .X(_07383_));
 sky130_fd_sc_hd__clkbuf_1 _12201_ (.A(_07383_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _12202_ (.A0(_05348_),
    .A1(\fifo_bank_register.bank[4][37] ),
    .S(_07376_),
    .X(_07384_));
 sky130_fd_sc_hd__clkbuf_1 _12203_ (.A(_07384_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _12204_ (.A0(_05350_),
    .A1(\fifo_bank_register.bank[4][38] ),
    .S(_07376_),
    .X(_07385_));
 sky130_fd_sc_hd__clkbuf_1 _12205_ (.A(_07385_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _12206_ (.A0(_05352_),
    .A1(\fifo_bank_register.bank[4][39] ),
    .S(_07376_),
    .X(_07386_));
 sky130_fd_sc_hd__clkbuf_1 _12207_ (.A(_07386_),
    .X(_00832_));
 sky130_fd_sc_hd__buf_4 _12208_ (.A(_07364_),
    .X(_07387_));
 sky130_fd_sc_hd__mux2_1 _12209_ (.A0(_05354_),
    .A1(\fifo_bank_register.bank[4][40] ),
    .S(_07387_),
    .X(_07388_));
 sky130_fd_sc_hd__clkbuf_1 _12210_ (.A(_07388_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _12211_ (.A0(_05357_),
    .A1(\fifo_bank_register.bank[4][41] ),
    .S(_07387_),
    .X(_07389_));
 sky130_fd_sc_hd__clkbuf_1 _12212_ (.A(_07389_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _12213_ (.A0(_05359_),
    .A1(\fifo_bank_register.bank[4][42] ),
    .S(_07387_),
    .X(_07390_));
 sky130_fd_sc_hd__clkbuf_1 _12214_ (.A(_07390_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _12215_ (.A0(_05361_),
    .A1(\fifo_bank_register.bank[4][43] ),
    .S(_07387_),
    .X(_07391_));
 sky130_fd_sc_hd__clkbuf_1 _12216_ (.A(_07391_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _12217_ (.A0(_05363_),
    .A1(\fifo_bank_register.bank[4][44] ),
    .S(_07387_),
    .X(_07392_));
 sky130_fd_sc_hd__clkbuf_1 _12218_ (.A(_07392_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _12219_ (.A0(_05365_),
    .A1(\fifo_bank_register.bank[4][45] ),
    .S(_07387_),
    .X(_07393_));
 sky130_fd_sc_hd__clkbuf_1 _12220_ (.A(_07393_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _12221_ (.A0(_05367_),
    .A1(\fifo_bank_register.bank[4][46] ),
    .S(_07387_),
    .X(_07394_));
 sky130_fd_sc_hd__clkbuf_1 _12222_ (.A(_07394_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _12223_ (.A0(_05369_),
    .A1(\fifo_bank_register.bank[4][47] ),
    .S(_07387_),
    .X(_07395_));
 sky130_fd_sc_hd__clkbuf_1 _12224_ (.A(_07395_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _12225_ (.A0(_05371_),
    .A1(\fifo_bank_register.bank[4][48] ),
    .S(_07387_),
    .X(_07396_));
 sky130_fd_sc_hd__clkbuf_1 _12226_ (.A(_07396_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _12227_ (.A0(_05373_),
    .A1(\fifo_bank_register.bank[4][49] ),
    .S(_07387_),
    .X(_07397_));
 sky130_fd_sc_hd__clkbuf_1 _12228_ (.A(_07397_),
    .X(_00842_));
 sky130_fd_sc_hd__buf_4 _12229_ (.A(_07364_),
    .X(_07398_));
 sky130_fd_sc_hd__mux2_1 _12230_ (.A0(_05375_),
    .A1(\fifo_bank_register.bank[4][50] ),
    .S(_07398_),
    .X(_07399_));
 sky130_fd_sc_hd__clkbuf_1 _12231_ (.A(_07399_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _12232_ (.A0(_05378_),
    .A1(\fifo_bank_register.bank[4][51] ),
    .S(_07398_),
    .X(_07400_));
 sky130_fd_sc_hd__clkbuf_1 _12233_ (.A(_07400_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _12234_ (.A0(_05380_),
    .A1(\fifo_bank_register.bank[4][52] ),
    .S(_07398_),
    .X(_07401_));
 sky130_fd_sc_hd__clkbuf_1 _12235_ (.A(_07401_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _12236_ (.A0(_05382_),
    .A1(\fifo_bank_register.bank[4][53] ),
    .S(_07398_),
    .X(_07402_));
 sky130_fd_sc_hd__clkbuf_1 _12237_ (.A(_07402_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _12238_ (.A0(_05384_),
    .A1(\fifo_bank_register.bank[4][54] ),
    .S(_07398_),
    .X(_07403_));
 sky130_fd_sc_hd__clkbuf_1 _12239_ (.A(_07403_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(_05386_),
    .A1(\fifo_bank_register.bank[4][55] ),
    .S(_07398_),
    .X(_07404_));
 sky130_fd_sc_hd__clkbuf_1 _12241_ (.A(_07404_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _12242_ (.A0(_05388_),
    .A1(\fifo_bank_register.bank[4][56] ),
    .S(_07398_),
    .X(_07405_));
 sky130_fd_sc_hd__clkbuf_1 _12243_ (.A(_07405_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _12244_ (.A0(_05390_),
    .A1(\fifo_bank_register.bank[4][57] ),
    .S(_07398_),
    .X(_07406_));
 sky130_fd_sc_hd__clkbuf_1 _12245_ (.A(_07406_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _12246_ (.A0(_05392_),
    .A1(\fifo_bank_register.bank[4][58] ),
    .S(_07398_),
    .X(_07407_));
 sky130_fd_sc_hd__clkbuf_1 _12247_ (.A(_07407_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _12248_ (.A0(_05394_),
    .A1(\fifo_bank_register.bank[4][59] ),
    .S(_07398_),
    .X(_07408_));
 sky130_fd_sc_hd__clkbuf_1 _12249_ (.A(_07408_),
    .X(_00852_));
 sky130_fd_sc_hd__buf_4 _12250_ (.A(_07364_),
    .X(_07409_));
 sky130_fd_sc_hd__mux2_1 _12251_ (.A0(_05396_),
    .A1(\fifo_bank_register.bank[4][60] ),
    .S(_07409_),
    .X(_07410_));
 sky130_fd_sc_hd__clkbuf_1 _12252_ (.A(_07410_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _12253_ (.A0(_05399_),
    .A1(\fifo_bank_register.bank[4][61] ),
    .S(_07409_),
    .X(_07411_));
 sky130_fd_sc_hd__clkbuf_1 _12254_ (.A(_07411_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _12255_ (.A0(_05401_),
    .A1(\fifo_bank_register.bank[4][62] ),
    .S(_07409_),
    .X(_07412_));
 sky130_fd_sc_hd__clkbuf_1 _12256_ (.A(_07412_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _12257_ (.A0(_05403_),
    .A1(\fifo_bank_register.bank[4][63] ),
    .S(_07409_),
    .X(_07413_));
 sky130_fd_sc_hd__clkbuf_1 _12258_ (.A(_07413_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _12259_ (.A0(_05405_),
    .A1(\fifo_bank_register.bank[4][64] ),
    .S(_07409_),
    .X(_07414_));
 sky130_fd_sc_hd__clkbuf_1 _12260_ (.A(_07414_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _12261_ (.A0(_05407_),
    .A1(\fifo_bank_register.bank[4][65] ),
    .S(_07409_),
    .X(_07415_));
 sky130_fd_sc_hd__clkbuf_1 _12262_ (.A(_07415_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _12263_ (.A0(_05409_),
    .A1(\fifo_bank_register.bank[4][66] ),
    .S(_07409_),
    .X(_07416_));
 sky130_fd_sc_hd__clkbuf_1 _12264_ (.A(_07416_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _12265_ (.A0(_05411_),
    .A1(\fifo_bank_register.bank[4][67] ),
    .S(_07409_),
    .X(_07417_));
 sky130_fd_sc_hd__clkbuf_1 _12266_ (.A(_07417_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _12267_ (.A0(_05413_),
    .A1(\fifo_bank_register.bank[4][68] ),
    .S(_07409_),
    .X(_07418_));
 sky130_fd_sc_hd__clkbuf_1 _12268_ (.A(_07418_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _12269_ (.A0(_05415_),
    .A1(\fifo_bank_register.bank[4][69] ),
    .S(_07409_),
    .X(_07419_));
 sky130_fd_sc_hd__clkbuf_1 _12270_ (.A(_07419_),
    .X(_00862_));
 sky130_fd_sc_hd__buf_4 _12271_ (.A(_07364_),
    .X(_07420_));
 sky130_fd_sc_hd__mux2_1 _12272_ (.A0(_05417_),
    .A1(\fifo_bank_register.bank[4][70] ),
    .S(_07420_),
    .X(_07421_));
 sky130_fd_sc_hd__clkbuf_1 _12273_ (.A(_07421_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _12274_ (.A0(_05420_),
    .A1(\fifo_bank_register.bank[4][71] ),
    .S(_07420_),
    .X(_07422_));
 sky130_fd_sc_hd__clkbuf_1 _12275_ (.A(_07422_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _12276_ (.A0(_05422_),
    .A1(\fifo_bank_register.bank[4][72] ),
    .S(_07420_),
    .X(_07423_));
 sky130_fd_sc_hd__clkbuf_1 _12277_ (.A(_07423_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _12278_ (.A0(_05424_),
    .A1(\fifo_bank_register.bank[4][73] ),
    .S(_07420_),
    .X(_07424_));
 sky130_fd_sc_hd__clkbuf_1 _12279_ (.A(_07424_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _12280_ (.A0(_05426_),
    .A1(\fifo_bank_register.bank[4][74] ),
    .S(_07420_),
    .X(_07425_));
 sky130_fd_sc_hd__clkbuf_1 _12281_ (.A(_07425_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _12282_ (.A0(_05428_),
    .A1(\fifo_bank_register.bank[4][75] ),
    .S(_07420_),
    .X(_07426_));
 sky130_fd_sc_hd__clkbuf_1 _12283_ (.A(_07426_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _12284_ (.A0(_05430_),
    .A1(\fifo_bank_register.bank[4][76] ),
    .S(_07420_),
    .X(_07427_));
 sky130_fd_sc_hd__clkbuf_1 _12285_ (.A(_07427_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _12286_ (.A0(_05432_),
    .A1(\fifo_bank_register.bank[4][77] ),
    .S(_07420_),
    .X(_07428_));
 sky130_fd_sc_hd__clkbuf_1 _12287_ (.A(_07428_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _12288_ (.A0(_05434_),
    .A1(\fifo_bank_register.bank[4][78] ),
    .S(_07420_),
    .X(_07429_));
 sky130_fd_sc_hd__clkbuf_1 _12289_ (.A(_07429_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _12290_ (.A0(_05436_),
    .A1(\fifo_bank_register.bank[4][79] ),
    .S(_07420_),
    .X(_07430_));
 sky130_fd_sc_hd__clkbuf_1 _12291_ (.A(_07430_),
    .X(_00872_));
 sky130_fd_sc_hd__buf_4 _12292_ (.A(_07364_),
    .X(_07431_));
 sky130_fd_sc_hd__mux2_1 _12293_ (.A0(_05438_),
    .A1(\fifo_bank_register.bank[4][80] ),
    .S(_07431_),
    .X(_07432_));
 sky130_fd_sc_hd__clkbuf_1 _12294_ (.A(_07432_),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _12295_ (.A0(_05441_),
    .A1(\fifo_bank_register.bank[4][81] ),
    .S(_07431_),
    .X(_07433_));
 sky130_fd_sc_hd__clkbuf_1 _12296_ (.A(_07433_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _12297_ (.A0(_05443_),
    .A1(\fifo_bank_register.bank[4][82] ),
    .S(_07431_),
    .X(_07434_));
 sky130_fd_sc_hd__clkbuf_1 _12298_ (.A(_07434_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _12299_ (.A0(_05445_),
    .A1(\fifo_bank_register.bank[4][83] ),
    .S(_07431_),
    .X(_07435_));
 sky130_fd_sc_hd__clkbuf_1 _12300_ (.A(_07435_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _12301_ (.A0(_05447_),
    .A1(\fifo_bank_register.bank[4][84] ),
    .S(_07431_),
    .X(_07436_));
 sky130_fd_sc_hd__clkbuf_1 _12302_ (.A(_07436_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _12303_ (.A0(_05449_),
    .A1(\fifo_bank_register.bank[4][85] ),
    .S(_07431_),
    .X(_07437_));
 sky130_fd_sc_hd__clkbuf_1 _12304_ (.A(_07437_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _12305_ (.A0(_05451_),
    .A1(\fifo_bank_register.bank[4][86] ),
    .S(_07431_),
    .X(_07438_));
 sky130_fd_sc_hd__clkbuf_1 _12306_ (.A(_07438_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _12307_ (.A0(_05453_),
    .A1(\fifo_bank_register.bank[4][87] ),
    .S(_07431_),
    .X(_07439_));
 sky130_fd_sc_hd__clkbuf_1 _12308_ (.A(_07439_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(_05455_),
    .A1(\fifo_bank_register.bank[4][88] ),
    .S(_07431_),
    .X(_07440_));
 sky130_fd_sc_hd__clkbuf_1 _12310_ (.A(_07440_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _12311_ (.A0(_05457_),
    .A1(\fifo_bank_register.bank[4][89] ),
    .S(_07431_),
    .X(_07441_));
 sky130_fd_sc_hd__clkbuf_1 _12312_ (.A(_07441_),
    .X(_00882_));
 sky130_fd_sc_hd__buf_4 _12313_ (.A(_07364_),
    .X(_07442_));
 sky130_fd_sc_hd__mux2_1 _12314_ (.A0(_05459_),
    .A1(\fifo_bank_register.bank[4][90] ),
    .S(_07442_),
    .X(_07443_));
 sky130_fd_sc_hd__clkbuf_1 _12315_ (.A(_07443_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _12316_ (.A0(_05462_),
    .A1(\fifo_bank_register.bank[4][91] ),
    .S(_07442_),
    .X(_07444_));
 sky130_fd_sc_hd__clkbuf_1 _12317_ (.A(_07444_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _12318_ (.A0(_05464_),
    .A1(\fifo_bank_register.bank[4][92] ),
    .S(_07442_),
    .X(_07445_));
 sky130_fd_sc_hd__clkbuf_1 _12319_ (.A(_07445_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _12320_ (.A0(_05466_),
    .A1(\fifo_bank_register.bank[4][93] ),
    .S(_07442_),
    .X(_07446_));
 sky130_fd_sc_hd__clkbuf_1 _12321_ (.A(_07446_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _12322_ (.A0(_05468_),
    .A1(\fifo_bank_register.bank[4][94] ),
    .S(_07442_),
    .X(_07447_));
 sky130_fd_sc_hd__clkbuf_1 _12323_ (.A(_07447_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _12324_ (.A0(_05470_),
    .A1(\fifo_bank_register.bank[4][95] ),
    .S(_07442_),
    .X(_07448_));
 sky130_fd_sc_hd__clkbuf_1 _12325_ (.A(_07448_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _12326_ (.A0(_05472_),
    .A1(\fifo_bank_register.bank[4][96] ),
    .S(_07442_),
    .X(_07449_));
 sky130_fd_sc_hd__clkbuf_1 _12327_ (.A(_07449_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _12328_ (.A0(_05474_),
    .A1(\fifo_bank_register.bank[4][97] ),
    .S(_07442_),
    .X(_07450_));
 sky130_fd_sc_hd__clkbuf_1 _12329_ (.A(_07450_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _12330_ (.A0(_05476_),
    .A1(\fifo_bank_register.bank[4][98] ),
    .S(_07442_),
    .X(_07451_));
 sky130_fd_sc_hd__clkbuf_1 _12331_ (.A(_07451_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _12332_ (.A0(_05478_),
    .A1(\fifo_bank_register.bank[4][99] ),
    .S(_07442_),
    .X(_07452_));
 sky130_fd_sc_hd__clkbuf_1 _12333_ (.A(_07452_),
    .X(_00892_));
 sky130_fd_sc_hd__buf_4 _12334_ (.A(_07364_),
    .X(_07453_));
 sky130_fd_sc_hd__mux2_1 _12335_ (.A0(_05480_),
    .A1(\fifo_bank_register.bank[4][100] ),
    .S(_07453_),
    .X(_07454_));
 sky130_fd_sc_hd__clkbuf_1 _12336_ (.A(_07454_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _12337_ (.A0(_05483_),
    .A1(\fifo_bank_register.bank[4][101] ),
    .S(_07453_),
    .X(_07455_));
 sky130_fd_sc_hd__clkbuf_1 _12338_ (.A(_07455_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _12339_ (.A0(_05485_),
    .A1(\fifo_bank_register.bank[4][102] ),
    .S(_07453_),
    .X(_07456_));
 sky130_fd_sc_hd__clkbuf_1 _12340_ (.A(_07456_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _12341_ (.A0(_05487_),
    .A1(\fifo_bank_register.bank[4][103] ),
    .S(_07453_),
    .X(_07457_));
 sky130_fd_sc_hd__clkbuf_1 _12342_ (.A(_07457_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _12343_ (.A0(_05489_),
    .A1(\fifo_bank_register.bank[4][104] ),
    .S(_07453_),
    .X(_07458_));
 sky130_fd_sc_hd__clkbuf_1 _12344_ (.A(_07458_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _12345_ (.A0(_05491_),
    .A1(\fifo_bank_register.bank[4][105] ),
    .S(_07453_),
    .X(_07459_));
 sky130_fd_sc_hd__clkbuf_1 _12346_ (.A(_07459_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _12347_ (.A0(_05493_),
    .A1(\fifo_bank_register.bank[4][106] ),
    .S(_07453_),
    .X(_07460_));
 sky130_fd_sc_hd__clkbuf_1 _12348_ (.A(_07460_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _12349_ (.A0(_05495_),
    .A1(\fifo_bank_register.bank[4][107] ),
    .S(_07453_),
    .X(_07461_));
 sky130_fd_sc_hd__clkbuf_1 _12350_ (.A(_07461_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _12351_ (.A0(_05497_),
    .A1(\fifo_bank_register.bank[4][108] ),
    .S(_07453_),
    .X(_07462_));
 sky130_fd_sc_hd__clkbuf_1 _12352_ (.A(_07462_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _12353_ (.A0(_05499_),
    .A1(\fifo_bank_register.bank[4][109] ),
    .S(_07453_),
    .X(_07463_));
 sky130_fd_sc_hd__clkbuf_1 _12354_ (.A(_07463_),
    .X(_00902_));
 sky130_fd_sc_hd__buf_4 _12355_ (.A(_07364_),
    .X(_07464_));
 sky130_fd_sc_hd__mux2_1 _12356_ (.A0(_05501_),
    .A1(\fifo_bank_register.bank[4][110] ),
    .S(_07464_),
    .X(_07465_));
 sky130_fd_sc_hd__clkbuf_1 _12357_ (.A(_07465_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _12358_ (.A0(_05504_),
    .A1(\fifo_bank_register.bank[4][111] ),
    .S(_07464_),
    .X(_07466_));
 sky130_fd_sc_hd__clkbuf_1 _12359_ (.A(_07466_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _12360_ (.A0(_05506_),
    .A1(\fifo_bank_register.bank[4][112] ),
    .S(_07464_),
    .X(_07467_));
 sky130_fd_sc_hd__clkbuf_1 _12361_ (.A(_07467_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _12362_ (.A0(_05508_),
    .A1(\fifo_bank_register.bank[4][113] ),
    .S(_07464_),
    .X(_07468_));
 sky130_fd_sc_hd__clkbuf_1 _12363_ (.A(_07468_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _12364_ (.A0(_05510_),
    .A1(\fifo_bank_register.bank[4][114] ),
    .S(_07464_),
    .X(_07469_));
 sky130_fd_sc_hd__clkbuf_1 _12365_ (.A(_07469_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _12366_ (.A0(_05512_),
    .A1(\fifo_bank_register.bank[4][115] ),
    .S(_07464_),
    .X(_07470_));
 sky130_fd_sc_hd__clkbuf_1 _12367_ (.A(_07470_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _12368_ (.A0(_05514_),
    .A1(\fifo_bank_register.bank[4][116] ),
    .S(_07464_),
    .X(_07471_));
 sky130_fd_sc_hd__clkbuf_1 _12369_ (.A(_07471_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _12370_ (.A0(_05516_),
    .A1(\fifo_bank_register.bank[4][117] ),
    .S(_07464_),
    .X(_07472_));
 sky130_fd_sc_hd__clkbuf_1 _12371_ (.A(_07472_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(_05518_),
    .A1(\fifo_bank_register.bank[4][118] ),
    .S(_07464_),
    .X(_07473_));
 sky130_fd_sc_hd__clkbuf_1 _12373_ (.A(_07473_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(_05520_),
    .A1(\fifo_bank_register.bank[4][119] ),
    .S(_07464_),
    .X(_07474_));
 sky130_fd_sc_hd__clkbuf_1 _12375_ (.A(_07474_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(_05522_),
    .A1(\fifo_bank_register.bank[4][120] ),
    .S(_07341_),
    .X(_07475_));
 sky130_fd_sc_hd__clkbuf_1 _12377_ (.A(_07475_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(_05524_),
    .A1(\fifo_bank_register.bank[4][121] ),
    .S(_07341_),
    .X(_07476_));
 sky130_fd_sc_hd__clkbuf_1 _12379_ (.A(_07476_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(_05526_),
    .A1(\fifo_bank_register.bank[4][122] ),
    .S(_07341_),
    .X(_07477_));
 sky130_fd_sc_hd__clkbuf_1 _12381_ (.A(_07477_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(_05528_),
    .A1(\fifo_bank_register.bank[4][123] ),
    .S(_07341_),
    .X(_07478_));
 sky130_fd_sc_hd__clkbuf_1 _12383_ (.A(_07478_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(_05530_),
    .A1(\fifo_bank_register.bank[4][124] ),
    .S(_07341_),
    .X(_07479_));
 sky130_fd_sc_hd__clkbuf_1 _12385_ (.A(_07479_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(_05532_),
    .A1(\fifo_bank_register.bank[4][125] ),
    .S(_07341_),
    .X(_07480_));
 sky130_fd_sc_hd__clkbuf_1 _12387_ (.A(_07480_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(_05534_),
    .A1(\fifo_bank_register.bank[4][126] ),
    .S(_07341_),
    .X(_07481_));
 sky130_fd_sc_hd__clkbuf_1 _12389_ (.A(_07481_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(_05536_),
    .A1(\fifo_bank_register.bank[4][127] ),
    .S(_07341_),
    .X(_07482_));
 sky130_fd_sc_hd__clkbuf_1 _12391_ (.A(_07482_),
    .X(_00920_));
 sky130_fd_sc_hd__and3b_1 _12392_ (.A_N(\fifo_bank_register.write_ptr[2] ),
    .B(_05254_),
    .C(_05266_),
    .X(_07483_));
 sky130_fd_sc_hd__and4_1 _12393_ (.A(net597),
    .B(_05249_),
    .C(_05250_),
    .D(_07483_),
    .X(_07484_));
 sky130_fd_sc_hd__buf_4 _12394_ (.A(_07484_),
    .X(_07485_));
 sky130_fd_sc_hd__buf_4 _12395_ (.A(_07485_),
    .X(_07486_));
 sky130_fd_sc_hd__mux2_1 _12396_ (.A0(\fifo_bank_register.bank[3][0] ),
    .A1(_05248_),
    .S(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__clkbuf_1 _12397_ (.A(_07487_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _12398_ (.A0(\fifo_bank_register.bank[3][1] ),
    .A1(_05272_),
    .S(_07486_),
    .X(_07488_));
 sky130_fd_sc_hd__clkbuf_1 _12399_ (.A(_07488_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _12400_ (.A0(\fifo_bank_register.bank[3][2] ),
    .A1(_05274_),
    .S(_07486_),
    .X(_07489_));
 sky130_fd_sc_hd__clkbuf_1 _12401_ (.A(_07489_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(\fifo_bank_register.bank[3][3] ),
    .A1(_05276_),
    .S(_07486_),
    .X(_07490_));
 sky130_fd_sc_hd__clkbuf_1 _12403_ (.A(_07490_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _12404_ (.A0(\fifo_bank_register.bank[3][4] ),
    .A1(_05278_),
    .S(_07486_),
    .X(_07491_));
 sky130_fd_sc_hd__clkbuf_1 _12405_ (.A(_07491_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _12406_ (.A0(\fifo_bank_register.bank[3][5] ),
    .A1(_05280_),
    .S(_07486_),
    .X(_07492_));
 sky130_fd_sc_hd__clkbuf_1 _12407_ (.A(_07492_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _12408_ (.A0(\fifo_bank_register.bank[3][6] ),
    .A1(_05282_),
    .S(_07486_),
    .X(_07493_));
 sky130_fd_sc_hd__clkbuf_1 _12409_ (.A(_07493_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(\fifo_bank_register.bank[3][7] ),
    .A1(_05284_),
    .S(_07486_),
    .X(_07494_));
 sky130_fd_sc_hd__clkbuf_1 _12411_ (.A(_07494_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _12412_ (.A0(\fifo_bank_register.bank[3][8] ),
    .A1(_05286_),
    .S(_07486_),
    .X(_07495_));
 sky130_fd_sc_hd__clkbuf_1 _12413_ (.A(_07495_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _12414_ (.A0(\fifo_bank_register.bank[3][9] ),
    .A1(_05288_),
    .S(_07486_),
    .X(_07496_));
 sky130_fd_sc_hd__clkbuf_1 _12415_ (.A(_07496_),
    .X(_00930_));
 sky130_fd_sc_hd__buf_4 _12416_ (.A(_07485_),
    .X(_07497_));
 sky130_fd_sc_hd__mux2_1 _12417_ (.A0(\fifo_bank_register.bank[3][10] ),
    .A1(_05290_),
    .S(_07497_),
    .X(_07498_));
 sky130_fd_sc_hd__clkbuf_1 _12418_ (.A(_07498_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _12419_ (.A0(\fifo_bank_register.bank[3][11] ),
    .A1(_05293_),
    .S(_07497_),
    .X(_07499_));
 sky130_fd_sc_hd__clkbuf_1 _12420_ (.A(_07499_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _12421_ (.A0(\fifo_bank_register.bank[3][12] ),
    .A1(_05295_),
    .S(_07497_),
    .X(_07500_));
 sky130_fd_sc_hd__clkbuf_1 _12422_ (.A(_07500_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _12423_ (.A0(\fifo_bank_register.bank[3][13] ),
    .A1(_05297_),
    .S(_07497_),
    .X(_07501_));
 sky130_fd_sc_hd__clkbuf_1 _12424_ (.A(_07501_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _12425_ (.A0(\fifo_bank_register.bank[3][14] ),
    .A1(_05299_),
    .S(_07497_),
    .X(_07502_));
 sky130_fd_sc_hd__clkbuf_1 _12426_ (.A(_07502_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _12427_ (.A0(\fifo_bank_register.bank[3][15] ),
    .A1(_05301_),
    .S(_07497_),
    .X(_07503_));
 sky130_fd_sc_hd__clkbuf_1 _12428_ (.A(_07503_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _12429_ (.A0(\fifo_bank_register.bank[3][16] ),
    .A1(_05303_),
    .S(_07497_),
    .X(_07504_));
 sky130_fd_sc_hd__clkbuf_1 _12430_ (.A(_07504_),
    .X(_00937_));
 sky130_fd_sc_hd__mux2_1 _12431_ (.A0(\fifo_bank_register.bank[3][17] ),
    .A1(_05305_),
    .S(_07497_),
    .X(_07505_));
 sky130_fd_sc_hd__clkbuf_1 _12432_ (.A(_07505_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _12433_ (.A0(\fifo_bank_register.bank[3][18] ),
    .A1(_05307_),
    .S(_07497_),
    .X(_07506_));
 sky130_fd_sc_hd__clkbuf_1 _12434_ (.A(_07506_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _12435_ (.A0(\fifo_bank_register.bank[3][19] ),
    .A1(_05309_),
    .S(_07497_),
    .X(_07507_));
 sky130_fd_sc_hd__clkbuf_1 _12436_ (.A(_07507_),
    .X(_00940_));
 sky130_fd_sc_hd__buf_6 _12437_ (.A(_07484_),
    .X(_07508_));
 sky130_fd_sc_hd__clkbuf_4 _12438_ (.A(_07508_),
    .X(_07509_));
 sky130_fd_sc_hd__mux2_1 _12439_ (.A0(\fifo_bank_register.bank[3][20] ),
    .A1(_05311_),
    .S(_07509_),
    .X(_07510_));
 sky130_fd_sc_hd__clkbuf_1 _12440_ (.A(_07510_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _12441_ (.A0(\fifo_bank_register.bank[3][21] ),
    .A1(_05315_),
    .S(_07509_),
    .X(_07511_));
 sky130_fd_sc_hd__clkbuf_1 _12442_ (.A(_07511_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _12443_ (.A0(\fifo_bank_register.bank[3][22] ),
    .A1(_05317_),
    .S(_07509_),
    .X(_07512_));
 sky130_fd_sc_hd__clkbuf_1 _12444_ (.A(_07512_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _12445_ (.A0(\fifo_bank_register.bank[3][23] ),
    .A1(_05319_),
    .S(_07509_),
    .X(_07513_));
 sky130_fd_sc_hd__clkbuf_1 _12446_ (.A(_07513_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _12447_ (.A0(\fifo_bank_register.bank[3][24] ),
    .A1(_05321_),
    .S(_07509_),
    .X(_07514_));
 sky130_fd_sc_hd__clkbuf_1 _12448_ (.A(_07514_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _12449_ (.A0(\fifo_bank_register.bank[3][25] ),
    .A1(_05323_),
    .S(_07509_),
    .X(_07515_));
 sky130_fd_sc_hd__clkbuf_1 _12450_ (.A(_07515_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(\fifo_bank_register.bank[3][26] ),
    .A1(_05325_),
    .S(_07509_),
    .X(_07516_));
 sky130_fd_sc_hd__clkbuf_1 _12452_ (.A(_07516_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(\fifo_bank_register.bank[3][27] ),
    .A1(_05327_),
    .S(_07509_),
    .X(_07517_));
 sky130_fd_sc_hd__clkbuf_1 _12454_ (.A(_07517_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(\fifo_bank_register.bank[3][28] ),
    .A1(_05329_),
    .S(_07509_),
    .X(_07518_));
 sky130_fd_sc_hd__clkbuf_1 _12456_ (.A(_07518_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _12457_ (.A0(\fifo_bank_register.bank[3][29] ),
    .A1(_05331_),
    .S(_07509_),
    .X(_07519_));
 sky130_fd_sc_hd__clkbuf_1 _12458_ (.A(_07519_),
    .X(_00950_));
 sky130_fd_sc_hd__buf_4 _12459_ (.A(_07508_),
    .X(_07520_));
 sky130_fd_sc_hd__mux2_1 _12460_ (.A0(\fifo_bank_register.bank[3][30] ),
    .A1(_05333_),
    .S(_07520_),
    .X(_07521_));
 sky130_fd_sc_hd__clkbuf_1 _12461_ (.A(_07521_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _12462_ (.A0(\fifo_bank_register.bank[3][31] ),
    .A1(_05336_),
    .S(_07520_),
    .X(_07522_));
 sky130_fd_sc_hd__clkbuf_1 _12463_ (.A(_07522_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _12464_ (.A0(\fifo_bank_register.bank[3][32] ),
    .A1(_05338_),
    .S(_07520_),
    .X(_07523_));
 sky130_fd_sc_hd__clkbuf_1 _12465_ (.A(_07523_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _12466_ (.A0(\fifo_bank_register.bank[3][33] ),
    .A1(_05340_),
    .S(_07520_),
    .X(_07524_));
 sky130_fd_sc_hd__clkbuf_1 _12467_ (.A(_07524_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _12468_ (.A0(\fifo_bank_register.bank[3][34] ),
    .A1(_05342_),
    .S(_07520_),
    .X(_07525_));
 sky130_fd_sc_hd__clkbuf_1 _12469_ (.A(_07525_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(\fifo_bank_register.bank[3][35] ),
    .A1(_05344_),
    .S(_07520_),
    .X(_07526_));
 sky130_fd_sc_hd__clkbuf_1 _12471_ (.A(_07526_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(\fifo_bank_register.bank[3][36] ),
    .A1(_05346_),
    .S(_07520_),
    .X(_07527_));
 sky130_fd_sc_hd__clkbuf_1 _12473_ (.A(_07527_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _12474_ (.A0(\fifo_bank_register.bank[3][37] ),
    .A1(_05348_),
    .S(_07520_),
    .X(_07528_));
 sky130_fd_sc_hd__clkbuf_1 _12475_ (.A(_07528_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(\fifo_bank_register.bank[3][38] ),
    .A1(_05350_),
    .S(_07520_),
    .X(_07529_));
 sky130_fd_sc_hd__clkbuf_1 _12477_ (.A(_07529_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _12478_ (.A0(\fifo_bank_register.bank[3][39] ),
    .A1(_05352_),
    .S(_07520_),
    .X(_07530_));
 sky130_fd_sc_hd__clkbuf_1 _12479_ (.A(_07530_),
    .X(_00960_));
 sky130_fd_sc_hd__buf_4 _12480_ (.A(_07508_),
    .X(_07531_));
 sky130_fd_sc_hd__mux2_1 _12481_ (.A0(\fifo_bank_register.bank[3][40] ),
    .A1(_05354_),
    .S(_07531_),
    .X(_07532_));
 sky130_fd_sc_hd__clkbuf_1 _12482_ (.A(_07532_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _12483_ (.A0(\fifo_bank_register.bank[3][41] ),
    .A1(_05357_),
    .S(_07531_),
    .X(_07533_));
 sky130_fd_sc_hd__clkbuf_1 _12484_ (.A(_07533_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _12485_ (.A0(\fifo_bank_register.bank[3][42] ),
    .A1(_05359_),
    .S(_07531_),
    .X(_07534_));
 sky130_fd_sc_hd__clkbuf_1 _12486_ (.A(_07534_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _12487_ (.A0(\fifo_bank_register.bank[3][43] ),
    .A1(_05361_),
    .S(_07531_),
    .X(_07535_));
 sky130_fd_sc_hd__clkbuf_1 _12488_ (.A(_07535_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _12489_ (.A0(\fifo_bank_register.bank[3][44] ),
    .A1(_05363_),
    .S(_07531_),
    .X(_07536_));
 sky130_fd_sc_hd__clkbuf_1 _12490_ (.A(_07536_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _12491_ (.A0(\fifo_bank_register.bank[3][45] ),
    .A1(_05365_),
    .S(_07531_),
    .X(_07537_));
 sky130_fd_sc_hd__clkbuf_1 _12492_ (.A(_07537_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _12493_ (.A0(\fifo_bank_register.bank[3][46] ),
    .A1(_05367_),
    .S(_07531_),
    .X(_07538_));
 sky130_fd_sc_hd__clkbuf_1 _12494_ (.A(_07538_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _12495_ (.A0(\fifo_bank_register.bank[3][47] ),
    .A1(_05369_),
    .S(_07531_),
    .X(_07539_));
 sky130_fd_sc_hd__clkbuf_1 _12496_ (.A(_07539_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _12497_ (.A0(\fifo_bank_register.bank[3][48] ),
    .A1(_05371_),
    .S(_07531_),
    .X(_07540_));
 sky130_fd_sc_hd__clkbuf_1 _12498_ (.A(_07540_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(\fifo_bank_register.bank[3][49] ),
    .A1(_05373_),
    .S(_07531_),
    .X(_07541_));
 sky130_fd_sc_hd__clkbuf_1 _12500_ (.A(_07541_),
    .X(_00970_));
 sky130_fd_sc_hd__buf_4 _12501_ (.A(_07508_),
    .X(_07542_));
 sky130_fd_sc_hd__mux2_1 _12502_ (.A0(\fifo_bank_register.bank[3][50] ),
    .A1(_05375_),
    .S(_07542_),
    .X(_07543_));
 sky130_fd_sc_hd__clkbuf_1 _12503_ (.A(_07543_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _12504_ (.A0(\fifo_bank_register.bank[3][51] ),
    .A1(_05378_),
    .S(_07542_),
    .X(_07544_));
 sky130_fd_sc_hd__clkbuf_1 _12505_ (.A(_07544_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _12506_ (.A0(\fifo_bank_register.bank[3][52] ),
    .A1(_05380_),
    .S(_07542_),
    .X(_07545_));
 sky130_fd_sc_hd__clkbuf_1 _12507_ (.A(_07545_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _12508_ (.A0(\fifo_bank_register.bank[3][53] ),
    .A1(_05382_),
    .S(_07542_),
    .X(_07546_));
 sky130_fd_sc_hd__clkbuf_1 _12509_ (.A(_07546_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _12510_ (.A0(\fifo_bank_register.bank[3][54] ),
    .A1(_05384_),
    .S(_07542_),
    .X(_07547_));
 sky130_fd_sc_hd__clkbuf_1 _12511_ (.A(_07547_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _12512_ (.A0(\fifo_bank_register.bank[3][55] ),
    .A1(_05386_),
    .S(_07542_),
    .X(_07548_));
 sky130_fd_sc_hd__clkbuf_1 _12513_ (.A(_07548_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _12514_ (.A0(\fifo_bank_register.bank[3][56] ),
    .A1(_05388_),
    .S(_07542_),
    .X(_07549_));
 sky130_fd_sc_hd__clkbuf_1 _12515_ (.A(_07549_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _12516_ (.A0(\fifo_bank_register.bank[3][57] ),
    .A1(_05390_),
    .S(_07542_),
    .X(_07550_));
 sky130_fd_sc_hd__clkbuf_1 _12517_ (.A(_07550_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _12518_ (.A0(\fifo_bank_register.bank[3][58] ),
    .A1(_05392_),
    .S(_07542_),
    .X(_07551_));
 sky130_fd_sc_hd__clkbuf_1 _12519_ (.A(_07551_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _12520_ (.A0(\fifo_bank_register.bank[3][59] ),
    .A1(_05394_),
    .S(_07542_),
    .X(_07552_));
 sky130_fd_sc_hd__clkbuf_1 _12521_ (.A(_07552_),
    .X(_00980_));
 sky130_fd_sc_hd__buf_4 _12522_ (.A(_07508_),
    .X(_07553_));
 sky130_fd_sc_hd__mux2_1 _12523_ (.A0(\fifo_bank_register.bank[3][60] ),
    .A1(_05396_),
    .S(_07553_),
    .X(_07554_));
 sky130_fd_sc_hd__clkbuf_1 _12524_ (.A(_07554_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _12525_ (.A0(\fifo_bank_register.bank[3][61] ),
    .A1(_05399_),
    .S(_07553_),
    .X(_07555_));
 sky130_fd_sc_hd__clkbuf_1 _12526_ (.A(_07555_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _12527_ (.A0(\fifo_bank_register.bank[3][62] ),
    .A1(_05401_),
    .S(_07553_),
    .X(_07556_));
 sky130_fd_sc_hd__clkbuf_1 _12528_ (.A(_07556_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _12529_ (.A0(\fifo_bank_register.bank[3][63] ),
    .A1(_05403_),
    .S(_07553_),
    .X(_07557_));
 sky130_fd_sc_hd__clkbuf_1 _12530_ (.A(_07557_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _12531_ (.A0(\fifo_bank_register.bank[3][64] ),
    .A1(_05405_),
    .S(_07553_),
    .X(_07558_));
 sky130_fd_sc_hd__clkbuf_1 _12532_ (.A(_07558_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _12533_ (.A0(\fifo_bank_register.bank[3][65] ),
    .A1(_05407_),
    .S(_07553_),
    .X(_07559_));
 sky130_fd_sc_hd__clkbuf_1 _12534_ (.A(_07559_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _12535_ (.A0(\fifo_bank_register.bank[3][66] ),
    .A1(_05409_),
    .S(_07553_),
    .X(_07560_));
 sky130_fd_sc_hd__clkbuf_1 _12536_ (.A(_07560_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _12537_ (.A0(\fifo_bank_register.bank[3][67] ),
    .A1(_05411_),
    .S(_07553_),
    .X(_07561_));
 sky130_fd_sc_hd__clkbuf_1 _12538_ (.A(_07561_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(\fifo_bank_register.bank[3][68] ),
    .A1(_05413_),
    .S(_07553_),
    .X(_07562_));
 sky130_fd_sc_hd__clkbuf_1 _12540_ (.A(_07562_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(\fifo_bank_register.bank[3][69] ),
    .A1(_05415_),
    .S(_07553_),
    .X(_07563_));
 sky130_fd_sc_hd__clkbuf_1 _12542_ (.A(_07563_),
    .X(_00990_));
 sky130_fd_sc_hd__clkbuf_4 _12543_ (.A(_07508_),
    .X(_07564_));
 sky130_fd_sc_hd__mux2_1 _12544_ (.A0(\fifo_bank_register.bank[3][70] ),
    .A1(_05417_),
    .S(_07564_),
    .X(_07565_));
 sky130_fd_sc_hd__clkbuf_1 _12545_ (.A(_07565_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _12546_ (.A0(\fifo_bank_register.bank[3][71] ),
    .A1(_05420_),
    .S(_07564_),
    .X(_07566_));
 sky130_fd_sc_hd__clkbuf_1 _12547_ (.A(_07566_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _12548_ (.A0(\fifo_bank_register.bank[3][72] ),
    .A1(_05422_),
    .S(_07564_),
    .X(_07567_));
 sky130_fd_sc_hd__clkbuf_1 _12549_ (.A(_07567_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _12550_ (.A0(\fifo_bank_register.bank[3][73] ),
    .A1(_05424_),
    .S(_07564_),
    .X(_07568_));
 sky130_fd_sc_hd__clkbuf_1 _12551_ (.A(_07568_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _12552_ (.A0(\fifo_bank_register.bank[3][74] ),
    .A1(_05426_),
    .S(_07564_),
    .X(_07569_));
 sky130_fd_sc_hd__clkbuf_1 _12553_ (.A(_07569_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _12554_ (.A0(\fifo_bank_register.bank[3][75] ),
    .A1(_05428_),
    .S(_07564_),
    .X(_07570_));
 sky130_fd_sc_hd__clkbuf_1 _12555_ (.A(_07570_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _12556_ (.A0(\fifo_bank_register.bank[3][76] ),
    .A1(_05430_),
    .S(_07564_),
    .X(_07571_));
 sky130_fd_sc_hd__clkbuf_1 _12557_ (.A(_07571_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _12558_ (.A0(\fifo_bank_register.bank[3][77] ),
    .A1(_05432_),
    .S(_07564_),
    .X(_07572_));
 sky130_fd_sc_hd__clkbuf_1 _12559_ (.A(_07572_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _12560_ (.A0(\fifo_bank_register.bank[3][78] ),
    .A1(_05434_),
    .S(_07564_),
    .X(_07573_));
 sky130_fd_sc_hd__clkbuf_1 _12561_ (.A(_07573_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(\fifo_bank_register.bank[3][79] ),
    .A1(_05436_),
    .S(_07564_),
    .X(_07574_));
 sky130_fd_sc_hd__clkbuf_1 _12563_ (.A(_07574_),
    .X(_01000_));
 sky130_fd_sc_hd__clkbuf_4 _12564_ (.A(_07508_),
    .X(_07575_));
 sky130_fd_sc_hd__mux2_1 _12565_ (.A0(\fifo_bank_register.bank[3][80] ),
    .A1(_05438_),
    .S(_07575_),
    .X(_07576_));
 sky130_fd_sc_hd__clkbuf_1 _12566_ (.A(_07576_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _12567_ (.A0(\fifo_bank_register.bank[3][81] ),
    .A1(_05441_),
    .S(_07575_),
    .X(_07577_));
 sky130_fd_sc_hd__clkbuf_1 _12568_ (.A(_07577_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _12569_ (.A0(\fifo_bank_register.bank[3][82] ),
    .A1(_05443_),
    .S(_07575_),
    .X(_07578_));
 sky130_fd_sc_hd__clkbuf_1 _12570_ (.A(_07578_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _12571_ (.A0(\fifo_bank_register.bank[3][83] ),
    .A1(_05445_),
    .S(_07575_),
    .X(_07579_));
 sky130_fd_sc_hd__clkbuf_1 _12572_ (.A(_07579_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _12573_ (.A0(\fifo_bank_register.bank[3][84] ),
    .A1(_05447_),
    .S(_07575_),
    .X(_07580_));
 sky130_fd_sc_hd__clkbuf_1 _12574_ (.A(_07580_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _12575_ (.A0(\fifo_bank_register.bank[3][85] ),
    .A1(_05449_),
    .S(_07575_),
    .X(_07581_));
 sky130_fd_sc_hd__clkbuf_1 _12576_ (.A(_07581_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _12577_ (.A0(\fifo_bank_register.bank[3][86] ),
    .A1(_05451_),
    .S(_07575_),
    .X(_07582_));
 sky130_fd_sc_hd__clkbuf_1 _12578_ (.A(_07582_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _12579_ (.A0(\fifo_bank_register.bank[3][87] ),
    .A1(_05453_),
    .S(_07575_),
    .X(_07583_));
 sky130_fd_sc_hd__clkbuf_1 _12580_ (.A(_07583_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _12581_ (.A0(\fifo_bank_register.bank[3][88] ),
    .A1(_05455_),
    .S(_07575_),
    .X(_07584_));
 sky130_fd_sc_hd__clkbuf_1 _12582_ (.A(_07584_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _12583_ (.A0(\fifo_bank_register.bank[3][89] ),
    .A1(_05457_),
    .S(_07575_),
    .X(_07585_));
 sky130_fd_sc_hd__clkbuf_1 _12584_ (.A(_07585_),
    .X(_01010_));
 sky130_fd_sc_hd__buf_4 _12585_ (.A(_07508_),
    .X(_07586_));
 sky130_fd_sc_hd__mux2_1 _12586_ (.A0(\fifo_bank_register.bank[3][90] ),
    .A1(_05459_),
    .S(_07586_),
    .X(_07587_));
 sky130_fd_sc_hd__clkbuf_1 _12587_ (.A(_07587_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _12588_ (.A0(\fifo_bank_register.bank[3][91] ),
    .A1(_05462_),
    .S(_07586_),
    .X(_07588_));
 sky130_fd_sc_hd__clkbuf_1 _12589_ (.A(_07588_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _12590_ (.A0(\fifo_bank_register.bank[3][92] ),
    .A1(_05464_),
    .S(_07586_),
    .X(_07589_));
 sky130_fd_sc_hd__clkbuf_1 _12591_ (.A(_07589_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _12592_ (.A0(\fifo_bank_register.bank[3][93] ),
    .A1(_05466_),
    .S(_07586_),
    .X(_07590_));
 sky130_fd_sc_hd__clkbuf_1 _12593_ (.A(_07590_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _12594_ (.A0(\fifo_bank_register.bank[3][94] ),
    .A1(_05468_),
    .S(_07586_),
    .X(_07591_));
 sky130_fd_sc_hd__clkbuf_1 _12595_ (.A(_07591_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(\fifo_bank_register.bank[3][95] ),
    .A1(_05470_),
    .S(_07586_),
    .X(_07592_));
 sky130_fd_sc_hd__clkbuf_1 _12597_ (.A(_07592_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(\fifo_bank_register.bank[3][96] ),
    .A1(_05472_),
    .S(_07586_),
    .X(_07593_));
 sky130_fd_sc_hd__clkbuf_1 _12599_ (.A(_07593_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(\fifo_bank_register.bank[3][97] ),
    .A1(_05474_),
    .S(_07586_),
    .X(_07594_));
 sky130_fd_sc_hd__clkbuf_1 _12601_ (.A(_07594_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(\fifo_bank_register.bank[3][98] ),
    .A1(_05476_),
    .S(_07586_),
    .X(_07595_));
 sky130_fd_sc_hd__clkbuf_1 _12603_ (.A(_07595_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _12604_ (.A0(\fifo_bank_register.bank[3][99] ),
    .A1(_05478_),
    .S(_07586_),
    .X(_07596_));
 sky130_fd_sc_hd__clkbuf_1 _12605_ (.A(_07596_),
    .X(_01020_));
 sky130_fd_sc_hd__buf_4 _12606_ (.A(_07508_),
    .X(_07597_));
 sky130_fd_sc_hd__mux2_1 _12607_ (.A0(\fifo_bank_register.bank[3][100] ),
    .A1(_05480_),
    .S(_07597_),
    .X(_07598_));
 sky130_fd_sc_hd__clkbuf_1 _12608_ (.A(_07598_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _12609_ (.A0(\fifo_bank_register.bank[3][101] ),
    .A1(_05483_),
    .S(_07597_),
    .X(_07599_));
 sky130_fd_sc_hd__clkbuf_1 _12610_ (.A(_07599_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _12611_ (.A0(\fifo_bank_register.bank[3][102] ),
    .A1(_05485_),
    .S(_07597_),
    .X(_07600_));
 sky130_fd_sc_hd__clkbuf_1 _12612_ (.A(_07600_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _12613_ (.A0(\fifo_bank_register.bank[3][103] ),
    .A1(_05487_),
    .S(_07597_),
    .X(_07601_));
 sky130_fd_sc_hd__clkbuf_1 _12614_ (.A(_07601_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _12615_ (.A0(\fifo_bank_register.bank[3][104] ),
    .A1(_05489_),
    .S(_07597_),
    .X(_07602_));
 sky130_fd_sc_hd__clkbuf_1 _12616_ (.A(_07602_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _12617_ (.A0(\fifo_bank_register.bank[3][105] ),
    .A1(_05491_),
    .S(_07597_),
    .X(_07603_));
 sky130_fd_sc_hd__clkbuf_1 _12618_ (.A(_07603_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _12619_ (.A0(\fifo_bank_register.bank[3][106] ),
    .A1(_05493_),
    .S(_07597_),
    .X(_07604_));
 sky130_fd_sc_hd__clkbuf_1 _12620_ (.A(_07604_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _12621_ (.A0(\fifo_bank_register.bank[3][107] ),
    .A1(_05495_),
    .S(_07597_),
    .X(_07605_));
 sky130_fd_sc_hd__clkbuf_1 _12622_ (.A(_07605_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _12623_ (.A0(\fifo_bank_register.bank[3][108] ),
    .A1(_05497_),
    .S(_07597_),
    .X(_07606_));
 sky130_fd_sc_hd__clkbuf_1 _12624_ (.A(_07606_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _12625_ (.A0(\fifo_bank_register.bank[3][109] ),
    .A1(_05499_),
    .S(_07597_),
    .X(_07607_));
 sky130_fd_sc_hd__clkbuf_1 _12626_ (.A(_07607_),
    .X(_01030_));
 sky130_fd_sc_hd__clkbuf_4 _12627_ (.A(_07508_),
    .X(_07608_));
 sky130_fd_sc_hd__mux2_1 _12628_ (.A0(\fifo_bank_register.bank[3][110] ),
    .A1(_05501_),
    .S(_07608_),
    .X(_07609_));
 sky130_fd_sc_hd__clkbuf_1 _12629_ (.A(_07609_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _12630_ (.A0(\fifo_bank_register.bank[3][111] ),
    .A1(_05504_),
    .S(_07608_),
    .X(_07610_));
 sky130_fd_sc_hd__clkbuf_1 _12631_ (.A(_07610_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _12632_ (.A0(\fifo_bank_register.bank[3][112] ),
    .A1(_05506_),
    .S(_07608_),
    .X(_07611_));
 sky130_fd_sc_hd__clkbuf_1 _12633_ (.A(_07611_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _12634_ (.A0(\fifo_bank_register.bank[3][113] ),
    .A1(_05508_),
    .S(_07608_),
    .X(_07612_));
 sky130_fd_sc_hd__clkbuf_1 _12635_ (.A(_07612_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _12636_ (.A0(\fifo_bank_register.bank[3][114] ),
    .A1(_05510_),
    .S(_07608_),
    .X(_07613_));
 sky130_fd_sc_hd__clkbuf_1 _12637_ (.A(_07613_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _12638_ (.A0(\fifo_bank_register.bank[3][115] ),
    .A1(_05512_),
    .S(_07608_),
    .X(_07614_));
 sky130_fd_sc_hd__clkbuf_1 _12639_ (.A(_07614_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _12640_ (.A0(\fifo_bank_register.bank[3][116] ),
    .A1(_05514_),
    .S(_07608_),
    .X(_07615_));
 sky130_fd_sc_hd__clkbuf_1 _12641_ (.A(_07615_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _12642_ (.A0(\fifo_bank_register.bank[3][117] ),
    .A1(_05516_),
    .S(_07608_),
    .X(_07616_));
 sky130_fd_sc_hd__clkbuf_1 _12643_ (.A(_07616_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _12644_ (.A0(\fifo_bank_register.bank[3][118] ),
    .A1(_05518_),
    .S(_07608_),
    .X(_07617_));
 sky130_fd_sc_hd__clkbuf_1 _12645_ (.A(_07617_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _12646_ (.A0(\fifo_bank_register.bank[3][119] ),
    .A1(_05520_),
    .S(_07608_),
    .X(_07618_));
 sky130_fd_sc_hd__clkbuf_1 _12647_ (.A(_07618_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _12648_ (.A0(\fifo_bank_register.bank[3][120] ),
    .A1(_05522_),
    .S(_07485_),
    .X(_07619_));
 sky130_fd_sc_hd__clkbuf_1 _12649_ (.A(_07619_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _12650_ (.A0(\fifo_bank_register.bank[3][121] ),
    .A1(_05524_),
    .S(_07485_),
    .X(_07620_));
 sky130_fd_sc_hd__clkbuf_1 _12651_ (.A(_07620_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(\fifo_bank_register.bank[3][122] ),
    .A1(_05526_),
    .S(_07485_),
    .X(_07621_));
 sky130_fd_sc_hd__clkbuf_1 _12653_ (.A(_07621_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _12654_ (.A0(\fifo_bank_register.bank[3][123] ),
    .A1(_05528_),
    .S(_07485_),
    .X(_07622_));
 sky130_fd_sc_hd__clkbuf_1 _12655_ (.A(_07622_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _12656_ (.A0(\fifo_bank_register.bank[3][124] ),
    .A1(_05530_),
    .S(_07485_),
    .X(_07623_));
 sky130_fd_sc_hd__clkbuf_1 _12657_ (.A(_07623_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _12658_ (.A0(\fifo_bank_register.bank[3][125] ),
    .A1(_05532_),
    .S(_07485_),
    .X(_07624_));
 sky130_fd_sc_hd__clkbuf_1 _12659_ (.A(_07624_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _12660_ (.A0(\fifo_bank_register.bank[3][126] ),
    .A1(_05534_),
    .S(_07485_),
    .X(_07625_));
 sky130_fd_sc_hd__clkbuf_1 _12661_ (.A(_07625_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _12662_ (.A0(\fifo_bank_register.bank[3][127] ),
    .A1(_05536_),
    .S(_07485_),
    .X(_07626_));
 sky130_fd_sc_hd__clkbuf_1 _12663_ (.A(_07626_),
    .X(_01048_));
 sky130_fd_sc_hd__and4b_1 _12664_ (.A_N(_05249_),
    .B(_05250_),
    .C(_07483_),
    .D(net597),
    .X(_07627_));
 sky130_fd_sc_hd__buf_4 _12665_ (.A(_07627_),
    .X(_07628_));
 sky130_fd_sc_hd__buf_4 _12666_ (.A(_07628_),
    .X(_07629_));
 sky130_fd_sc_hd__mux2_1 _12667_ (.A0(\fifo_bank_register.bank[2][0] ),
    .A1(_05248_),
    .S(_07629_),
    .X(_07630_));
 sky130_fd_sc_hd__clkbuf_1 _12668_ (.A(_07630_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _12669_ (.A0(\fifo_bank_register.bank[2][1] ),
    .A1(_05272_),
    .S(_07629_),
    .X(_07631_));
 sky130_fd_sc_hd__clkbuf_1 _12670_ (.A(_07631_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _12671_ (.A0(\fifo_bank_register.bank[2][2] ),
    .A1(_05274_),
    .S(_07629_),
    .X(_07632_));
 sky130_fd_sc_hd__clkbuf_1 _12672_ (.A(_07632_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _12673_ (.A0(\fifo_bank_register.bank[2][3] ),
    .A1(_05276_),
    .S(_07629_),
    .X(_07633_));
 sky130_fd_sc_hd__clkbuf_1 _12674_ (.A(_07633_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _12675_ (.A0(\fifo_bank_register.bank[2][4] ),
    .A1(_05278_),
    .S(_07629_),
    .X(_07634_));
 sky130_fd_sc_hd__clkbuf_1 _12676_ (.A(_07634_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _12677_ (.A0(\fifo_bank_register.bank[2][5] ),
    .A1(_05280_),
    .S(_07629_),
    .X(_07635_));
 sky130_fd_sc_hd__clkbuf_1 _12678_ (.A(_07635_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _12679_ (.A0(\fifo_bank_register.bank[2][6] ),
    .A1(_05282_),
    .S(_07629_),
    .X(_07636_));
 sky130_fd_sc_hd__clkbuf_1 _12680_ (.A(_07636_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _12681_ (.A0(\fifo_bank_register.bank[2][7] ),
    .A1(_05284_),
    .S(_07629_),
    .X(_07637_));
 sky130_fd_sc_hd__clkbuf_1 _12682_ (.A(_07637_),
    .X(_01056_));
 sky130_fd_sc_hd__mux2_1 _12683_ (.A0(\fifo_bank_register.bank[2][8] ),
    .A1(_05286_),
    .S(_07629_),
    .X(_07638_));
 sky130_fd_sc_hd__clkbuf_1 _12684_ (.A(_07638_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _12685_ (.A0(\fifo_bank_register.bank[2][9] ),
    .A1(_05288_),
    .S(_07629_),
    .X(_07639_));
 sky130_fd_sc_hd__clkbuf_1 _12686_ (.A(_07639_),
    .X(_01058_));
 sky130_fd_sc_hd__buf_4 _12687_ (.A(_07628_),
    .X(_07640_));
 sky130_fd_sc_hd__mux2_1 _12688_ (.A0(\fifo_bank_register.bank[2][10] ),
    .A1(_05290_),
    .S(_07640_),
    .X(_07641_));
 sky130_fd_sc_hd__clkbuf_1 _12689_ (.A(_07641_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _12690_ (.A0(\fifo_bank_register.bank[2][11] ),
    .A1(_05293_),
    .S(_07640_),
    .X(_07642_));
 sky130_fd_sc_hd__clkbuf_1 _12691_ (.A(_07642_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _12692_ (.A0(\fifo_bank_register.bank[2][12] ),
    .A1(_05295_),
    .S(_07640_),
    .X(_07643_));
 sky130_fd_sc_hd__clkbuf_1 _12693_ (.A(_07643_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _12694_ (.A0(\fifo_bank_register.bank[2][13] ),
    .A1(_05297_),
    .S(_07640_),
    .X(_07644_));
 sky130_fd_sc_hd__clkbuf_1 _12695_ (.A(_07644_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _12696_ (.A0(\fifo_bank_register.bank[2][14] ),
    .A1(_05299_),
    .S(_07640_),
    .X(_07645_));
 sky130_fd_sc_hd__clkbuf_1 _12697_ (.A(_07645_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _12698_ (.A0(\fifo_bank_register.bank[2][15] ),
    .A1(_05301_),
    .S(_07640_),
    .X(_07646_));
 sky130_fd_sc_hd__clkbuf_1 _12699_ (.A(_07646_),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _12700_ (.A0(\fifo_bank_register.bank[2][16] ),
    .A1(_05303_),
    .S(_07640_),
    .X(_07647_));
 sky130_fd_sc_hd__clkbuf_1 _12701_ (.A(_07647_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _12702_ (.A0(\fifo_bank_register.bank[2][17] ),
    .A1(_05305_),
    .S(_07640_),
    .X(_07648_));
 sky130_fd_sc_hd__clkbuf_1 _12703_ (.A(_07648_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _12704_ (.A0(\fifo_bank_register.bank[2][18] ),
    .A1(_05307_),
    .S(_07640_),
    .X(_07649_));
 sky130_fd_sc_hd__clkbuf_1 _12705_ (.A(_07649_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _12706_ (.A0(\fifo_bank_register.bank[2][19] ),
    .A1(_05309_),
    .S(_07640_),
    .X(_07650_));
 sky130_fd_sc_hd__clkbuf_1 _12707_ (.A(_07650_),
    .X(_01068_));
 sky130_fd_sc_hd__buf_6 _12708_ (.A(_07627_),
    .X(_07651_));
 sky130_fd_sc_hd__buf_4 _12709_ (.A(_07651_),
    .X(_07652_));
 sky130_fd_sc_hd__mux2_1 _12710_ (.A0(\fifo_bank_register.bank[2][20] ),
    .A1(_05311_),
    .S(_07652_),
    .X(_07653_));
 sky130_fd_sc_hd__clkbuf_1 _12711_ (.A(_07653_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _12712_ (.A0(\fifo_bank_register.bank[2][21] ),
    .A1(_05315_),
    .S(_07652_),
    .X(_07654_));
 sky130_fd_sc_hd__clkbuf_1 _12713_ (.A(_07654_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(\fifo_bank_register.bank[2][22] ),
    .A1(_05317_),
    .S(_07652_),
    .X(_07655_));
 sky130_fd_sc_hd__clkbuf_1 _12715_ (.A(_07655_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _12716_ (.A0(\fifo_bank_register.bank[2][23] ),
    .A1(_05319_),
    .S(_07652_),
    .X(_07656_));
 sky130_fd_sc_hd__clkbuf_1 _12717_ (.A(_07656_),
    .X(_01072_));
 sky130_fd_sc_hd__mux2_1 _12718_ (.A0(\fifo_bank_register.bank[2][24] ),
    .A1(_05321_),
    .S(_07652_),
    .X(_07657_));
 sky130_fd_sc_hd__clkbuf_1 _12719_ (.A(_07657_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _12720_ (.A0(\fifo_bank_register.bank[2][25] ),
    .A1(_05323_),
    .S(_07652_),
    .X(_07658_));
 sky130_fd_sc_hd__clkbuf_1 _12721_ (.A(_07658_),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _12722_ (.A0(\fifo_bank_register.bank[2][26] ),
    .A1(_05325_),
    .S(_07652_),
    .X(_07659_));
 sky130_fd_sc_hd__clkbuf_1 _12723_ (.A(_07659_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _12724_ (.A0(\fifo_bank_register.bank[2][27] ),
    .A1(_05327_),
    .S(_07652_),
    .X(_07660_));
 sky130_fd_sc_hd__clkbuf_1 _12725_ (.A(_07660_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _12726_ (.A0(\fifo_bank_register.bank[2][28] ),
    .A1(_05329_),
    .S(_07652_),
    .X(_07661_));
 sky130_fd_sc_hd__clkbuf_1 _12727_ (.A(_07661_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _12728_ (.A0(\fifo_bank_register.bank[2][29] ),
    .A1(_05331_),
    .S(_07652_),
    .X(_07662_));
 sky130_fd_sc_hd__clkbuf_1 _12729_ (.A(_07662_),
    .X(_01078_));
 sky130_fd_sc_hd__buf_4 _12730_ (.A(_07651_),
    .X(_07663_));
 sky130_fd_sc_hd__mux2_1 _12731_ (.A0(\fifo_bank_register.bank[2][30] ),
    .A1(_05333_),
    .S(_07663_),
    .X(_07664_));
 sky130_fd_sc_hd__clkbuf_1 _12732_ (.A(_07664_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _12733_ (.A0(\fifo_bank_register.bank[2][31] ),
    .A1(_05336_),
    .S(_07663_),
    .X(_07665_));
 sky130_fd_sc_hd__clkbuf_1 _12734_ (.A(_07665_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _12735_ (.A0(\fifo_bank_register.bank[2][32] ),
    .A1(_05338_),
    .S(_07663_),
    .X(_07666_));
 sky130_fd_sc_hd__clkbuf_1 _12736_ (.A(_07666_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _12737_ (.A0(\fifo_bank_register.bank[2][33] ),
    .A1(_05340_),
    .S(_07663_),
    .X(_07667_));
 sky130_fd_sc_hd__clkbuf_1 _12738_ (.A(_07667_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _12739_ (.A0(\fifo_bank_register.bank[2][34] ),
    .A1(_05342_),
    .S(_07663_),
    .X(_07668_));
 sky130_fd_sc_hd__clkbuf_1 _12740_ (.A(_07668_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _12741_ (.A0(\fifo_bank_register.bank[2][35] ),
    .A1(_05344_),
    .S(_07663_),
    .X(_07669_));
 sky130_fd_sc_hd__clkbuf_1 _12742_ (.A(_07669_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _12743_ (.A0(\fifo_bank_register.bank[2][36] ),
    .A1(_05346_),
    .S(_07663_),
    .X(_07670_));
 sky130_fd_sc_hd__clkbuf_1 _12744_ (.A(_07670_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _12745_ (.A0(\fifo_bank_register.bank[2][37] ),
    .A1(_05348_),
    .S(_07663_),
    .X(_07671_));
 sky130_fd_sc_hd__clkbuf_1 _12746_ (.A(_07671_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _12747_ (.A0(\fifo_bank_register.bank[2][38] ),
    .A1(_05350_),
    .S(_07663_),
    .X(_07672_));
 sky130_fd_sc_hd__clkbuf_1 _12748_ (.A(_07672_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _12749_ (.A0(\fifo_bank_register.bank[2][39] ),
    .A1(_05352_),
    .S(_07663_),
    .X(_07673_));
 sky130_fd_sc_hd__clkbuf_1 _12750_ (.A(_07673_),
    .X(_01088_));
 sky130_fd_sc_hd__buf_4 _12751_ (.A(_07651_),
    .X(_07674_));
 sky130_fd_sc_hd__mux2_1 _12752_ (.A0(\fifo_bank_register.bank[2][40] ),
    .A1(_05354_),
    .S(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__clkbuf_1 _12753_ (.A(_07675_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _12754_ (.A0(\fifo_bank_register.bank[2][41] ),
    .A1(_05357_),
    .S(_07674_),
    .X(_07676_));
 sky130_fd_sc_hd__clkbuf_1 _12755_ (.A(_07676_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _12756_ (.A0(\fifo_bank_register.bank[2][42] ),
    .A1(_05359_),
    .S(_07674_),
    .X(_07677_));
 sky130_fd_sc_hd__clkbuf_1 _12757_ (.A(_07677_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _12758_ (.A0(\fifo_bank_register.bank[2][43] ),
    .A1(_05361_),
    .S(_07674_),
    .X(_07678_));
 sky130_fd_sc_hd__clkbuf_1 _12759_ (.A(_07678_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _12760_ (.A0(\fifo_bank_register.bank[2][44] ),
    .A1(_05363_),
    .S(_07674_),
    .X(_07679_));
 sky130_fd_sc_hd__clkbuf_1 _12761_ (.A(_07679_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _12762_ (.A0(\fifo_bank_register.bank[2][45] ),
    .A1(_05365_),
    .S(_07674_),
    .X(_07680_));
 sky130_fd_sc_hd__clkbuf_1 _12763_ (.A(_07680_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _12764_ (.A0(\fifo_bank_register.bank[2][46] ),
    .A1(_05367_),
    .S(_07674_),
    .X(_07681_));
 sky130_fd_sc_hd__clkbuf_1 _12765_ (.A(_07681_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _12766_ (.A0(\fifo_bank_register.bank[2][47] ),
    .A1(_05369_),
    .S(_07674_),
    .X(_07682_));
 sky130_fd_sc_hd__clkbuf_1 _12767_ (.A(_07682_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _12768_ (.A0(\fifo_bank_register.bank[2][48] ),
    .A1(_05371_),
    .S(_07674_),
    .X(_07683_));
 sky130_fd_sc_hd__clkbuf_1 _12769_ (.A(_07683_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _12770_ (.A0(\fifo_bank_register.bank[2][49] ),
    .A1(_05373_),
    .S(_07674_),
    .X(_07684_));
 sky130_fd_sc_hd__clkbuf_1 _12771_ (.A(_07684_),
    .X(_01098_));
 sky130_fd_sc_hd__buf_4 _12772_ (.A(_07651_),
    .X(_07685_));
 sky130_fd_sc_hd__mux2_1 _12773_ (.A0(\fifo_bank_register.bank[2][50] ),
    .A1(_05375_),
    .S(_07685_),
    .X(_07686_));
 sky130_fd_sc_hd__clkbuf_1 _12774_ (.A(_07686_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _12775_ (.A0(\fifo_bank_register.bank[2][51] ),
    .A1(_05378_),
    .S(_07685_),
    .X(_07687_));
 sky130_fd_sc_hd__clkbuf_1 _12776_ (.A(_07687_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _12777_ (.A0(\fifo_bank_register.bank[2][52] ),
    .A1(_05380_),
    .S(_07685_),
    .X(_07688_));
 sky130_fd_sc_hd__clkbuf_1 _12778_ (.A(_07688_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _12779_ (.A0(\fifo_bank_register.bank[2][53] ),
    .A1(_05382_),
    .S(_07685_),
    .X(_07689_));
 sky130_fd_sc_hd__clkbuf_1 _12780_ (.A(_07689_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _12781_ (.A0(\fifo_bank_register.bank[2][54] ),
    .A1(_05384_),
    .S(_07685_),
    .X(_07690_));
 sky130_fd_sc_hd__clkbuf_1 _12782_ (.A(_07690_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _12783_ (.A0(\fifo_bank_register.bank[2][55] ),
    .A1(_05386_),
    .S(_07685_),
    .X(_07691_));
 sky130_fd_sc_hd__clkbuf_1 _12784_ (.A(_07691_),
    .X(_01104_));
 sky130_fd_sc_hd__mux2_1 _12785_ (.A0(\fifo_bank_register.bank[2][56] ),
    .A1(_05388_),
    .S(_07685_),
    .X(_07692_));
 sky130_fd_sc_hd__clkbuf_1 _12786_ (.A(_07692_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _12787_ (.A0(\fifo_bank_register.bank[2][57] ),
    .A1(_05390_),
    .S(_07685_),
    .X(_07693_));
 sky130_fd_sc_hd__clkbuf_1 _12788_ (.A(_07693_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _12789_ (.A0(\fifo_bank_register.bank[2][58] ),
    .A1(_05392_),
    .S(_07685_),
    .X(_07694_));
 sky130_fd_sc_hd__clkbuf_1 _12790_ (.A(_07694_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _12791_ (.A0(\fifo_bank_register.bank[2][59] ),
    .A1(_05394_),
    .S(_07685_),
    .X(_07695_));
 sky130_fd_sc_hd__clkbuf_1 _12792_ (.A(_07695_),
    .X(_01108_));
 sky130_fd_sc_hd__buf_4 _12793_ (.A(_07651_),
    .X(_07696_));
 sky130_fd_sc_hd__mux2_1 _12794_ (.A0(\fifo_bank_register.bank[2][60] ),
    .A1(_05396_),
    .S(_07696_),
    .X(_07697_));
 sky130_fd_sc_hd__clkbuf_1 _12795_ (.A(_07697_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _12796_ (.A0(\fifo_bank_register.bank[2][61] ),
    .A1(_05399_),
    .S(_07696_),
    .X(_07698_));
 sky130_fd_sc_hd__clkbuf_1 _12797_ (.A(_07698_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _12798_ (.A0(\fifo_bank_register.bank[2][62] ),
    .A1(_05401_),
    .S(_07696_),
    .X(_07699_));
 sky130_fd_sc_hd__clkbuf_1 _12799_ (.A(_07699_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _12800_ (.A0(\fifo_bank_register.bank[2][63] ),
    .A1(_05403_),
    .S(_07696_),
    .X(_07700_));
 sky130_fd_sc_hd__clkbuf_1 _12801_ (.A(_07700_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _12802_ (.A0(\fifo_bank_register.bank[2][64] ),
    .A1(_05405_),
    .S(_07696_),
    .X(_07701_));
 sky130_fd_sc_hd__clkbuf_1 _12803_ (.A(_07701_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _12804_ (.A0(\fifo_bank_register.bank[2][65] ),
    .A1(_05407_),
    .S(_07696_),
    .X(_07702_));
 sky130_fd_sc_hd__clkbuf_1 _12805_ (.A(_07702_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _12806_ (.A0(\fifo_bank_register.bank[2][66] ),
    .A1(_05409_),
    .S(_07696_),
    .X(_07703_));
 sky130_fd_sc_hd__clkbuf_1 _12807_ (.A(_07703_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _12808_ (.A0(\fifo_bank_register.bank[2][67] ),
    .A1(_05411_),
    .S(_07696_),
    .X(_07704_));
 sky130_fd_sc_hd__clkbuf_1 _12809_ (.A(_07704_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _12810_ (.A0(\fifo_bank_register.bank[2][68] ),
    .A1(_05413_),
    .S(_07696_),
    .X(_07705_));
 sky130_fd_sc_hd__clkbuf_1 _12811_ (.A(_07705_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _12812_ (.A0(\fifo_bank_register.bank[2][69] ),
    .A1(_05415_),
    .S(_07696_),
    .X(_07706_));
 sky130_fd_sc_hd__clkbuf_1 _12813_ (.A(_07706_),
    .X(_01118_));
 sky130_fd_sc_hd__clkbuf_4 _12814_ (.A(_07651_),
    .X(_07707_));
 sky130_fd_sc_hd__mux2_1 _12815_ (.A0(\fifo_bank_register.bank[2][70] ),
    .A1(_05417_),
    .S(_07707_),
    .X(_07708_));
 sky130_fd_sc_hd__clkbuf_1 _12816_ (.A(_07708_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _12817_ (.A0(\fifo_bank_register.bank[2][71] ),
    .A1(_05420_),
    .S(_07707_),
    .X(_07709_));
 sky130_fd_sc_hd__clkbuf_1 _12818_ (.A(_07709_),
    .X(_01120_));
 sky130_fd_sc_hd__mux2_1 _12819_ (.A0(\fifo_bank_register.bank[2][72] ),
    .A1(_05422_),
    .S(_07707_),
    .X(_07710_));
 sky130_fd_sc_hd__clkbuf_1 _12820_ (.A(_07710_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _12821_ (.A0(\fifo_bank_register.bank[2][73] ),
    .A1(_05424_),
    .S(_07707_),
    .X(_07711_));
 sky130_fd_sc_hd__clkbuf_1 _12822_ (.A(_07711_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _12823_ (.A0(\fifo_bank_register.bank[2][74] ),
    .A1(_05426_),
    .S(_07707_),
    .X(_07712_));
 sky130_fd_sc_hd__clkbuf_1 _12824_ (.A(_07712_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _12825_ (.A0(\fifo_bank_register.bank[2][75] ),
    .A1(_05428_),
    .S(_07707_),
    .X(_07713_));
 sky130_fd_sc_hd__clkbuf_1 _12826_ (.A(_07713_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _12827_ (.A0(\fifo_bank_register.bank[2][76] ),
    .A1(_05430_),
    .S(_07707_),
    .X(_07714_));
 sky130_fd_sc_hd__clkbuf_1 _12828_ (.A(_07714_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _12829_ (.A0(\fifo_bank_register.bank[2][77] ),
    .A1(_05432_),
    .S(_07707_),
    .X(_07715_));
 sky130_fd_sc_hd__clkbuf_1 _12830_ (.A(_07715_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _12831_ (.A0(\fifo_bank_register.bank[2][78] ),
    .A1(_05434_),
    .S(_07707_),
    .X(_07716_));
 sky130_fd_sc_hd__clkbuf_1 _12832_ (.A(_07716_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _12833_ (.A0(\fifo_bank_register.bank[2][79] ),
    .A1(_05436_),
    .S(_07707_),
    .X(_07717_));
 sky130_fd_sc_hd__clkbuf_1 _12834_ (.A(_07717_),
    .X(_01128_));
 sky130_fd_sc_hd__clkbuf_4 _12835_ (.A(_07651_),
    .X(_07718_));
 sky130_fd_sc_hd__mux2_1 _12836_ (.A0(\fifo_bank_register.bank[2][80] ),
    .A1(_05438_),
    .S(_07718_),
    .X(_07719_));
 sky130_fd_sc_hd__clkbuf_1 _12837_ (.A(_07719_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _12838_ (.A0(\fifo_bank_register.bank[2][81] ),
    .A1(_05441_),
    .S(_07718_),
    .X(_07720_));
 sky130_fd_sc_hd__clkbuf_1 _12839_ (.A(_07720_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _12840_ (.A0(\fifo_bank_register.bank[2][82] ),
    .A1(_05443_),
    .S(_07718_),
    .X(_07721_));
 sky130_fd_sc_hd__clkbuf_1 _12841_ (.A(_07721_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _12842_ (.A0(\fifo_bank_register.bank[2][83] ),
    .A1(_05445_),
    .S(_07718_),
    .X(_07722_));
 sky130_fd_sc_hd__clkbuf_1 _12843_ (.A(_07722_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _12844_ (.A0(\fifo_bank_register.bank[2][84] ),
    .A1(_05447_),
    .S(_07718_),
    .X(_07723_));
 sky130_fd_sc_hd__clkbuf_1 _12845_ (.A(_07723_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _12846_ (.A0(\fifo_bank_register.bank[2][85] ),
    .A1(_05449_),
    .S(_07718_),
    .X(_07724_));
 sky130_fd_sc_hd__clkbuf_1 _12847_ (.A(_07724_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _12848_ (.A0(\fifo_bank_register.bank[2][86] ),
    .A1(_05451_),
    .S(_07718_),
    .X(_07725_));
 sky130_fd_sc_hd__clkbuf_1 _12849_ (.A(_07725_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _12850_ (.A0(\fifo_bank_register.bank[2][87] ),
    .A1(_05453_),
    .S(_07718_),
    .X(_07726_));
 sky130_fd_sc_hd__clkbuf_1 _12851_ (.A(_07726_),
    .X(_01136_));
 sky130_fd_sc_hd__mux2_1 _12852_ (.A0(\fifo_bank_register.bank[2][88] ),
    .A1(_05455_),
    .S(_07718_),
    .X(_07727_));
 sky130_fd_sc_hd__clkbuf_1 _12853_ (.A(_07727_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _12854_ (.A0(\fifo_bank_register.bank[2][89] ),
    .A1(_05457_),
    .S(_07718_),
    .X(_07728_));
 sky130_fd_sc_hd__clkbuf_1 _12855_ (.A(_07728_),
    .X(_01138_));
 sky130_fd_sc_hd__buf_4 _12856_ (.A(_07651_),
    .X(_07729_));
 sky130_fd_sc_hd__mux2_1 _12857_ (.A0(\fifo_bank_register.bank[2][90] ),
    .A1(_05459_),
    .S(_07729_),
    .X(_07730_));
 sky130_fd_sc_hd__clkbuf_1 _12858_ (.A(_07730_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _12859_ (.A0(\fifo_bank_register.bank[2][91] ),
    .A1(_05462_),
    .S(_07729_),
    .X(_07731_));
 sky130_fd_sc_hd__clkbuf_1 _12860_ (.A(_07731_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _12861_ (.A0(\fifo_bank_register.bank[2][92] ),
    .A1(_05464_),
    .S(_07729_),
    .X(_07732_));
 sky130_fd_sc_hd__clkbuf_1 _12862_ (.A(_07732_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _12863_ (.A0(\fifo_bank_register.bank[2][93] ),
    .A1(_05466_),
    .S(_07729_),
    .X(_07733_));
 sky130_fd_sc_hd__clkbuf_1 _12864_ (.A(_07733_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _12865_ (.A0(\fifo_bank_register.bank[2][94] ),
    .A1(_05468_),
    .S(_07729_),
    .X(_07734_));
 sky130_fd_sc_hd__clkbuf_1 _12866_ (.A(_07734_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _12867_ (.A0(\fifo_bank_register.bank[2][95] ),
    .A1(_05470_),
    .S(_07729_),
    .X(_07735_));
 sky130_fd_sc_hd__clkbuf_1 _12868_ (.A(_07735_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _12869_ (.A0(\fifo_bank_register.bank[2][96] ),
    .A1(_05472_),
    .S(_07729_),
    .X(_07736_));
 sky130_fd_sc_hd__clkbuf_1 _12870_ (.A(_07736_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _12871_ (.A0(\fifo_bank_register.bank[2][97] ),
    .A1(_05474_),
    .S(_07729_),
    .X(_07737_));
 sky130_fd_sc_hd__clkbuf_1 _12872_ (.A(_07737_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _12873_ (.A0(\fifo_bank_register.bank[2][98] ),
    .A1(_05476_),
    .S(_07729_),
    .X(_07738_));
 sky130_fd_sc_hd__clkbuf_1 _12874_ (.A(_07738_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _12875_ (.A0(\fifo_bank_register.bank[2][99] ),
    .A1(_05478_),
    .S(_07729_),
    .X(_07739_));
 sky130_fd_sc_hd__clkbuf_1 _12876_ (.A(_07739_),
    .X(_01148_));
 sky130_fd_sc_hd__buf_4 _12877_ (.A(_07651_),
    .X(_07740_));
 sky130_fd_sc_hd__mux2_1 _12878_ (.A0(\fifo_bank_register.bank[2][100] ),
    .A1(_05480_),
    .S(_07740_),
    .X(_07741_));
 sky130_fd_sc_hd__clkbuf_1 _12879_ (.A(_07741_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _12880_ (.A0(\fifo_bank_register.bank[2][101] ),
    .A1(_05483_),
    .S(_07740_),
    .X(_07742_));
 sky130_fd_sc_hd__clkbuf_1 _12881_ (.A(_07742_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _12882_ (.A0(\fifo_bank_register.bank[2][102] ),
    .A1(_05485_),
    .S(_07740_),
    .X(_07743_));
 sky130_fd_sc_hd__clkbuf_1 _12883_ (.A(_07743_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _12884_ (.A0(\fifo_bank_register.bank[2][103] ),
    .A1(_05487_),
    .S(_07740_),
    .X(_07744_));
 sky130_fd_sc_hd__clkbuf_1 _12885_ (.A(_07744_),
    .X(_01152_));
 sky130_fd_sc_hd__mux2_1 _12886_ (.A0(\fifo_bank_register.bank[2][104] ),
    .A1(_05489_),
    .S(_07740_),
    .X(_07745_));
 sky130_fd_sc_hd__clkbuf_1 _12887_ (.A(_07745_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _12888_ (.A0(\fifo_bank_register.bank[2][105] ),
    .A1(_05491_),
    .S(_07740_),
    .X(_07746_));
 sky130_fd_sc_hd__clkbuf_1 _12889_ (.A(_07746_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _12890_ (.A0(\fifo_bank_register.bank[2][106] ),
    .A1(_05493_),
    .S(_07740_),
    .X(_07747_));
 sky130_fd_sc_hd__clkbuf_1 _12891_ (.A(_07747_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _12892_ (.A0(\fifo_bank_register.bank[2][107] ),
    .A1(_05495_),
    .S(_07740_),
    .X(_07748_));
 sky130_fd_sc_hd__clkbuf_1 _12893_ (.A(_07748_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _12894_ (.A0(\fifo_bank_register.bank[2][108] ),
    .A1(_05497_),
    .S(_07740_),
    .X(_07749_));
 sky130_fd_sc_hd__clkbuf_1 _12895_ (.A(_07749_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _12896_ (.A0(\fifo_bank_register.bank[2][109] ),
    .A1(_05499_),
    .S(_07740_),
    .X(_07750_));
 sky130_fd_sc_hd__clkbuf_1 _12897_ (.A(_07750_),
    .X(_01158_));
 sky130_fd_sc_hd__clkbuf_4 _12898_ (.A(_07651_),
    .X(_07751_));
 sky130_fd_sc_hd__mux2_1 _12899_ (.A0(\fifo_bank_register.bank[2][110] ),
    .A1(_05501_),
    .S(_07751_),
    .X(_07752_));
 sky130_fd_sc_hd__clkbuf_1 _12900_ (.A(_07752_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _12901_ (.A0(\fifo_bank_register.bank[2][111] ),
    .A1(_05504_),
    .S(_07751_),
    .X(_07753_));
 sky130_fd_sc_hd__clkbuf_1 _12902_ (.A(_07753_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _12903_ (.A0(\fifo_bank_register.bank[2][112] ),
    .A1(_05506_),
    .S(_07751_),
    .X(_07754_));
 sky130_fd_sc_hd__clkbuf_1 _12904_ (.A(_07754_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _12905_ (.A0(\fifo_bank_register.bank[2][113] ),
    .A1(_05508_),
    .S(_07751_),
    .X(_07755_));
 sky130_fd_sc_hd__clkbuf_1 _12906_ (.A(_07755_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _12907_ (.A0(\fifo_bank_register.bank[2][114] ),
    .A1(_05510_),
    .S(_07751_),
    .X(_07756_));
 sky130_fd_sc_hd__clkbuf_1 _12908_ (.A(_07756_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _12909_ (.A0(\fifo_bank_register.bank[2][115] ),
    .A1(_05512_),
    .S(_07751_),
    .X(_07757_));
 sky130_fd_sc_hd__clkbuf_1 _12910_ (.A(_07757_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _12911_ (.A0(\fifo_bank_register.bank[2][116] ),
    .A1(_05514_),
    .S(_07751_),
    .X(_07758_));
 sky130_fd_sc_hd__clkbuf_1 _12912_ (.A(_07758_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _12913_ (.A0(\fifo_bank_register.bank[2][117] ),
    .A1(_05516_),
    .S(_07751_),
    .X(_07759_));
 sky130_fd_sc_hd__clkbuf_1 _12914_ (.A(_07759_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _12915_ (.A0(\fifo_bank_register.bank[2][118] ),
    .A1(_05518_),
    .S(_07751_),
    .X(_07760_));
 sky130_fd_sc_hd__clkbuf_1 _12916_ (.A(_07760_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _12917_ (.A0(\fifo_bank_register.bank[2][119] ),
    .A1(_05520_),
    .S(_07751_),
    .X(_07761_));
 sky130_fd_sc_hd__clkbuf_1 _12918_ (.A(_07761_),
    .X(_01168_));
 sky130_fd_sc_hd__mux2_1 _12919_ (.A0(\fifo_bank_register.bank[2][120] ),
    .A1(_05522_),
    .S(_07628_),
    .X(_07762_));
 sky130_fd_sc_hd__clkbuf_1 _12920_ (.A(_07762_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _12921_ (.A0(\fifo_bank_register.bank[2][121] ),
    .A1(_05524_),
    .S(_07628_),
    .X(_07763_));
 sky130_fd_sc_hd__clkbuf_1 _12922_ (.A(_07763_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _12923_ (.A0(\fifo_bank_register.bank[2][122] ),
    .A1(_05526_),
    .S(_07628_),
    .X(_07764_));
 sky130_fd_sc_hd__clkbuf_1 _12924_ (.A(_07764_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _12925_ (.A0(\fifo_bank_register.bank[2][123] ),
    .A1(_05528_),
    .S(_07628_),
    .X(_07765_));
 sky130_fd_sc_hd__clkbuf_1 _12926_ (.A(_07765_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _12927_ (.A0(\fifo_bank_register.bank[2][124] ),
    .A1(_05530_),
    .S(_07628_),
    .X(_07766_));
 sky130_fd_sc_hd__clkbuf_1 _12928_ (.A(_07766_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _12929_ (.A0(\fifo_bank_register.bank[2][125] ),
    .A1(_05532_),
    .S(_07628_),
    .X(_07767_));
 sky130_fd_sc_hd__clkbuf_1 _12930_ (.A(_07767_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _12931_ (.A0(\fifo_bank_register.bank[2][126] ),
    .A1(_05534_),
    .S(_07628_),
    .X(_07768_));
 sky130_fd_sc_hd__clkbuf_1 _12932_ (.A(_07768_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _12933_ (.A0(\fifo_bank_register.bank[2][127] ),
    .A1(_05536_),
    .S(_07628_),
    .X(_07769_));
 sky130_fd_sc_hd__clkbuf_1 _12934_ (.A(_07769_),
    .X(_01176_));
 sky130_fd_sc_hd__and2_1 _12935_ (.A(_05267_),
    .B(_07483_),
    .X(_07770_));
 sky130_fd_sc_hd__buf_4 _12936_ (.A(_07770_),
    .X(_07771_));
 sky130_fd_sc_hd__buf_4 _12937_ (.A(_07771_),
    .X(_07772_));
 sky130_fd_sc_hd__mux2_1 _12938_ (.A0(\fifo_bank_register.bank[1][0] ),
    .A1(_05248_),
    .S(_07772_),
    .X(_07773_));
 sky130_fd_sc_hd__clkbuf_1 _12939_ (.A(_07773_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _12940_ (.A0(\fifo_bank_register.bank[1][1] ),
    .A1(_05272_),
    .S(_07772_),
    .X(_07774_));
 sky130_fd_sc_hd__clkbuf_1 _12941_ (.A(_07774_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _12942_ (.A0(\fifo_bank_register.bank[1][2] ),
    .A1(_05274_),
    .S(_07772_),
    .X(_07775_));
 sky130_fd_sc_hd__clkbuf_1 _12943_ (.A(_07775_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _12944_ (.A0(\fifo_bank_register.bank[1][3] ),
    .A1(_05276_),
    .S(_07772_),
    .X(_07776_));
 sky130_fd_sc_hd__clkbuf_1 _12945_ (.A(_07776_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _12946_ (.A0(\fifo_bank_register.bank[1][4] ),
    .A1(_05278_),
    .S(_07772_),
    .X(_07777_));
 sky130_fd_sc_hd__clkbuf_1 _12947_ (.A(_07777_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _12948_ (.A0(\fifo_bank_register.bank[1][5] ),
    .A1(_05280_),
    .S(_07772_),
    .X(_07778_));
 sky130_fd_sc_hd__clkbuf_1 _12949_ (.A(_07778_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _12950_ (.A0(\fifo_bank_register.bank[1][6] ),
    .A1(_05282_),
    .S(_07772_),
    .X(_07779_));
 sky130_fd_sc_hd__clkbuf_1 _12951_ (.A(_07779_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _12952_ (.A0(\fifo_bank_register.bank[1][7] ),
    .A1(_05284_),
    .S(_07772_),
    .X(_07780_));
 sky130_fd_sc_hd__clkbuf_1 _12953_ (.A(_07780_),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _12954_ (.A0(\fifo_bank_register.bank[1][8] ),
    .A1(_05286_),
    .S(_07772_),
    .X(_07781_));
 sky130_fd_sc_hd__clkbuf_1 _12955_ (.A(_07781_),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _12956_ (.A0(\fifo_bank_register.bank[1][9] ),
    .A1(_05288_),
    .S(_07772_),
    .X(_07782_));
 sky130_fd_sc_hd__clkbuf_1 _12957_ (.A(_07782_),
    .X(_01186_));
 sky130_fd_sc_hd__buf_4 _12958_ (.A(_07771_),
    .X(_07783_));
 sky130_fd_sc_hd__mux2_1 _12959_ (.A0(\fifo_bank_register.bank[1][10] ),
    .A1(_05290_),
    .S(_07783_),
    .X(_07784_));
 sky130_fd_sc_hd__clkbuf_1 _12960_ (.A(_07784_),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _12961_ (.A0(\fifo_bank_register.bank[1][11] ),
    .A1(_05293_),
    .S(_07783_),
    .X(_07785_));
 sky130_fd_sc_hd__clkbuf_1 _12962_ (.A(_07785_),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _12963_ (.A0(\fifo_bank_register.bank[1][12] ),
    .A1(_05295_),
    .S(_07783_),
    .X(_07786_));
 sky130_fd_sc_hd__clkbuf_1 _12964_ (.A(_07786_),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _12965_ (.A0(\fifo_bank_register.bank[1][13] ),
    .A1(_05297_),
    .S(_07783_),
    .X(_07787_));
 sky130_fd_sc_hd__clkbuf_1 _12966_ (.A(_07787_),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _12967_ (.A0(\fifo_bank_register.bank[1][14] ),
    .A1(_05299_),
    .S(_07783_),
    .X(_07788_));
 sky130_fd_sc_hd__clkbuf_1 _12968_ (.A(_07788_),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _12969_ (.A0(\fifo_bank_register.bank[1][15] ),
    .A1(_05301_),
    .S(_07783_),
    .X(_07789_));
 sky130_fd_sc_hd__clkbuf_1 _12970_ (.A(_07789_),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _12971_ (.A0(\fifo_bank_register.bank[1][16] ),
    .A1(_05303_),
    .S(_07783_),
    .X(_07790_));
 sky130_fd_sc_hd__clkbuf_1 _12972_ (.A(_07790_),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _12973_ (.A0(\fifo_bank_register.bank[1][17] ),
    .A1(_05305_),
    .S(_07783_),
    .X(_07791_));
 sky130_fd_sc_hd__clkbuf_1 _12974_ (.A(_07791_),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _12975_ (.A0(\fifo_bank_register.bank[1][18] ),
    .A1(_05307_),
    .S(_07783_),
    .X(_07792_));
 sky130_fd_sc_hd__clkbuf_1 _12976_ (.A(_07792_),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _12977_ (.A0(\fifo_bank_register.bank[1][19] ),
    .A1(_05309_),
    .S(_07783_),
    .X(_07793_));
 sky130_fd_sc_hd__clkbuf_1 _12978_ (.A(_07793_),
    .X(_01196_));
 sky130_fd_sc_hd__buf_8 _12979_ (.A(_07770_),
    .X(_07794_));
 sky130_fd_sc_hd__buf_4 _12980_ (.A(_07794_),
    .X(_07795_));
 sky130_fd_sc_hd__mux2_1 _12981_ (.A0(\fifo_bank_register.bank[1][20] ),
    .A1(_05311_),
    .S(_07795_),
    .X(_07796_));
 sky130_fd_sc_hd__clkbuf_1 _12982_ (.A(_07796_),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _12983_ (.A0(\fifo_bank_register.bank[1][21] ),
    .A1(_05315_),
    .S(_07795_),
    .X(_07797_));
 sky130_fd_sc_hd__clkbuf_1 _12984_ (.A(_07797_),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _12985_ (.A0(\fifo_bank_register.bank[1][22] ),
    .A1(_05317_),
    .S(_07795_),
    .X(_07798_));
 sky130_fd_sc_hd__clkbuf_1 _12986_ (.A(_07798_),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _12987_ (.A0(\fifo_bank_register.bank[1][23] ),
    .A1(_05319_),
    .S(_07795_),
    .X(_07799_));
 sky130_fd_sc_hd__clkbuf_1 _12988_ (.A(_07799_),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _12989_ (.A0(\fifo_bank_register.bank[1][24] ),
    .A1(_05321_),
    .S(_07795_),
    .X(_07800_));
 sky130_fd_sc_hd__clkbuf_1 _12990_ (.A(_07800_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _12991_ (.A0(\fifo_bank_register.bank[1][25] ),
    .A1(_05323_),
    .S(_07795_),
    .X(_07801_));
 sky130_fd_sc_hd__clkbuf_1 _12992_ (.A(_07801_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _12993_ (.A0(\fifo_bank_register.bank[1][26] ),
    .A1(_05325_),
    .S(_07795_),
    .X(_07802_));
 sky130_fd_sc_hd__clkbuf_1 _12994_ (.A(_07802_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _12995_ (.A0(\fifo_bank_register.bank[1][27] ),
    .A1(_05327_),
    .S(_07795_),
    .X(_07803_));
 sky130_fd_sc_hd__clkbuf_1 _12996_ (.A(_07803_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _12997_ (.A0(\fifo_bank_register.bank[1][28] ),
    .A1(_05329_),
    .S(_07795_),
    .X(_07804_));
 sky130_fd_sc_hd__clkbuf_1 _12998_ (.A(_07804_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _12999_ (.A0(\fifo_bank_register.bank[1][29] ),
    .A1(_05331_),
    .S(_07795_),
    .X(_07805_));
 sky130_fd_sc_hd__clkbuf_1 _13000_ (.A(_07805_),
    .X(_01206_));
 sky130_fd_sc_hd__buf_4 _13001_ (.A(_07794_),
    .X(_07806_));
 sky130_fd_sc_hd__mux2_1 _13002_ (.A0(\fifo_bank_register.bank[1][30] ),
    .A1(_05333_),
    .S(_07806_),
    .X(_07807_));
 sky130_fd_sc_hd__clkbuf_1 _13003_ (.A(_07807_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _13004_ (.A0(\fifo_bank_register.bank[1][31] ),
    .A1(_05336_),
    .S(_07806_),
    .X(_07808_));
 sky130_fd_sc_hd__clkbuf_1 _13005_ (.A(_07808_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _13006_ (.A0(\fifo_bank_register.bank[1][32] ),
    .A1(_05338_),
    .S(_07806_),
    .X(_07809_));
 sky130_fd_sc_hd__clkbuf_1 _13007_ (.A(_07809_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _13008_ (.A0(\fifo_bank_register.bank[1][33] ),
    .A1(_05340_),
    .S(_07806_),
    .X(_07810_));
 sky130_fd_sc_hd__clkbuf_1 _13009_ (.A(_07810_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _13010_ (.A0(\fifo_bank_register.bank[1][34] ),
    .A1(_05342_),
    .S(_07806_),
    .X(_07811_));
 sky130_fd_sc_hd__clkbuf_1 _13011_ (.A(_07811_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _13012_ (.A0(\fifo_bank_register.bank[1][35] ),
    .A1(_05344_),
    .S(_07806_),
    .X(_07812_));
 sky130_fd_sc_hd__clkbuf_1 _13013_ (.A(_07812_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _13014_ (.A0(\fifo_bank_register.bank[1][36] ),
    .A1(_05346_),
    .S(_07806_),
    .X(_07813_));
 sky130_fd_sc_hd__clkbuf_1 _13015_ (.A(_07813_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _13016_ (.A0(\fifo_bank_register.bank[1][37] ),
    .A1(_05348_),
    .S(_07806_),
    .X(_07814_));
 sky130_fd_sc_hd__clkbuf_1 _13017_ (.A(_07814_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _13018_ (.A0(\fifo_bank_register.bank[1][38] ),
    .A1(_05350_),
    .S(_07806_),
    .X(_07815_));
 sky130_fd_sc_hd__clkbuf_1 _13019_ (.A(_07815_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _13020_ (.A0(\fifo_bank_register.bank[1][39] ),
    .A1(_05352_),
    .S(_07806_),
    .X(_07816_));
 sky130_fd_sc_hd__clkbuf_1 _13021_ (.A(_07816_),
    .X(_01216_));
 sky130_fd_sc_hd__buf_4 _13022_ (.A(_07794_),
    .X(_07817_));
 sky130_fd_sc_hd__mux2_1 _13023_ (.A0(\fifo_bank_register.bank[1][40] ),
    .A1(_05354_),
    .S(_07817_),
    .X(_07818_));
 sky130_fd_sc_hd__clkbuf_1 _13024_ (.A(_07818_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _13025_ (.A0(\fifo_bank_register.bank[1][41] ),
    .A1(_05357_),
    .S(_07817_),
    .X(_07819_));
 sky130_fd_sc_hd__clkbuf_1 _13026_ (.A(_07819_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _13027_ (.A0(\fifo_bank_register.bank[1][42] ),
    .A1(_05359_),
    .S(_07817_),
    .X(_07820_));
 sky130_fd_sc_hd__clkbuf_1 _13028_ (.A(_07820_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _13029_ (.A0(\fifo_bank_register.bank[1][43] ),
    .A1(_05361_),
    .S(_07817_),
    .X(_07821_));
 sky130_fd_sc_hd__clkbuf_1 _13030_ (.A(_07821_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _13031_ (.A0(\fifo_bank_register.bank[1][44] ),
    .A1(_05363_),
    .S(_07817_),
    .X(_07822_));
 sky130_fd_sc_hd__clkbuf_1 _13032_ (.A(_07822_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _13033_ (.A0(\fifo_bank_register.bank[1][45] ),
    .A1(_05365_),
    .S(_07817_),
    .X(_07823_));
 sky130_fd_sc_hd__clkbuf_1 _13034_ (.A(_07823_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _13035_ (.A0(\fifo_bank_register.bank[1][46] ),
    .A1(_05367_),
    .S(_07817_),
    .X(_07824_));
 sky130_fd_sc_hd__clkbuf_1 _13036_ (.A(_07824_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _13037_ (.A0(\fifo_bank_register.bank[1][47] ),
    .A1(_05369_),
    .S(_07817_),
    .X(_07825_));
 sky130_fd_sc_hd__clkbuf_1 _13038_ (.A(_07825_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _13039_ (.A0(\fifo_bank_register.bank[1][48] ),
    .A1(_05371_),
    .S(_07817_),
    .X(_07826_));
 sky130_fd_sc_hd__clkbuf_1 _13040_ (.A(_07826_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _13041_ (.A0(\fifo_bank_register.bank[1][49] ),
    .A1(_05373_),
    .S(_07817_),
    .X(_07827_));
 sky130_fd_sc_hd__clkbuf_1 _13042_ (.A(_07827_),
    .X(_01226_));
 sky130_fd_sc_hd__buf_4 _13043_ (.A(_07794_),
    .X(_07828_));
 sky130_fd_sc_hd__mux2_1 _13044_ (.A0(\fifo_bank_register.bank[1][50] ),
    .A1(_05375_),
    .S(_07828_),
    .X(_07829_));
 sky130_fd_sc_hd__clkbuf_1 _13045_ (.A(_07829_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _13046_ (.A0(\fifo_bank_register.bank[1][51] ),
    .A1(_05378_),
    .S(_07828_),
    .X(_07830_));
 sky130_fd_sc_hd__clkbuf_1 _13047_ (.A(_07830_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _13048_ (.A0(\fifo_bank_register.bank[1][52] ),
    .A1(_05380_),
    .S(_07828_),
    .X(_07831_));
 sky130_fd_sc_hd__clkbuf_1 _13049_ (.A(_07831_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _13050_ (.A0(\fifo_bank_register.bank[1][53] ),
    .A1(_05382_),
    .S(_07828_),
    .X(_07832_));
 sky130_fd_sc_hd__clkbuf_1 _13051_ (.A(_07832_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _13052_ (.A0(\fifo_bank_register.bank[1][54] ),
    .A1(_05384_),
    .S(_07828_),
    .X(_07833_));
 sky130_fd_sc_hd__clkbuf_1 _13053_ (.A(_07833_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _13054_ (.A0(\fifo_bank_register.bank[1][55] ),
    .A1(_05386_),
    .S(_07828_),
    .X(_07834_));
 sky130_fd_sc_hd__clkbuf_1 _13055_ (.A(_07834_),
    .X(_01232_));
 sky130_fd_sc_hd__mux2_1 _13056_ (.A0(\fifo_bank_register.bank[1][56] ),
    .A1(_05388_),
    .S(_07828_),
    .X(_07835_));
 sky130_fd_sc_hd__clkbuf_1 _13057_ (.A(_07835_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _13058_ (.A0(\fifo_bank_register.bank[1][57] ),
    .A1(_05390_),
    .S(_07828_),
    .X(_07836_));
 sky130_fd_sc_hd__clkbuf_1 _13059_ (.A(_07836_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _13060_ (.A0(\fifo_bank_register.bank[1][58] ),
    .A1(_05392_),
    .S(_07828_),
    .X(_07837_));
 sky130_fd_sc_hd__clkbuf_1 _13061_ (.A(_07837_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _13062_ (.A0(\fifo_bank_register.bank[1][59] ),
    .A1(_05394_),
    .S(_07828_),
    .X(_07838_));
 sky130_fd_sc_hd__clkbuf_1 _13063_ (.A(_07838_),
    .X(_01236_));
 sky130_fd_sc_hd__buf_4 _13064_ (.A(_07794_),
    .X(_07839_));
 sky130_fd_sc_hd__mux2_1 _13065_ (.A0(\fifo_bank_register.bank[1][60] ),
    .A1(_05396_),
    .S(_07839_),
    .X(_07840_));
 sky130_fd_sc_hd__clkbuf_1 _13066_ (.A(_07840_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _13067_ (.A0(\fifo_bank_register.bank[1][61] ),
    .A1(_05399_),
    .S(_07839_),
    .X(_07841_));
 sky130_fd_sc_hd__clkbuf_1 _13068_ (.A(_07841_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _13069_ (.A0(\fifo_bank_register.bank[1][62] ),
    .A1(_05401_),
    .S(_07839_),
    .X(_07842_));
 sky130_fd_sc_hd__clkbuf_1 _13070_ (.A(_07842_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _13071_ (.A0(\fifo_bank_register.bank[1][63] ),
    .A1(_05403_),
    .S(_07839_),
    .X(_07843_));
 sky130_fd_sc_hd__clkbuf_1 _13072_ (.A(_07843_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _13073_ (.A0(\fifo_bank_register.bank[1][64] ),
    .A1(_05405_),
    .S(_07839_),
    .X(_07844_));
 sky130_fd_sc_hd__clkbuf_1 _13074_ (.A(_07844_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _13075_ (.A0(\fifo_bank_register.bank[1][65] ),
    .A1(_05407_),
    .S(_07839_),
    .X(_07845_));
 sky130_fd_sc_hd__clkbuf_1 _13076_ (.A(_07845_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _13077_ (.A0(\fifo_bank_register.bank[1][66] ),
    .A1(_05409_),
    .S(_07839_),
    .X(_07846_));
 sky130_fd_sc_hd__clkbuf_1 _13078_ (.A(_07846_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _13079_ (.A0(\fifo_bank_register.bank[1][67] ),
    .A1(_05411_),
    .S(_07839_),
    .X(_07847_));
 sky130_fd_sc_hd__clkbuf_1 _13080_ (.A(_07847_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _13081_ (.A0(\fifo_bank_register.bank[1][68] ),
    .A1(_05413_),
    .S(_07839_),
    .X(_07848_));
 sky130_fd_sc_hd__clkbuf_1 _13082_ (.A(_07848_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _13083_ (.A0(\fifo_bank_register.bank[1][69] ),
    .A1(_05415_),
    .S(_07839_),
    .X(_07849_));
 sky130_fd_sc_hd__clkbuf_1 _13084_ (.A(_07849_),
    .X(_01246_));
 sky130_fd_sc_hd__buf_4 _13085_ (.A(_07794_),
    .X(_07850_));
 sky130_fd_sc_hd__mux2_1 _13086_ (.A0(\fifo_bank_register.bank[1][70] ),
    .A1(_05417_),
    .S(_07850_),
    .X(_07851_));
 sky130_fd_sc_hd__clkbuf_1 _13087_ (.A(_07851_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _13088_ (.A0(\fifo_bank_register.bank[1][71] ),
    .A1(_05420_),
    .S(_07850_),
    .X(_07852_));
 sky130_fd_sc_hd__clkbuf_1 _13089_ (.A(_07852_),
    .X(_01248_));
 sky130_fd_sc_hd__mux2_1 _13090_ (.A0(\fifo_bank_register.bank[1][72] ),
    .A1(_05422_),
    .S(_07850_),
    .X(_07853_));
 sky130_fd_sc_hd__clkbuf_1 _13091_ (.A(_07853_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _13092_ (.A0(\fifo_bank_register.bank[1][73] ),
    .A1(_05424_),
    .S(_07850_),
    .X(_07854_));
 sky130_fd_sc_hd__clkbuf_1 _13093_ (.A(_07854_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _13094_ (.A0(\fifo_bank_register.bank[1][74] ),
    .A1(_05426_),
    .S(_07850_),
    .X(_07855_));
 sky130_fd_sc_hd__clkbuf_1 _13095_ (.A(_07855_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _13096_ (.A0(\fifo_bank_register.bank[1][75] ),
    .A1(_05428_),
    .S(_07850_),
    .X(_07856_));
 sky130_fd_sc_hd__clkbuf_1 _13097_ (.A(_07856_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _13098_ (.A0(\fifo_bank_register.bank[1][76] ),
    .A1(_05430_),
    .S(_07850_),
    .X(_07857_));
 sky130_fd_sc_hd__clkbuf_1 _13099_ (.A(_07857_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _13100_ (.A0(\fifo_bank_register.bank[1][77] ),
    .A1(_05432_),
    .S(_07850_),
    .X(_07858_));
 sky130_fd_sc_hd__clkbuf_1 _13101_ (.A(_07858_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _13102_ (.A0(\fifo_bank_register.bank[1][78] ),
    .A1(_05434_),
    .S(_07850_),
    .X(_07859_));
 sky130_fd_sc_hd__clkbuf_1 _13103_ (.A(_07859_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _13104_ (.A0(\fifo_bank_register.bank[1][79] ),
    .A1(_05436_),
    .S(_07850_),
    .X(_07860_));
 sky130_fd_sc_hd__clkbuf_1 _13105_ (.A(_07860_),
    .X(_01256_));
 sky130_fd_sc_hd__buf_4 _13106_ (.A(_07794_),
    .X(_07861_));
 sky130_fd_sc_hd__mux2_1 _13107_ (.A0(\fifo_bank_register.bank[1][80] ),
    .A1(_05438_),
    .S(_07861_),
    .X(_07862_));
 sky130_fd_sc_hd__clkbuf_1 _13108_ (.A(_07862_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _13109_ (.A0(\fifo_bank_register.bank[1][81] ),
    .A1(_05441_),
    .S(_07861_),
    .X(_07863_));
 sky130_fd_sc_hd__clkbuf_1 _13110_ (.A(_07863_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _13111_ (.A0(\fifo_bank_register.bank[1][82] ),
    .A1(_05443_),
    .S(_07861_),
    .X(_07864_));
 sky130_fd_sc_hd__clkbuf_1 _13112_ (.A(_07864_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _13113_ (.A0(\fifo_bank_register.bank[1][83] ),
    .A1(_05445_),
    .S(_07861_),
    .X(_07865_));
 sky130_fd_sc_hd__clkbuf_1 _13114_ (.A(_07865_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _13115_ (.A0(\fifo_bank_register.bank[1][84] ),
    .A1(_05447_),
    .S(_07861_),
    .X(_07866_));
 sky130_fd_sc_hd__clkbuf_1 _13116_ (.A(_07866_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _13117_ (.A0(\fifo_bank_register.bank[1][85] ),
    .A1(_05449_),
    .S(_07861_),
    .X(_07867_));
 sky130_fd_sc_hd__clkbuf_1 _13118_ (.A(_07867_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _13119_ (.A0(\fifo_bank_register.bank[1][86] ),
    .A1(_05451_),
    .S(_07861_),
    .X(_07868_));
 sky130_fd_sc_hd__clkbuf_1 _13120_ (.A(_07868_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _13121_ (.A0(\fifo_bank_register.bank[1][87] ),
    .A1(_05453_),
    .S(_07861_),
    .X(_07869_));
 sky130_fd_sc_hd__clkbuf_1 _13122_ (.A(_07869_),
    .X(_01264_));
 sky130_fd_sc_hd__mux2_1 _13123_ (.A0(\fifo_bank_register.bank[1][88] ),
    .A1(_05455_),
    .S(_07861_),
    .X(_07870_));
 sky130_fd_sc_hd__clkbuf_1 _13124_ (.A(_07870_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _13125_ (.A0(\fifo_bank_register.bank[1][89] ),
    .A1(_05457_),
    .S(_07861_),
    .X(_07871_));
 sky130_fd_sc_hd__clkbuf_1 _13126_ (.A(_07871_),
    .X(_01266_));
 sky130_fd_sc_hd__buf_4 _13127_ (.A(_07794_),
    .X(_07872_));
 sky130_fd_sc_hd__mux2_1 _13128_ (.A0(\fifo_bank_register.bank[1][90] ),
    .A1(_05459_),
    .S(_07872_),
    .X(_07873_));
 sky130_fd_sc_hd__clkbuf_1 _13129_ (.A(_07873_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _13130_ (.A0(\fifo_bank_register.bank[1][91] ),
    .A1(_05462_),
    .S(_07872_),
    .X(_07874_));
 sky130_fd_sc_hd__clkbuf_1 _13131_ (.A(_07874_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _13132_ (.A0(\fifo_bank_register.bank[1][92] ),
    .A1(_05464_),
    .S(_07872_),
    .X(_07875_));
 sky130_fd_sc_hd__clkbuf_1 _13133_ (.A(_07875_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _13134_ (.A0(\fifo_bank_register.bank[1][93] ),
    .A1(_05466_),
    .S(_07872_),
    .X(_07876_));
 sky130_fd_sc_hd__clkbuf_1 _13135_ (.A(_07876_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _13136_ (.A0(\fifo_bank_register.bank[1][94] ),
    .A1(_05468_),
    .S(_07872_),
    .X(_07877_));
 sky130_fd_sc_hd__clkbuf_1 _13137_ (.A(_07877_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _13138_ (.A0(\fifo_bank_register.bank[1][95] ),
    .A1(_05470_),
    .S(_07872_),
    .X(_07878_));
 sky130_fd_sc_hd__clkbuf_1 _13139_ (.A(_07878_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _13140_ (.A0(\fifo_bank_register.bank[1][96] ),
    .A1(_05472_),
    .S(_07872_),
    .X(_07879_));
 sky130_fd_sc_hd__clkbuf_1 _13141_ (.A(_07879_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _13142_ (.A0(\fifo_bank_register.bank[1][97] ),
    .A1(_05474_),
    .S(_07872_),
    .X(_07880_));
 sky130_fd_sc_hd__clkbuf_1 _13143_ (.A(_07880_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _13144_ (.A0(\fifo_bank_register.bank[1][98] ),
    .A1(_05476_),
    .S(_07872_),
    .X(_07881_));
 sky130_fd_sc_hd__clkbuf_1 _13145_ (.A(_07881_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _13146_ (.A0(\fifo_bank_register.bank[1][99] ),
    .A1(_05478_),
    .S(_07872_),
    .X(_07882_));
 sky130_fd_sc_hd__clkbuf_1 _13147_ (.A(_07882_),
    .X(_01276_));
 sky130_fd_sc_hd__buf_4 _13148_ (.A(_07794_),
    .X(_07883_));
 sky130_fd_sc_hd__mux2_1 _13149_ (.A0(\fifo_bank_register.bank[1][100] ),
    .A1(_05480_),
    .S(_07883_),
    .X(_07884_));
 sky130_fd_sc_hd__clkbuf_1 _13150_ (.A(_07884_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _13151_ (.A0(\fifo_bank_register.bank[1][101] ),
    .A1(_05483_),
    .S(_07883_),
    .X(_07885_));
 sky130_fd_sc_hd__clkbuf_1 _13152_ (.A(_07885_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _13153_ (.A0(\fifo_bank_register.bank[1][102] ),
    .A1(_05485_),
    .S(_07883_),
    .X(_07886_));
 sky130_fd_sc_hd__clkbuf_1 _13154_ (.A(_07886_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _13155_ (.A0(\fifo_bank_register.bank[1][103] ),
    .A1(_05487_),
    .S(_07883_),
    .X(_07887_));
 sky130_fd_sc_hd__clkbuf_1 _13156_ (.A(_07887_),
    .X(_01280_));
 sky130_fd_sc_hd__mux2_1 _13157_ (.A0(\fifo_bank_register.bank[1][104] ),
    .A1(_05489_),
    .S(_07883_),
    .X(_07888_));
 sky130_fd_sc_hd__clkbuf_1 _13158_ (.A(_07888_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _13159_ (.A0(\fifo_bank_register.bank[1][105] ),
    .A1(_05491_),
    .S(_07883_),
    .X(_07889_));
 sky130_fd_sc_hd__clkbuf_1 _13160_ (.A(_07889_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _13161_ (.A0(\fifo_bank_register.bank[1][106] ),
    .A1(_05493_),
    .S(_07883_),
    .X(_07890_));
 sky130_fd_sc_hd__clkbuf_1 _13162_ (.A(_07890_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _13163_ (.A0(\fifo_bank_register.bank[1][107] ),
    .A1(_05495_),
    .S(_07883_),
    .X(_07891_));
 sky130_fd_sc_hd__clkbuf_1 _13164_ (.A(_07891_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _13165_ (.A0(\fifo_bank_register.bank[1][108] ),
    .A1(_05497_),
    .S(_07883_),
    .X(_07892_));
 sky130_fd_sc_hd__clkbuf_1 _13166_ (.A(_07892_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _13167_ (.A0(\fifo_bank_register.bank[1][109] ),
    .A1(_05499_),
    .S(_07883_),
    .X(_07893_));
 sky130_fd_sc_hd__clkbuf_1 _13168_ (.A(_07893_),
    .X(_01286_));
 sky130_fd_sc_hd__buf_4 _13169_ (.A(_07794_),
    .X(_07894_));
 sky130_fd_sc_hd__mux2_1 _13170_ (.A0(\fifo_bank_register.bank[1][110] ),
    .A1(_05501_),
    .S(_07894_),
    .X(_07895_));
 sky130_fd_sc_hd__clkbuf_1 _13171_ (.A(_07895_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _13172_ (.A0(\fifo_bank_register.bank[1][111] ),
    .A1(_05504_),
    .S(_07894_),
    .X(_07896_));
 sky130_fd_sc_hd__clkbuf_1 _13173_ (.A(_07896_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _13174_ (.A0(\fifo_bank_register.bank[1][112] ),
    .A1(_05506_),
    .S(_07894_),
    .X(_07897_));
 sky130_fd_sc_hd__clkbuf_1 _13175_ (.A(_07897_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _13176_ (.A0(\fifo_bank_register.bank[1][113] ),
    .A1(_05508_),
    .S(_07894_),
    .X(_07898_));
 sky130_fd_sc_hd__clkbuf_1 _13177_ (.A(_07898_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _13178_ (.A0(\fifo_bank_register.bank[1][114] ),
    .A1(_05510_),
    .S(_07894_),
    .X(_07899_));
 sky130_fd_sc_hd__clkbuf_1 _13179_ (.A(_07899_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _13180_ (.A0(\fifo_bank_register.bank[1][115] ),
    .A1(_05512_),
    .S(_07894_),
    .X(_07900_));
 sky130_fd_sc_hd__clkbuf_1 _13181_ (.A(_07900_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _13182_ (.A0(\fifo_bank_register.bank[1][116] ),
    .A1(_05514_),
    .S(_07894_),
    .X(_07901_));
 sky130_fd_sc_hd__clkbuf_1 _13183_ (.A(_07901_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _13184_ (.A0(\fifo_bank_register.bank[1][117] ),
    .A1(_05516_),
    .S(_07894_),
    .X(_07902_));
 sky130_fd_sc_hd__clkbuf_1 _13185_ (.A(_07902_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _13186_ (.A0(\fifo_bank_register.bank[1][118] ),
    .A1(_05518_),
    .S(_07894_),
    .X(_07903_));
 sky130_fd_sc_hd__clkbuf_1 _13187_ (.A(_07903_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _13188_ (.A0(\fifo_bank_register.bank[1][119] ),
    .A1(_05520_),
    .S(_07894_),
    .X(_07904_));
 sky130_fd_sc_hd__clkbuf_1 _13189_ (.A(_07904_),
    .X(_01296_));
 sky130_fd_sc_hd__mux2_1 _13190_ (.A0(\fifo_bank_register.bank[1][120] ),
    .A1(_05522_),
    .S(_07771_),
    .X(_07905_));
 sky130_fd_sc_hd__clkbuf_1 _13191_ (.A(_07905_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _13192_ (.A0(\fifo_bank_register.bank[1][121] ),
    .A1(_05524_),
    .S(_07771_),
    .X(_07906_));
 sky130_fd_sc_hd__clkbuf_1 _13193_ (.A(_07906_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _13194_ (.A0(\fifo_bank_register.bank[1][122] ),
    .A1(_05526_),
    .S(_07771_),
    .X(_07907_));
 sky130_fd_sc_hd__clkbuf_1 _13195_ (.A(_07907_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _13196_ (.A0(\fifo_bank_register.bank[1][123] ),
    .A1(_05528_),
    .S(_07771_),
    .X(_07908_));
 sky130_fd_sc_hd__clkbuf_1 _13197_ (.A(_07908_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _13198_ (.A0(\fifo_bank_register.bank[1][124] ),
    .A1(_05530_),
    .S(_07771_),
    .X(_07909_));
 sky130_fd_sc_hd__clkbuf_1 _13199_ (.A(_07909_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _13200_ (.A0(\fifo_bank_register.bank[1][125] ),
    .A1(_05532_),
    .S(_07771_),
    .X(_07910_));
 sky130_fd_sc_hd__clkbuf_1 _13201_ (.A(_07910_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _13202_ (.A0(\fifo_bank_register.bank[1][126] ),
    .A1(_05534_),
    .S(_07771_),
    .X(_07911_));
 sky130_fd_sc_hd__clkbuf_1 _13203_ (.A(_07911_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _13204_ (.A0(\fifo_bank_register.bank[1][127] ),
    .A1(_05536_),
    .S(_07771_),
    .X(_07912_));
 sky130_fd_sc_hd__clkbuf_1 _13205_ (.A(_07912_),
    .X(_01304_));
 sky130_fd_sc_hd__or2b_1 _13206_ (.A(_06766_),
    .B_N(_07483_),
    .X(_07913_));
 sky130_fd_sc_hd__buf_4 _13207_ (.A(_07913_),
    .X(_07914_));
 sky130_fd_sc_hd__clkbuf_4 _13208_ (.A(_07914_),
    .X(_07915_));
 sky130_fd_sc_hd__mux2_1 _13209_ (.A0(_05248_),
    .A1(\fifo_bank_register.bank[0][0] ),
    .S(_07915_),
    .X(_07916_));
 sky130_fd_sc_hd__clkbuf_1 _13210_ (.A(_07916_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _13211_ (.A0(_05272_),
    .A1(\fifo_bank_register.bank[0][1] ),
    .S(_07915_),
    .X(_07917_));
 sky130_fd_sc_hd__clkbuf_1 _13212_ (.A(_07917_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _13213_ (.A0(_05274_),
    .A1(\fifo_bank_register.bank[0][2] ),
    .S(_07915_),
    .X(_07918_));
 sky130_fd_sc_hd__clkbuf_1 _13214_ (.A(_07918_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _13215_ (.A0(_05276_),
    .A1(\fifo_bank_register.bank[0][3] ),
    .S(_07915_),
    .X(_07919_));
 sky130_fd_sc_hd__clkbuf_1 _13216_ (.A(_07919_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(_05278_),
    .A1(\fifo_bank_register.bank[0][4] ),
    .S(_07915_),
    .X(_07920_));
 sky130_fd_sc_hd__clkbuf_1 _13218_ (.A(_07920_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _13219_ (.A0(_05280_),
    .A1(\fifo_bank_register.bank[0][5] ),
    .S(_07915_),
    .X(_07921_));
 sky130_fd_sc_hd__clkbuf_1 _13220_ (.A(_07921_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _13221_ (.A0(_05282_),
    .A1(\fifo_bank_register.bank[0][6] ),
    .S(_07915_),
    .X(_07922_));
 sky130_fd_sc_hd__clkbuf_1 _13222_ (.A(_07922_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _13223_ (.A0(_05284_),
    .A1(\fifo_bank_register.bank[0][7] ),
    .S(_07915_),
    .X(_07923_));
 sky130_fd_sc_hd__clkbuf_1 _13224_ (.A(_07923_),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _13225_ (.A0(_05286_),
    .A1(\fifo_bank_register.bank[0][8] ),
    .S(_07915_),
    .X(_07924_));
 sky130_fd_sc_hd__clkbuf_1 _13226_ (.A(_07924_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _13227_ (.A0(_05288_),
    .A1(\fifo_bank_register.bank[0][9] ),
    .S(_07915_),
    .X(_07925_));
 sky130_fd_sc_hd__clkbuf_1 _13228_ (.A(_07925_),
    .X(_01314_));
 sky130_fd_sc_hd__buf_4 _13229_ (.A(_07914_),
    .X(_07926_));
 sky130_fd_sc_hd__mux2_1 _13230_ (.A0(_05290_),
    .A1(\fifo_bank_register.bank[0][10] ),
    .S(_07926_),
    .X(_07927_));
 sky130_fd_sc_hd__clkbuf_1 _13231_ (.A(_07927_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _13232_ (.A0(_05293_),
    .A1(\fifo_bank_register.bank[0][11] ),
    .S(_07926_),
    .X(_07928_));
 sky130_fd_sc_hd__clkbuf_1 _13233_ (.A(_07928_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _13234_ (.A0(_05295_),
    .A1(\fifo_bank_register.bank[0][12] ),
    .S(_07926_),
    .X(_07929_));
 sky130_fd_sc_hd__clkbuf_1 _13235_ (.A(_07929_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _13236_ (.A0(_05297_),
    .A1(\fifo_bank_register.bank[0][13] ),
    .S(_07926_),
    .X(_07930_));
 sky130_fd_sc_hd__clkbuf_1 _13237_ (.A(_07930_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _13238_ (.A0(_05299_),
    .A1(\fifo_bank_register.bank[0][14] ),
    .S(_07926_),
    .X(_07931_));
 sky130_fd_sc_hd__clkbuf_1 _13239_ (.A(_07931_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _13240_ (.A0(_05301_),
    .A1(\fifo_bank_register.bank[0][15] ),
    .S(_07926_),
    .X(_07932_));
 sky130_fd_sc_hd__clkbuf_1 _13241_ (.A(_07932_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _13242_ (.A0(_05303_),
    .A1(\fifo_bank_register.bank[0][16] ),
    .S(_07926_),
    .X(_07933_));
 sky130_fd_sc_hd__clkbuf_1 _13243_ (.A(_07933_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _13244_ (.A0(_05305_),
    .A1(\fifo_bank_register.bank[0][17] ),
    .S(_07926_),
    .X(_07934_));
 sky130_fd_sc_hd__clkbuf_1 _13245_ (.A(_07934_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _13246_ (.A0(_05307_),
    .A1(\fifo_bank_register.bank[0][18] ),
    .S(_07926_),
    .X(_07935_));
 sky130_fd_sc_hd__clkbuf_1 _13247_ (.A(_07935_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _13248_ (.A0(_05309_),
    .A1(\fifo_bank_register.bank[0][19] ),
    .S(_07926_),
    .X(_07936_));
 sky130_fd_sc_hd__clkbuf_1 _13249_ (.A(_07936_),
    .X(_01324_));
 sky130_fd_sc_hd__clkbuf_8 _13250_ (.A(_07913_),
    .X(_07937_));
 sky130_fd_sc_hd__buf_4 _13251_ (.A(_07937_),
    .X(_07938_));
 sky130_fd_sc_hd__mux2_1 _13252_ (.A0(_05311_),
    .A1(\fifo_bank_register.bank[0][20] ),
    .S(_07938_),
    .X(_07939_));
 sky130_fd_sc_hd__clkbuf_1 _13253_ (.A(_07939_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _13254_ (.A0(_05315_),
    .A1(\fifo_bank_register.bank[0][21] ),
    .S(_07938_),
    .X(_07940_));
 sky130_fd_sc_hd__clkbuf_1 _13255_ (.A(_07940_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _13256_ (.A0(_05317_),
    .A1(\fifo_bank_register.bank[0][22] ),
    .S(_07938_),
    .X(_07941_));
 sky130_fd_sc_hd__clkbuf_1 _13257_ (.A(_07941_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _13258_ (.A0(_05319_),
    .A1(\fifo_bank_register.bank[0][23] ),
    .S(_07938_),
    .X(_07942_));
 sky130_fd_sc_hd__clkbuf_1 _13259_ (.A(_07942_),
    .X(_01328_));
 sky130_fd_sc_hd__mux2_1 _13260_ (.A0(_05321_),
    .A1(\fifo_bank_register.bank[0][24] ),
    .S(_07938_),
    .X(_07943_));
 sky130_fd_sc_hd__clkbuf_1 _13261_ (.A(_07943_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _13262_ (.A0(_05323_),
    .A1(\fifo_bank_register.bank[0][25] ),
    .S(_07938_),
    .X(_07944_));
 sky130_fd_sc_hd__clkbuf_1 _13263_ (.A(_07944_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _13264_ (.A0(_05325_),
    .A1(\fifo_bank_register.bank[0][26] ),
    .S(_07938_),
    .X(_07945_));
 sky130_fd_sc_hd__clkbuf_1 _13265_ (.A(_07945_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _13266_ (.A0(_05327_),
    .A1(\fifo_bank_register.bank[0][27] ),
    .S(_07938_),
    .X(_07946_));
 sky130_fd_sc_hd__clkbuf_1 _13267_ (.A(_07946_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _13268_ (.A0(_05329_),
    .A1(\fifo_bank_register.bank[0][28] ),
    .S(_07938_),
    .X(_07947_));
 sky130_fd_sc_hd__clkbuf_1 _13269_ (.A(_07947_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _13270_ (.A0(_05331_),
    .A1(\fifo_bank_register.bank[0][29] ),
    .S(_07938_),
    .X(_07948_));
 sky130_fd_sc_hd__clkbuf_1 _13271_ (.A(_07948_),
    .X(_01334_));
 sky130_fd_sc_hd__buf_4 _13272_ (.A(_07937_),
    .X(_07949_));
 sky130_fd_sc_hd__mux2_1 _13273_ (.A0(_05333_),
    .A1(\fifo_bank_register.bank[0][30] ),
    .S(_07949_),
    .X(_07950_));
 sky130_fd_sc_hd__clkbuf_1 _13274_ (.A(_07950_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _13275_ (.A0(_05336_),
    .A1(\fifo_bank_register.bank[0][31] ),
    .S(_07949_),
    .X(_07951_));
 sky130_fd_sc_hd__clkbuf_1 _13276_ (.A(_07951_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _13277_ (.A0(_05338_),
    .A1(\fifo_bank_register.bank[0][32] ),
    .S(_07949_),
    .X(_07952_));
 sky130_fd_sc_hd__clkbuf_1 _13278_ (.A(_07952_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _13279_ (.A0(_05340_),
    .A1(\fifo_bank_register.bank[0][33] ),
    .S(_07949_),
    .X(_07953_));
 sky130_fd_sc_hd__clkbuf_1 _13280_ (.A(_07953_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _13281_ (.A0(_05342_),
    .A1(\fifo_bank_register.bank[0][34] ),
    .S(_07949_),
    .X(_07954_));
 sky130_fd_sc_hd__clkbuf_1 _13282_ (.A(_07954_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _13283_ (.A0(_05344_),
    .A1(\fifo_bank_register.bank[0][35] ),
    .S(_07949_),
    .X(_07955_));
 sky130_fd_sc_hd__clkbuf_1 _13284_ (.A(_07955_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _13285_ (.A0(_05346_),
    .A1(\fifo_bank_register.bank[0][36] ),
    .S(_07949_),
    .X(_07956_));
 sky130_fd_sc_hd__clkbuf_1 _13286_ (.A(_07956_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _13287_ (.A0(_05348_),
    .A1(\fifo_bank_register.bank[0][37] ),
    .S(_07949_),
    .X(_07957_));
 sky130_fd_sc_hd__clkbuf_1 _13288_ (.A(_07957_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _13289_ (.A0(_05350_),
    .A1(\fifo_bank_register.bank[0][38] ),
    .S(_07949_),
    .X(_07958_));
 sky130_fd_sc_hd__clkbuf_1 _13290_ (.A(_07958_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _13291_ (.A0(_05352_),
    .A1(\fifo_bank_register.bank[0][39] ),
    .S(_07949_),
    .X(_07959_));
 sky130_fd_sc_hd__clkbuf_1 _13292_ (.A(_07959_),
    .X(_01344_));
 sky130_fd_sc_hd__buf_4 _13293_ (.A(_07937_),
    .X(_07960_));
 sky130_fd_sc_hd__mux2_1 _13294_ (.A0(_05354_),
    .A1(\fifo_bank_register.bank[0][40] ),
    .S(_07960_),
    .X(_07961_));
 sky130_fd_sc_hd__clkbuf_1 _13295_ (.A(_07961_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _13296_ (.A0(_05357_),
    .A1(\fifo_bank_register.bank[0][41] ),
    .S(_07960_),
    .X(_07962_));
 sky130_fd_sc_hd__clkbuf_1 _13297_ (.A(_07962_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _13298_ (.A0(_05359_),
    .A1(\fifo_bank_register.bank[0][42] ),
    .S(_07960_),
    .X(_07963_));
 sky130_fd_sc_hd__clkbuf_1 _13299_ (.A(_07963_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _13300_ (.A0(_05361_),
    .A1(\fifo_bank_register.bank[0][43] ),
    .S(_07960_),
    .X(_07964_));
 sky130_fd_sc_hd__clkbuf_1 _13301_ (.A(_07964_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _13302_ (.A0(_05363_),
    .A1(\fifo_bank_register.bank[0][44] ),
    .S(_07960_),
    .X(_07965_));
 sky130_fd_sc_hd__clkbuf_1 _13303_ (.A(_07965_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _13304_ (.A0(_05365_),
    .A1(\fifo_bank_register.bank[0][45] ),
    .S(_07960_),
    .X(_07966_));
 sky130_fd_sc_hd__clkbuf_1 _13305_ (.A(_07966_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _13306_ (.A0(_05367_),
    .A1(\fifo_bank_register.bank[0][46] ),
    .S(_07960_),
    .X(_07967_));
 sky130_fd_sc_hd__clkbuf_1 _13307_ (.A(_07967_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _13308_ (.A0(_05369_),
    .A1(\fifo_bank_register.bank[0][47] ),
    .S(_07960_),
    .X(_07968_));
 sky130_fd_sc_hd__clkbuf_1 _13309_ (.A(_07968_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _13310_ (.A0(_05371_),
    .A1(\fifo_bank_register.bank[0][48] ),
    .S(_07960_),
    .X(_07969_));
 sky130_fd_sc_hd__clkbuf_1 _13311_ (.A(_07969_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _13312_ (.A0(_05373_),
    .A1(\fifo_bank_register.bank[0][49] ),
    .S(_07960_),
    .X(_07970_));
 sky130_fd_sc_hd__clkbuf_1 _13313_ (.A(_07970_),
    .X(_01354_));
 sky130_fd_sc_hd__buf_4 _13314_ (.A(_07937_),
    .X(_07971_));
 sky130_fd_sc_hd__mux2_1 _13315_ (.A0(_05375_),
    .A1(\fifo_bank_register.bank[0][50] ),
    .S(_07971_),
    .X(_07972_));
 sky130_fd_sc_hd__clkbuf_1 _13316_ (.A(_07972_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _13317_ (.A0(_05378_),
    .A1(\fifo_bank_register.bank[0][51] ),
    .S(_07971_),
    .X(_07973_));
 sky130_fd_sc_hd__clkbuf_1 _13318_ (.A(_07973_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _13319_ (.A0(_05380_),
    .A1(\fifo_bank_register.bank[0][52] ),
    .S(_07971_),
    .X(_07974_));
 sky130_fd_sc_hd__clkbuf_1 _13320_ (.A(_07974_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _13321_ (.A0(_05382_),
    .A1(\fifo_bank_register.bank[0][53] ),
    .S(_07971_),
    .X(_07975_));
 sky130_fd_sc_hd__clkbuf_1 _13322_ (.A(_07975_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _13323_ (.A0(_05384_),
    .A1(\fifo_bank_register.bank[0][54] ),
    .S(_07971_),
    .X(_07976_));
 sky130_fd_sc_hd__clkbuf_1 _13324_ (.A(_07976_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _13325_ (.A0(_05386_),
    .A1(\fifo_bank_register.bank[0][55] ),
    .S(_07971_),
    .X(_07977_));
 sky130_fd_sc_hd__clkbuf_1 _13326_ (.A(_07977_),
    .X(_01360_));
 sky130_fd_sc_hd__mux2_1 _13327_ (.A0(_05388_),
    .A1(\fifo_bank_register.bank[0][56] ),
    .S(_07971_),
    .X(_07978_));
 sky130_fd_sc_hd__clkbuf_1 _13328_ (.A(_07978_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _13329_ (.A0(_05390_),
    .A1(\fifo_bank_register.bank[0][57] ),
    .S(_07971_),
    .X(_07979_));
 sky130_fd_sc_hd__clkbuf_1 _13330_ (.A(_07979_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _13331_ (.A0(_05392_),
    .A1(\fifo_bank_register.bank[0][58] ),
    .S(_07971_),
    .X(_07980_));
 sky130_fd_sc_hd__clkbuf_1 _13332_ (.A(_07980_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _13333_ (.A0(_05394_),
    .A1(\fifo_bank_register.bank[0][59] ),
    .S(_07971_),
    .X(_07981_));
 sky130_fd_sc_hd__clkbuf_1 _13334_ (.A(_07981_),
    .X(_01364_));
 sky130_fd_sc_hd__buf_4 _13335_ (.A(_07937_),
    .X(_07982_));
 sky130_fd_sc_hd__mux2_1 _13336_ (.A0(_05396_),
    .A1(\fifo_bank_register.bank[0][60] ),
    .S(_07982_),
    .X(_07983_));
 sky130_fd_sc_hd__clkbuf_1 _13337_ (.A(_07983_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _13338_ (.A0(_05399_),
    .A1(\fifo_bank_register.bank[0][61] ),
    .S(_07982_),
    .X(_07984_));
 sky130_fd_sc_hd__clkbuf_1 _13339_ (.A(_07984_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _13340_ (.A0(_05401_),
    .A1(\fifo_bank_register.bank[0][62] ),
    .S(_07982_),
    .X(_07985_));
 sky130_fd_sc_hd__clkbuf_1 _13341_ (.A(_07985_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _13342_ (.A0(_05403_),
    .A1(\fifo_bank_register.bank[0][63] ),
    .S(_07982_),
    .X(_07986_));
 sky130_fd_sc_hd__clkbuf_1 _13343_ (.A(_07986_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _13344_ (.A0(_05405_),
    .A1(\fifo_bank_register.bank[0][64] ),
    .S(_07982_),
    .X(_07987_));
 sky130_fd_sc_hd__clkbuf_1 _13345_ (.A(_07987_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _13346_ (.A0(_05407_),
    .A1(\fifo_bank_register.bank[0][65] ),
    .S(_07982_),
    .X(_07988_));
 sky130_fd_sc_hd__clkbuf_1 _13347_ (.A(_07988_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _13348_ (.A0(_05409_),
    .A1(\fifo_bank_register.bank[0][66] ),
    .S(_07982_),
    .X(_07989_));
 sky130_fd_sc_hd__clkbuf_1 _13349_ (.A(_07989_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _13350_ (.A0(_05411_),
    .A1(\fifo_bank_register.bank[0][67] ),
    .S(_07982_),
    .X(_07990_));
 sky130_fd_sc_hd__clkbuf_1 _13351_ (.A(_07990_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _13352_ (.A0(_05413_),
    .A1(\fifo_bank_register.bank[0][68] ),
    .S(_07982_),
    .X(_07991_));
 sky130_fd_sc_hd__clkbuf_1 _13353_ (.A(_07991_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _13354_ (.A0(_05415_),
    .A1(\fifo_bank_register.bank[0][69] ),
    .S(_07982_),
    .X(_07992_));
 sky130_fd_sc_hd__clkbuf_1 _13355_ (.A(_07992_),
    .X(_01374_));
 sky130_fd_sc_hd__buf_4 _13356_ (.A(_07937_),
    .X(_07993_));
 sky130_fd_sc_hd__mux2_1 _13357_ (.A0(_05417_),
    .A1(\fifo_bank_register.bank[0][70] ),
    .S(_07993_),
    .X(_07994_));
 sky130_fd_sc_hd__clkbuf_1 _13358_ (.A(_07994_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _13359_ (.A0(_05420_),
    .A1(\fifo_bank_register.bank[0][71] ),
    .S(_07993_),
    .X(_07995_));
 sky130_fd_sc_hd__clkbuf_1 _13360_ (.A(_07995_),
    .X(_01376_));
 sky130_fd_sc_hd__mux2_1 _13361_ (.A0(_05422_),
    .A1(\fifo_bank_register.bank[0][72] ),
    .S(_07993_),
    .X(_07996_));
 sky130_fd_sc_hd__clkbuf_1 _13362_ (.A(_07996_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _13363_ (.A0(_05424_),
    .A1(\fifo_bank_register.bank[0][73] ),
    .S(_07993_),
    .X(_07997_));
 sky130_fd_sc_hd__clkbuf_1 _13364_ (.A(_07997_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _13365_ (.A0(_05426_),
    .A1(\fifo_bank_register.bank[0][74] ),
    .S(_07993_),
    .X(_07998_));
 sky130_fd_sc_hd__clkbuf_1 _13366_ (.A(_07998_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _13367_ (.A0(_05428_),
    .A1(\fifo_bank_register.bank[0][75] ),
    .S(_07993_),
    .X(_07999_));
 sky130_fd_sc_hd__clkbuf_1 _13368_ (.A(_07999_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _13369_ (.A0(_05430_),
    .A1(\fifo_bank_register.bank[0][76] ),
    .S(_07993_),
    .X(_08000_));
 sky130_fd_sc_hd__clkbuf_1 _13370_ (.A(_08000_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _13371_ (.A0(_05432_),
    .A1(\fifo_bank_register.bank[0][77] ),
    .S(_07993_),
    .X(_08001_));
 sky130_fd_sc_hd__clkbuf_1 _13372_ (.A(_08001_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _13373_ (.A0(_05434_),
    .A1(\fifo_bank_register.bank[0][78] ),
    .S(_07993_),
    .X(_08002_));
 sky130_fd_sc_hd__clkbuf_1 _13374_ (.A(_08002_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _13375_ (.A0(_05436_),
    .A1(\fifo_bank_register.bank[0][79] ),
    .S(_07993_),
    .X(_08003_));
 sky130_fd_sc_hd__clkbuf_1 _13376_ (.A(_08003_),
    .X(_01384_));
 sky130_fd_sc_hd__buf_4 _13377_ (.A(_07937_),
    .X(_08004_));
 sky130_fd_sc_hd__mux2_1 _13378_ (.A0(_05438_),
    .A1(\fifo_bank_register.bank[0][80] ),
    .S(_08004_),
    .X(_08005_));
 sky130_fd_sc_hd__clkbuf_1 _13379_ (.A(_08005_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _13380_ (.A0(_05441_),
    .A1(\fifo_bank_register.bank[0][81] ),
    .S(_08004_),
    .X(_08006_));
 sky130_fd_sc_hd__clkbuf_1 _13381_ (.A(_08006_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _13382_ (.A0(_05443_),
    .A1(\fifo_bank_register.bank[0][82] ),
    .S(_08004_),
    .X(_08007_));
 sky130_fd_sc_hd__clkbuf_1 _13383_ (.A(_08007_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _13384_ (.A0(_05445_),
    .A1(\fifo_bank_register.bank[0][83] ),
    .S(_08004_),
    .X(_08008_));
 sky130_fd_sc_hd__clkbuf_1 _13385_ (.A(_08008_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _13386_ (.A0(_05447_),
    .A1(\fifo_bank_register.bank[0][84] ),
    .S(_08004_),
    .X(_08009_));
 sky130_fd_sc_hd__clkbuf_1 _13387_ (.A(_08009_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _13388_ (.A0(_05449_),
    .A1(\fifo_bank_register.bank[0][85] ),
    .S(_08004_),
    .X(_08010_));
 sky130_fd_sc_hd__clkbuf_1 _13389_ (.A(_08010_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _13390_ (.A0(_05451_),
    .A1(\fifo_bank_register.bank[0][86] ),
    .S(_08004_),
    .X(_08011_));
 sky130_fd_sc_hd__clkbuf_1 _13391_ (.A(_08011_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _13392_ (.A0(_05453_),
    .A1(\fifo_bank_register.bank[0][87] ),
    .S(_08004_),
    .X(_08012_));
 sky130_fd_sc_hd__clkbuf_1 _13393_ (.A(_08012_),
    .X(_01392_));
 sky130_fd_sc_hd__mux2_1 _13394_ (.A0(_05455_),
    .A1(\fifo_bank_register.bank[0][88] ),
    .S(_08004_),
    .X(_08013_));
 sky130_fd_sc_hd__clkbuf_1 _13395_ (.A(_08013_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _13396_ (.A0(_05457_),
    .A1(\fifo_bank_register.bank[0][89] ),
    .S(_08004_),
    .X(_08014_));
 sky130_fd_sc_hd__clkbuf_1 _13397_ (.A(_08014_),
    .X(_01394_));
 sky130_fd_sc_hd__buf_4 _13398_ (.A(_07937_),
    .X(_08015_));
 sky130_fd_sc_hd__mux2_1 _13399_ (.A0(_05459_),
    .A1(\fifo_bank_register.bank[0][90] ),
    .S(_08015_),
    .X(_08016_));
 sky130_fd_sc_hd__clkbuf_1 _13400_ (.A(_08016_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _13401_ (.A0(_05462_),
    .A1(\fifo_bank_register.bank[0][91] ),
    .S(_08015_),
    .X(_08017_));
 sky130_fd_sc_hd__clkbuf_1 _13402_ (.A(_08017_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _13403_ (.A0(_05464_),
    .A1(\fifo_bank_register.bank[0][92] ),
    .S(_08015_),
    .X(_08018_));
 sky130_fd_sc_hd__clkbuf_1 _13404_ (.A(_08018_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _13405_ (.A0(_05466_),
    .A1(\fifo_bank_register.bank[0][93] ),
    .S(_08015_),
    .X(_08019_));
 sky130_fd_sc_hd__clkbuf_1 _13406_ (.A(_08019_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _13407_ (.A0(_05468_),
    .A1(\fifo_bank_register.bank[0][94] ),
    .S(_08015_),
    .X(_08020_));
 sky130_fd_sc_hd__clkbuf_1 _13408_ (.A(_08020_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _13409_ (.A0(_05470_),
    .A1(\fifo_bank_register.bank[0][95] ),
    .S(_08015_),
    .X(_08021_));
 sky130_fd_sc_hd__clkbuf_1 _13410_ (.A(_08021_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _13411_ (.A0(_05472_),
    .A1(\fifo_bank_register.bank[0][96] ),
    .S(_08015_),
    .X(_08022_));
 sky130_fd_sc_hd__clkbuf_1 _13412_ (.A(_08022_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _13413_ (.A0(_05474_),
    .A1(\fifo_bank_register.bank[0][97] ),
    .S(_08015_),
    .X(_08023_));
 sky130_fd_sc_hd__clkbuf_1 _13414_ (.A(_08023_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _13415_ (.A0(_05476_),
    .A1(\fifo_bank_register.bank[0][98] ),
    .S(_08015_),
    .X(_08024_));
 sky130_fd_sc_hd__clkbuf_1 _13416_ (.A(_08024_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _13417_ (.A0(_05478_),
    .A1(\fifo_bank_register.bank[0][99] ),
    .S(_08015_),
    .X(_08025_));
 sky130_fd_sc_hd__clkbuf_1 _13418_ (.A(_08025_),
    .X(_01404_));
 sky130_fd_sc_hd__buf_4 _13419_ (.A(_07937_),
    .X(_08026_));
 sky130_fd_sc_hd__mux2_1 _13420_ (.A0(_05480_),
    .A1(\fifo_bank_register.bank[0][100] ),
    .S(_08026_),
    .X(_08027_));
 sky130_fd_sc_hd__clkbuf_1 _13421_ (.A(_08027_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _13422_ (.A0(_05483_),
    .A1(\fifo_bank_register.bank[0][101] ),
    .S(_08026_),
    .X(_08028_));
 sky130_fd_sc_hd__clkbuf_1 _13423_ (.A(_08028_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _13424_ (.A0(_05485_),
    .A1(\fifo_bank_register.bank[0][102] ),
    .S(_08026_),
    .X(_08029_));
 sky130_fd_sc_hd__clkbuf_1 _13425_ (.A(_08029_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _13426_ (.A0(_05487_),
    .A1(\fifo_bank_register.bank[0][103] ),
    .S(_08026_),
    .X(_08030_));
 sky130_fd_sc_hd__clkbuf_1 _13427_ (.A(_08030_),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _13428_ (.A0(_05489_),
    .A1(\fifo_bank_register.bank[0][104] ),
    .S(_08026_),
    .X(_08031_));
 sky130_fd_sc_hd__clkbuf_1 _13429_ (.A(_08031_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _13430_ (.A0(_05491_),
    .A1(\fifo_bank_register.bank[0][105] ),
    .S(_08026_),
    .X(_08032_));
 sky130_fd_sc_hd__clkbuf_1 _13431_ (.A(_08032_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _13432_ (.A0(_05493_),
    .A1(\fifo_bank_register.bank[0][106] ),
    .S(_08026_),
    .X(_08033_));
 sky130_fd_sc_hd__clkbuf_1 _13433_ (.A(_08033_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _13434_ (.A0(_05495_),
    .A1(\fifo_bank_register.bank[0][107] ),
    .S(_08026_),
    .X(_08034_));
 sky130_fd_sc_hd__clkbuf_1 _13435_ (.A(_08034_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _13436_ (.A0(_05497_),
    .A1(\fifo_bank_register.bank[0][108] ),
    .S(_08026_),
    .X(_08035_));
 sky130_fd_sc_hd__clkbuf_1 _13437_ (.A(_08035_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _13438_ (.A0(_05499_),
    .A1(\fifo_bank_register.bank[0][109] ),
    .S(_08026_),
    .X(_08036_));
 sky130_fd_sc_hd__clkbuf_1 _13439_ (.A(_08036_),
    .X(_01414_));
 sky130_fd_sc_hd__buf_4 _13440_ (.A(_07937_),
    .X(_08037_));
 sky130_fd_sc_hd__mux2_1 _13441_ (.A0(_05501_),
    .A1(\fifo_bank_register.bank[0][110] ),
    .S(_08037_),
    .X(_08038_));
 sky130_fd_sc_hd__clkbuf_1 _13442_ (.A(_08038_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _13443_ (.A0(_05504_),
    .A1(\fifo_bank_register.bank[0][111] ),
    .S(_08037_),
    .X(_08039_));
 sky130_fd_sc_hd__clkbuf_1 _13444_ (.A(_08039_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _13445_ (.A0(_05506_),
    .A1(\fifo_bank_register.bank[0][112] ),
    .S(_08037_),
    .X(_08040_));
 sky130_fd_sc_hd__clkbuf_1 _13446_ (.A(_08040_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _13447_ (.A0(_05508_),
    .A1(\fifo_bank_register.bank[0][113] ),
    .S(_08037_),
    .X(_08041_));
 sky130_fd_sc_hd__clkbuf_1 _13448_ (.A(_08041_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _13449_ (.A0(_05510_),
    .A1(\fifo_bank_register.bank[0][114] ),
    .S(_08037_),
    .X(_08042_));
 sky130_fd_sc_hd__clkbuf_1 _13450_ (.A(_08042_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _13451_ (.A0(_05512_),
    .A1(\fifo_bank_register.bank[0][115] ),
    .S(_08037_),
    .X(_08043_));
 sky130_fd_sc_hd__clkbuf_1 _13452_ (.A(_08043_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _13453_ (.A0(_05514_),
    .A1(\fifo_bank_register.bank[0][116] ),
    .S(_08037_),
    .X(_08044_));
 sky130_fd_sc_hd__clkbuf_1 _13454_ (.A(_08044_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _13455_ (.A0(_05516_),
    .A1(\fifo_bank_register.bank[0][117] ),
    .S(_08037_),
    .X(_08045_));
 sky130_fd_sc_hd__clkbuf_1 _13456_ (.A(_08045_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _13457_ (.A0(_05518_),
    .A1(\fifo_bank_register.bank[0][118] ),
    .S(_08037_),
    .X(_08046_));
 sky130_fd_sc_hd__clkbuf_1 _13458_ (.A(_08046_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _13459_ (.A0(_05520_),
    .A1(\fifo_bank_register.bank[0][119] ),
    .S(_08037_),
    .X(_08047_));
 sky130_fd_sc_hd__clkbuf_1 _13460_ (.A(_08047_),
    .X(_01424_));
 sky130_fd_sc_hd__mux2_1 _13461_ (.A0(_05522_),
    .A1(\fifo_bank_register.bank[0][120] ),
    .S(_07914_),
    .X(_08048_));
 sky130_fd_sc_hd__clkbuf_1 _13462_ (.A(_08048_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _13463_ (.A0(_05524_),
    .A1(\fifo_bank_register.bank[0][121] ),
    .S(_07914_),
    .X(_08049_));
 sky130_fd_sc_hd__clkbuf_1 _13464_ (.A(_08049_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _13465_ (.A0(_05526_),
    .A1(\fifo_bank_register.bank[0][122] ),
    .S(_07914_),
    .X(_08050_));
 sky130_fd_sc_hd__clkbuf_1 _13466_ (.A(_08050_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _13467_ (.A0(_05528_),
    .A1(\fifo_bank_register.bank[0][123] ),
    .S(_07914_),
    .X(_08051_));
 sky130_fd_sc_hd__clkbuf_1 _13468_ (.A(_08051_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _13469_ (.A0(_05530_),
    .A1(\fifo_bank_register.bank[0][124] ),
    .S(_07914_),
    .X(_08052_));
 sky130_fd_sc_hd__clkbuf_1 _13470_ (.A(_08052_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _13471_ (.A0(_05532_),
    .A1(\fifo_bank_register.bank[0][125] ),
    .S(_07914_),
    .X(_08053_));
 sky130_fd_sc_hd__clkbuf_1 _13472_ (.A(_08053_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _13473_ (.A0(_05534_),
    .A1(\fifo_bank_register.bank[0][126] ),
    .S(_07914_),
    .X(_08054_));
 sky130_fd_sc_hd__clkbuf_1 _13474_ (.A(_08054_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _13475_ (.A0(_05536_),
    .A1(\fifo_bank_register.bank[0][127] ),
    .S(_07914_),
    .X(_08055_));
 sky130_fd_sc_hd__clkbuf_1 _13476_ (.A(_08055_),
    .X(_01432_));
 sky130_fd_sc_hd__buf_2 _13477_ (.A(\fifo_bank_register.read_ptr[3] ),
    .X(_08056_));
 sky130_fd_sc_hd__or2_1 _13478_ (.A(_08056_),
    .B(\fifo_bank_register.write_ptr[3] ),
    .X(_08057_));
 sky130_fd_sc_hd__nand2_1 _13479_ (.A(_08056_),
    .B(\fifo_bank_register.write_ptr[3] ),
    .Y(_08058_));
 sky130_fd_sc_hd__or2_1 _13480_ (.A(_05262_),
    .B(\fifo_bank_register.write_ptr[2] ),
    .X(_08059_));
 sky130_fd_sc_hd__nand2_1 _13481_ (.A(_05262_),
    .B(\fifo_bank_register.write_ptr[2] ),
    .Y(_08060_));
 sky130_fd_sc_hd__xor2_1 _13482_ (.A(\fifo_bank_register.read_ptr[1] ),
    .B(_05250_),
    .X(_08061_));
 sky130_fd_sc_hd__a221o_1 _13483_ (.A1(_08057_),
    .A2(_08058_),
    .B1(_08059_),
    .B2(_08060_),
    .C1(_08061_),
    .X(_08062_));
 sky130_fd_sc_hd__o21ai_4 _13484_ (.A1(_05258_),
    .A2(_08062_),
    .B1(_04466_),
    .Y(_08063_));
 sky130_fd_sc_hd__buf_4 _13485_ (.A(_08063_),
    .X(_08064_));
 sky130_fd_sc_hd__xnor2_1 _13486_ (.A(\fifo_bank_register.read_ptr[0] ),
    .B(_08064_),
    .Y(_01433_));
 sky130_fd_sc_hd__or2b_1 _13487_ (.A(\fifo_bank_register.read_ptr[1] ),
    .B_N(\fifo_bank_register.read_ptr[0] ),
    .X(_08065_));
 sky130_fd_sc_hd__or2b_1 _13488_ (.A(\fifo_bank_register.read_ptr[0] ),
    .B_N(\fifo_bank_register.read_ptr[1] ),
    .X(_08066_));
 sky130_fd_sc_hd__nand2_1 _13489_ (.A(_08065_),
    .B(_08066_),
    .Y(_08067_));
 sky130_fd_sc_hd__clkbuf_8 _13490_ (.A(_08063_),
    .X(_08068_));
 sky130_fd_sc_hd__or2_1 _13491_ (.A(\fifo_bank_register.read_ptr[0] ),
    .B(\fifo_bank_register.read_ptr[1] ),
    .X(_08069_));
 sky130_fd_sc_hd__nor2_1 _13492_ (.A(_05262_),
    .B(_08069_),
    .Y(_08070_));
 sky130_fd_sc_hd__inv_2 _13493_ (.A(_08063_),
    .Y(_08071_));
 sky130_fd_sc_hd__and3b_1 _13494_ (.A_N(_08070_),
    .B(_08071_),
    .C(_08056_),
    .X(_08072_));
 sky130_fd_sc_hd__a21oi_1 _13495_ (.A1(\fifo_bank_register.read_ptr[0] ),
    .A2(_08068_),
    .B1(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__xnor2_1 _13496_ (.A(_08067_),
    .B(_08073_),
    .Y(_01434_));
 sky130_fd_sc_hd__and3_1 _13497_ (.A(\fifo_bank_register.read_ptr[0] ),
    .B(\fifo_bank_register.read_ptr[1] ),
    .C(_05262_),
    .X(_08074_));
 sky130_fd_sc_hd__nor2_1 _13498_ (.A(_08067_),
    .B(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__nor2b_1 _13499_ (.A(\fifo_bank_register.read_ptr[3] ),
    .B_N(_08074_),
    .Y(_08076_));
 sky130_fd_sc_hd__clkbuf_4 _13500_ (.A(_08076_),
    .X(_08077_));
 sky130_fd_sc_hd__clkbuf_4 _13501_ (.A(_08077_),
    .X(_08078_));
 sky130_fd_sc_hd__a21oi_1 _13502_ (.A1(\fifo_bank_register.read_ptr[0] ),
    .A2(\fifo_bank_register.read_ptr[1] ),
    .B1(_05262_),
    .Y(_08079_));
 sky130_fd_sc_hd__a2111o_1 _13503_ (.A1(_08056_),
    .A2(_08075_),
    .B1(_08078_),
    .C1(_08079_),
    .D1(_08064_),
    .X(_08080_));
 sky130_fd_sc_hd__a21bo_1 _13504_ (.A1(_05262_),
    .A2(_08064_),
    .B1_N(_08080_),
    .X(_01435_));
 sky130_fd_sc_hd__a21oi_1 _13505_ (.A1(_08071_),
    .A2(_08074_),
    .B1(_08056_),
    .Y(_08081_));
 sky130_fd_sc_hd__nor2_1 _13506_ (.A(_08072_),
    .B(_08081_),
    .Y(_01436_));
 sky130_fd_sc_hd__xor2_1 _13507_ (.A(_05249_),
    .B(_05266_),
    .X(_01437_));
 sky130_fd_sc_hd__inv_2 _13508_ (.A(_05260_),
    .Y(_08082_));
 sky130_fd_sc_hd__mux2_1 _13509_ (.A0(_05250_),
    .A1(_08082_),
    .S(_05266_),
    .X(_08083_));
 sky130_fd_sc_hd__clkbuf_1 _13510_ (.A(_08083_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _13511_ (.A0(\fifo_bank_register.write_ptr[2] ),
    .A1(_05264_),
    .S(_05266_),
    .X(_08084_));
 sky130_fd_sc_hd__clkbuf_1 _13512_ (.A(_08084_),
    .X(_01439_));
 sky130_fd_sc_hd__inv_2 _13513_ (.A(_05256_),
    .Y(_08085_));
 sky130_fd_sc_hd__mux2_1 _13514_ (.A0(\fifo_bank_register.write_ptr[3] ),
    .A1(_08085_),
    .S(_05266_),
    .X(_08086_));
 sky130_fd_sc_hd__clkbuf_1 _13515_ (.A(_08086_),
    .X(_01440_));
 sky130_fd_sc_hd__nor2_1 _13516_ (.A(_05262_),
    .B(_08065_),
    .Y(_08087_));
 sky130_fd_sc_hd__and2_1 _13517_ (.A(_08056_),
    .B(_08087_),
    .X(_08088_));
 sky130_fd_sc_hd__clkbuf_4 _13518_ (.A(_08088_),
    .X(_08089_));
 sky130_fd_sc_hd__buf_2 _13519_ (.A(_08089_),
    .X(_08090_));
 sky130_fd_sc_hd__nor3_1 _13520_ (.A(_05262_),
    .B(_08056_),
    .C(_08066_),
    .Y(_08091_));
 sky130_fd_sc_hd__clkbuf_4 _13521_ (.A(_08091_),
    .X(_08092_));
 sky130_fd_sc_hd__clkbuf_4 _13522_ (.A(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__or2b_1 _13523_ (.A(\fifo_bank_register.read_ptr[3] ),
    .B_N(\fifo_bank_register.read_ptr[2] ),
    .X(_08094_));
 sky130_fd_sc_hd__nor2_1 _13524_ (.A(_08065_),
    .B(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__clkbuf_4 _13525_ (.A(_08095_),
    .X(_08096_));
 sky130_fd_sc_hd__clkbuf_4 _13526_ (.A(_08096_),
    .X(_08097_));
 sky130_fd_sc_hd__and4bb_1 _13527_ (.A_N(_05262_),
    .B_N(\fifo_bank_register.read_ptr[3] ),
    .C(\fifo_bank_register.read_ptr[0] ),
    .D(\fifo_bank_register.read_ptr[1] ),
    .X(_08098_));
 sky130_fd_sc_hd__clkbuf_4 _13528_ (.A(_08098_),
    .X(_08099_));
 sky130_fd_sc_hd__clkbuf_4 _13529_ (.A(_08099_),
    .X(_08100_));
 sky130_fd_sc_hd__a22o_1 _13530_ (.A1(\fifo_bank_register.bank[5][0] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][0] ),
    .X(_08101_));
 sky130_fd_sc_hd__a221o_1 _13531_ (.A1(\fifo_bank_register.bank[7][0] ),
    .A2(_08078_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][0] ),
    .C1(_08101_),
    .X(_08102_));
 sky130_fd_sc_hd__nor2_1 _13532_ (.A(_08066_),
    .B(_08094_),
    .Y(_08103_));
 sky130_fd_sc_hd__clkbuf_4 _13533_ (.A(_08103_),
    .X(_08104_));
 sky130_fd_sc_hd__clkbuf_4 _13534_ (.A(_08104_),
    .X(_08105_));
 sky130_fd_sc_hd__nor2_1 _13535_ (.A(_08069_),
    .B(_08094_),
    .Y(_08106_));
 sky130_fd_sc_hd__clkbuf_4 _13536_ (.A(_08106_),
    .X(_08107_));
 sky130_fd_sc_hd__clkbuf_4 _13537_ (.A(_08107_),
    .X(_08108_));
 sky130_fd_sc_hd__a22o_1 _13538_ (.A1(\fifo_bank_register.bank[6][0] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][0] ),
    .X(_08109_));
 sky130_fd_sc_hd__and2b_1 _13539_ (.A_N(_08056_),
    .B(_08087_),
    .X(_08110_));
 sky130_fd_sc_hd__clkbuf_4 _13540_ (.A(_08110_),
    .X(_08111_));
 sky130_fd_sc_hd__buf_2 _13541_ (.A(_08111_),
    .X(_08112_));
 sky130_fd_sc_hd__and2_1 _13542_ (.A(_08056_),
    .B(_08070_),
    .X(_08113_));
 sky130_fd_sc_hd__clkbuf_4 _13543_ (.A(_08113_),
    .X(_08114_));
 sky130_fd_sc_hd__clkbuf_4 _13544_ (.A(_08114_),
    .X(_08115_));
 sky130_fd_sc_hd__a22o_1 _13545_ (.A1(\fifo_bank_register.bank[1][0] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][0] ),
    .X(_08116_));
 sky130_fd_sc_hd__a2111o_1 _13546_ (.A1(\fifo_bank_register.bank[9][0] ),
    .A2(_08090_),
    .B1(_08102_),
    .C1(_08109_),
    .D1(_08116_),
    .X(_08117_));
 sky130_fd_sc_hd__nor2_1 _13547_ (.A(_08056_),
    .B(_08070_),
    .Y(_08118_));
 sky130_fd_sc_hd__or3_1 _13548_ (.A(_08087_),
    .B(_08113_),
    .C(_08118_),
    .X(_08119_));
 sky130_fd_sc_hd__buf_4 _13549_ (.A(_08119_),
    .X(_08120_));
 sky130_fd_sc_hd__clkbuf_4 _13550_ (.A(_08120_),
    .X(_08121_));
 sky130_fd_sc_hd__mux2_1 _13551_ (.A0(\fifo_bank_register.bank[0][0] ),
    .A1(_08117_),
    .S(_08121_),
    .X(_08122_));
 sky130_fd_sc_hd__mux2_1 _13552_ (.A0(_08122_),
    .A1(\fifo_bank_register.data_out[0] ),
    .S(_08064_),
    .X(_08123_));
 sky130_fd_sc_hd__clkbuf_1 _13553_ (.A(_08123_),
    .X(_01441_));
 sky130_fd_sc_hd__a22o_1 _13554_ (.A1(\fifo_bank_register.bank[5][1] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][1] ),
    .X(_08124_));
 sky130_fd_sc_hd__a221o_1 _13555_ (.A1(\fifo_bank_register.bank[7][1] ),
    .A2(_08078_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][1] ),
    .C1(_08124_),
    .X(_08125_));
 sky130_fd_sc_hd__a22o_1 _13556_ (.A1(\fifo_bank_register.bank[6][1] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][1] ),
    .X(_08126_));
 sky130_fd_sc_hd__a22o_1 _13557_ (.A1(\fifo_bank_register.bank[1][1] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][1] ),
    .X(_08127_));
 sky130_fd_sc_hd__a2111o_1 _13558_ (.A1(\fifo_bank_register.bank[9][1] ),
    .A2(_08090_),
    .B1(_08125_),
    .C1(_08126_),
    .D1(_08127_),
    .X(_08128_));
 sky130_fd_sc_hd__mux2_1 _13559_ (.A0(\fifo_bank_register.bank[0][1] ),
    .A1(_08128_),
    .S(_08121_),
    .X(_08129_));
 sky130_fd_sc_hd__mux2_1 _13560_ (.A0(_08129_),
    .A1(\fifo_bank_register.data_out[1] ),
    .S(_08064_),
    .X(_08130_));
 sky130_fd_sc_hd__clkbuf_1 _13561_ (.A(_08130_),
    .X(_01442_));
 sky130_fd_sc_hd__a22o_1 _13562_ (.A1(\fifo_bank_register.bank[5][2] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][2] ),
    .X(_08131_));
 sky130_fd_sc_hd__a221o_1 _13563_ (.A1(\fifo_bank_register.bank[7][2] ),
    .A2(_08078_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][2] ),
    .C1(_08131_),
    .X(_08132_));
 sky130_fd_sc_hd__a22o_1 _13564_ (.A1(\fifo_bank_register.bank[6][2] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][2] ),
    .X(_08133_));
 sky130_fd_sc_hd__a22o_1 _13565_ (.A1(\fifo_bank_register.bank[1][2] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][2] ),
    .X(_08134_));
 sky130_fd_sc_hd__a2111o_1 _13566_ (.A1(\fifo_bank_register.bank[9][2] ),
    .A2(_08090_),
    .B1(_08132_),
    .C1(_08133_),
    .D1(_08134_),
    .X(_08135_));
 sky130_fd_sc_hd__mux2_1 _13567_ (.A0(\fifo_bank_register.bank[0][2] ),
    .A1(_08135_),
    .S(_08121_),
    .X(_08136_));
 sky130_fd_sc_hd__mux2_1 _13568_ (.A0(_08136_),
    .A1(\fifo_bank_register.data_out[2] ),
    .S(_08064_),
    .X(_08137_));
 sky130_fd_sc_hd__clkbuf_1 _13569_ (.A(_08137_),
    .X(_01443_));
 sky130_fd_sc_hd__a22o_1 _13570_ (.A1(\fifo_bank_register.bank[5][3] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][3] ),
    .X(_08138_));
 sky130_fd_sc_hd__a221o_1 _13571_ (.A1(\fifo_bank_register.bank[7][3] ),
    .A2(_08078_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][3] ),
    .C1(_08138_),
    .X(_08139_));
 sky130_fd_sc_hd__a22o_1 _13572_ (.A1(\fifo_bank_register.bank[6][3] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][3] ),
    .X(_08140_));
 sky130_fd_sc_hd__a22o_1 _13573_ (.A1(\fifo_bank_register.bank[1][3] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][3] ),
    .X(_08141_));
 sky130_fd_sc_hd__a2111o_1 _13574_ (.A1(\fifo_bank_register.bank[9][3] ),
    .A2(_08090_),
    .B1(_08139_),
    .C1(_08140_),
    .D1(_08141_),
    .X(_08142_));
 sky130_fd_sc_hd__mux2_1 _13575_ (.A0(\fifo_bank_register.bank[0][3] ),
    .A1(_08142_),
    .S(_08121_),
    .X(_08143_));
 sky130_fd_sc_hd__mux2_1 _13576_ (.A0(_08143_),
    .A1(\fifo_bank_register.data_out[3] ),
    .S(_08064_),
    .X(_08144_));
 sky130_fd_sc_hd__clkbuf_1 _13577_ (.A(_08144_),
    .X(_01444_));
 sky130_fd_sc_hd__a22o_1 _13578_ (.A1(\fifo_bank_register.bank[5][4] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][4] ),
    .X(_08145_));
 sky130_fd_sc_hd__a221o_1 _13579_ (.A1(\fifo_bank_register.bank[7][4] ),
    .A2(_08078_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][4] ),
    .C1(_08145_),
    .X(_08146_));
 sky130_fd_sc_hd__a22o_1 _13580_ (.A1(\fifo_bank_register.bank[6][4] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][4] ),
    .X(_08147_));
 sky130_fd_sc_hd__a22o_1 _13581_ (.A1(\fifo_bank_register.bank[1][4] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][4] ),
    .X(_08148_));
 sky130_fd_sc_hd__a2111o_1 _13582_ (.A1(\fifo_bank_register.bank[9][4] ),
    .A2(_08090_),
    .B1(_08146_),
    .C1(_08147_),
    .D1(_08148_),
    .X(_08149_));
 sky130_fd_sc_hd__mux2_1 _13583_ (.A0(\fifo_bank_register.bank[0][4] ),
    .A1(_08149_),
    .S(_08121_),
    .X(_08150_));
 sky130_fd_sc_hd__mux2_1 _13584_ (.A0(_08150_),
    .A1(\fifo_bank_register.data_out[4] ),
    .S(_08064_),
    .X(_08151_));
 sky130_fd_sc_hd__clkbuf_1 _13585_ (.A(_08151_),
    .X(_01445_));
 sky130_fd_sc_hd__a22o_1 _13586_ (.A1(\fifo_bank_register.bank[5][5] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][5] ),
    .X(_08152_));
 sky130_fd_sc_hd__a221o_1 _13587_ (.A1(\fifo_bank_register.bank[7][5] ),
    .A2(_08078_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][5] ),
    .C1(_08152_),
    .X(_08153_));
 sky130_fd_sc_hd__a22o_1 _13588_ (.A1(\fifo_bank_register.bank[6][5] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][5] ),
    .X(_08154_));
 sky130_fd_sc_hd__a22o_1 _13589_ (.A1(\fifo_bank_register.bank[1][5] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][5] ),
    .X(_08155_));
 sky130_fd_sc_hd__a2111o_1 _13590_ (.A1(\fifo_bank_register.bank[9][5] ),
    .A2(_08090_),
    .B1(_08153_),
    .C1(_08154_),
    .D1(_08155_),
    .X(_08156_));
 sky130_fd_sc_hd__mux2_1 _13591_ (.A0(\fifo_bank_register.bank[0][5] ),
    .A1(_08156_),
    .S(_08121_),
    .X(_08157_));
 sky130_fd_sc_hd__mux2_1 _13592_ (.A0(_08157_),
    .A1(\fifo_bank_register.data_out[5] ),
    .S(_08064_),
    .X(_08158_));
 sky130_fd_sc_hd__clkbuf_1 _13593_ (.A(_08158_),
    .X(_01446_));
 sky130_fd_sc_hd__a22o_1 _13594_ (.A1(\fifo_bank_register.bank[5][6] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][6] ),
    .X(_08159_));
 sky130_fd_sc_hd__a221o_1 _13595_ (.A1(\fifo_bank_register.bank[7][6] ),
    .A2(_08078_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][6] ),
    .C1(_08159_),
    .X(_08160_));
 sky130_fd_sc_hd__a22o_1 _13596_ (.A1(\fifo_bank_register.bank[6][6] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][6] ),
    .X(_08161_));
 sky130_fd_sc_hd__a22o_1 _13597_ (.A1(\fifo_bank_register.bank[1][6] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][6] ),
    .X(_08162_));
 sky130_fd_sc_hd__a2111o_1 _13598_ (.A1(\fifo_bank_register.bank[9][6] ),
    .A2(_08090_),
    .B1(_08160_),
    .C1(_08161_),
    .D1(_08162_),
    .X(_08163_));
 sky130_fd_sc_hd__mux2_1 _13599_ (.A0(\fifo_bank_register.bank[0][6] ),
    .A1(_08163_),
    .S(_08121_),
    .X(_08164_));
 sky130_fd_sc_hd__mux2_1 _13600_ (.A0(_08164_),
    .A1(\fifo_bank_register.data_out[6] ),
    .S(_08064_),
    .X(_08165_));
 sky130_fd_sc_hd__clkbuf_1 _13601_ (.A(_08165_),
    .X(_01447_));
 sky130_fd_sc_hd__a22o_1 _13602_ (.A1(\fifo_bank_register.bank[5][7] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][7] ),
    .X(_08166_));
 sky130_fd_sc_hd__a221o_1 _13603_ (.A1(\fifo_bank_register.bank[7][7] ),
    .A2(_08078_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][7] ),
    .C1(_08166_),
    .X(_08167_));
 sky130_fd_sc_hd__a22o_1 _13604_ (.A1(\fifo_bank_register.bank[6][7] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][7] ),
    .X(_08168_));
 sky130_fd_sc_hd__a22o_1 _13605_ (.A1(\fifo_bank_register.bank[1][7] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][7] ),
    .X(_08169_));
 sky130_fd_sc_hd__a2111o_1 _13606_ (.A1(\fifo_bank_register.bank[9][7] ),
    .A2(_08090_),
    .B1(_08167_),
    .C1(_08168_),
    .D1(_08169_),
    .X(_08170_));
 sky130_fd_sc_hd__mux2_1 _13607_ (.A0(\fifo_bank_register.bank[0][7] ),
    .A1(_08170_),
    .S(_08121_),
    .X(_08171_));
 sky130_fd_sc_hd__clkbuf_8 _13608_ (.A(_08068_),
    .X(_08172_));
 sky130_fd_sc_hd__mux2_1 _13609_ (.A0(_08171_),
    .A1(\fifo_bank_register.data_out[7] ),
    .S(_08172_),
    .X(_08173_));
 sky130_fd_sc_hd__clkbuf_1 _13610_ (.A(_08173_),
    .X(_01448_));
 sky130_fd_sc_hd__a22o_1 _13611_ (.A1(\fifo_bank_register.bank[5][8] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][8] ),
    .X(_08174_));
 sky130_fd_sc_hd__a221o_1 _13612_ (.A1(\fifo_bank_register.bank[7][8] ),
    .A2(_08078_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][8] ),
    .C1(_08174_),
    .X(_08175_));
 sky130_fd_sc_hd__a22o_1 _13613_ (.A1(\fifo_bank_register.bank[6][8] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][8] ),
    .X(_08176_));
 sky130_fd_sc_hd__a22o_1 _13614_ (.A1(\fifo_bank_register.bank[1][8] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][8] ),
    .X(_08177_));
 sky130_fd_sc_hd__a2111o_1 _13615_ (.A1(\fifo_bank_register.bank[9][8] ),
    .A2(_08090_),
    .B1(_08175_),
    .C1(_08176_),
    .D1(_08177_),
    .X(_08178_));
 sky130_fd_sc_hd__mux2_1 _13616_ (.A0(\fifo_bank_register.bank[0][8] ),
    .A1(_08178_),
    .S(_08121_),
    .X(_08179_));
 sky130_fd_sc_hd__mux2_1 _13617_ (.A0(_08179_),
    .A1(\fifo_bank_register.data_out[8] ),
    .S(_08172_),
    .X(_08180_));
 sky130_fd_sc_hd__clkbuf_1 _13618_ (.A(_08180_),
    .X(_01449_));
 sky130_fd_sc_hd__buf_6 _13619_ (.A(_08076_),
    .X(_08181_));
 sky130_fd_sc_hd__buf_4 _13620_ (.A(_08181_),
    .X(_08182_));
 sky130_fd_sc_hd__a22o_1 _13621_ (.A1(\fifo_bank_register.bank[5][9] ),
    .A2(_08097_),
    .B1(_08100_),
    .B2(\fifo_bank_register.bank[3][9] ),
    .X(_08183_));
 sky130_fd_sc_hd__a221o_1 _13622_ (.A1(\fifo_bank_register.bank[7][9] ),
    .A2(_08182_),
    .B1(_08093_),
    .B2(\fifo_bank_register.bank[2][9] ),
    .C1(_08183_),
    .X(_08184_));
 sky130_fd_sc_hd__a22o_1 _13623_ (.A1(\fifo_bank_register.bank[6][9] ),
    .A2(_08105_),
    .B1(_08108_),
    .B2(\fifo_bank_register.bank[4][9] ),
    .X(_08185_));
 sky130_fd_sc_hd__a22o_1 _13624_ (.A1(\fifo_bank_register.bank[1][9] ),
    .A2(_08112_),
    .B1(_08115_),
    .B2(\fifo_bank_register.bank[8][9] ),
    .X(_08186_));
 sky130_fd_sc_hd__a2111o_1 _13625_ (.A1(\fifo_bank_register.bank[9][9] ),
    .A2(_08090_),
    .B1(_08184_),
    .C1(_08185_),
    .D1(_08186_),
    .X(_08187_));
 sky130_fd_sc_hd__mux2_1 _13626_ (.A0(\fifo_bank_register.bank[0][9] ),
    .A1(_08187_),
    .S(_08121_),
    .X(_08188_));
 sky130_fd_sc_hd__mux2_1 _13627_ (.A0(_08188_),
    .A1(\fifo_bank_register.data_out[9] ),
    .S(_08172_),
    .X(_08189_));
 sky130_fd_sc_hd__clkbuf_1 _13628_ (.A(_08189_),
    .X(_01450_));
 sky130_fd_sc_hd__clkbuf_4 _13629_ (.A(_08089_),
    .X(_08190_));
 sky130_fd_sc_hd__clkbuf_4 _13630_ (.A(_08092_),
    .X(_08191_));
 sky130_fd_sc_hd__clkbuf_4 _13631_ (.A(_08096_),
    .X(_08192_));
 sky130_fd_sc_hd__clkbuf_4 _13632_ (.A(_08099_),
    .X(_08193_));
 sky130_fd_sc_hd__a22o_1 _13633_ (.A1(\fifo_bank_register.bank[5][10] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][10] ),
    .X(_08194_));
 sky130_fd_sc_hd__a221o_1 _13634_ (.A1(\fifo_bank_register.bank[7][10] ),
    .A2(_08182_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][10] ),
    .C1(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__clkbuf_4 _13635_ (.A(_08104_),
    .X(_08196_));
 sky130_fd_sc_hd__clkbuf_4 _13636_ (.A(_08107_),
    .X(_08197_));
 sky130_fd_sc_hd__a22o_1 _13637_ (.A1(\fifo_bank_register.bank[6][10] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][10] ),
    .X(_08198_));
 sky130_fd_sc_hd__clkbuf_4 _13638_ (.A(_08111_),
    .X(_08199_));
 sky130_fd_sc_hd__clkbuf_4 _13639_ (.A(_08114_),
    .X(_08200_));
 sky130_fd_sc_hd__a22o_1 _13640_ (.A1(\fifo_bank_register.bank[1][10] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][10] ),
    .X(_08201_));
 sky130_fd_sc_hd__a2111o_1 _13641_ (.A1(\fifo_bank_register.bank[9][10] ),
    .A2(_08190_),
    .B1(_08195_),
    .C1(_08198_),
    .D1(_08201_),
    .X(_02067_));
 sky130_fd_sc_hd__buf_4 _13642_ (.A(_08120_),
    .X(_02068_));
 sky130_fd_sc_hd__mux2_1 _13643_ (.A0(\fifo_bank_register.bank[0][10] ),
    .A1(_02067_),
    .S(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_1 _13644_ (.A0(_02069_),
    .A1(\fifo_bank_register.data_out[10] ),
    .S(_08172_),
    .X(_02070_));
 sky130_fd_sc_hd__clkbuf_1 _13645_ (.A(_02070_),
    .X(_01451_));
 sky130_fd_sc_hd__a22o_1 _13646_ (.A1(\fifo_bank_register.bank[5][11] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][11] ),
    .X(_02071_));
 sky130_fd_sc_hd__a221o_1 _13647_ (.A1(\fifo_bank_register.bank[7][11] ),
    .A2(_08182_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][11] ),
    .C1(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__a22o_1 _13648_ (.A1(\fifo_bank_register.bank[6][11] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][11] ),
    .X(_02073_));
 sky130_fd_sc_hd__a22o_1 _13649_ (.A1(\fifo_bank_register.bank[1][11] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][11] ),
    .X(_02074_));
 sky130_fd_sc_hd__a2111o_1 _13650_ (.A1(\fifo_bank_register.bank[9][11] ),
    .A2(_08190_),
    .B1(_02072_),
    .C1(_02073_),
    .D1(_02074_),
    .X(_02075_));
 sky130_fd_sc_hd__mux2_1 _13651_ (.A0(\fifo_bank_register.bank[0][11] ),
    .A1(_02075_),
    .S(_02068_),
    .X(_02076_));
 sky130_fd_sc_hd__mux2_1 _13652_ (.A0(_02076_),
    .A1(\fifo_bank_register.data_out[11] ),
    .S(_08172_),
    .X(_02077_));
 sky130_fd_sc_hd__clkbuf_1 _13653_ (.A(_02077_),
    .X(_01452_));
 sky130_fd_sc_hd__a22o_1 _13654_ (.A1(\fifo_bank_register.bank[5][12] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][12] ),
    .X(_02078_));
 sky130_fd_sc_hd__a221o_1 _13655_ (.A1(\fifo_bank_register.bank[7][12] ),
    .A2(_08182_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][12] ),
    .C1(_02078_),
    .X(_02079_));
 sky130_fd_sc_hd__a22o_1 _13656_ (.A1(\fifo_bank_register.bank[6][12] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][12] ),
    .X(_02080_));
 sky130_fd_sc_hd__a22o_1 _13657_ (.A1(\fifo_bank_register.bank[1][12] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][12] ),
    .X(_02081_));
 sky130_fd_sc_hd__a2111o_1 _13658_ (.A1(\fifo_bank_register.bank[9][12] ),
    .A2(_08190_),
    .B1(_02079_),
    .C1(_02080_),
    .D1(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__mux2_1 _13659_ (.A0(\fifo_bank_register.bank[0][12] ),
    .A1(_02082_),
    .S(_02068_),
    .X(_02083_));
 sky130_fd_sc_hd__mux2_1 _13660_ (.A0(_02083_),
    .A1(\fifo_bank_register.data_out[12] ),
    .S(_08172_),
    .X(_02084_));
 sky130_fd_sc_hd__clkbuf_1 _13661_ (.A(_02084_),
    .X(_01453_));
 sky130_fd_sc_hd__a22o_1 _13662_ (.A1(\fifo_bank_register.bank[5][13] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][13] ),
    .X(_02085_));
 sky130_fd_sc_hd__a221o_1 _13663_ (.A1(\fifo_bank_register.bank[7][13] ),
    .A2(_08182_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][13] ),
    .C1(_02085_),
    .X(_02086_));
 sky130_fd_sc_hd__a22o_1 _13664_ (.A1(\fifo_bank_register.bank[6][13] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][13] ),
    .X(_02087_));
 sky130_fd_sc_hd__a22o_1 _13665_ (.A1(\fifo_bank_register.bank[1][13] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][13] ),
    .X(_02088_));
 sky130_fd_sc_hd__a2111o_1 _13666_ (.A1(\fifo_bank_register.bank[9][13] ),
    .A2(_08190_),
    .B1(_02086_),
    .C1(_02087_),
    .D1(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__mux2_1 _13667_ (.A0(\fifo_bank_register.bank[0][13] ),
    .A1(_02089_),
    .S(_02068_),
    .X(_02090_));
 sky130_fd_sc_hd__mux2_1 _13668_ (.A0(_02090_),
    .A1(\fifo_bank_register.data_out[13] ),
    .S(_08172_),
    .X(_02091_));
 sky130_fd_sc_hd__clkbuf_1 _13669_ (.A(_02091_),
    .X(_01454_));
 sky130_fd_sc_hd__a22o_1 _13670_ (.A1(\fifo_bank_register.bank[5][14] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][14] ),
    .X(_02092_));
 sky130_fd_sc_hd__a221o_1 _13671_ (.A1(\fifo_bank_register.bank[7][14] ),
    .A2(_08182_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][14] ),
    .C1(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__a22o_1 _13672_ (.A1(\fifo_bank_register.bank[6][14] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][14] ),
    .X(_02094_));
 sky130_fd_sc_hd__a22o_1 _13673_ (.A1(\fifo_bank_register.bank[1][14] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][14] ),
    .X(_02095_));
 sky130_fd_sc_hd__a2111o_1 _13674_ (.A1(\fifo_bank_register.bank[9][14] ),
    .A2(_08190_),
    .B1(_02093_),
    .C1(_02094_),
    .D1(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__mux2_1 _13675_ (.A0(\fifo_bank_register.bank[0][14] ),
    .A1(_02096_),
    .S(_02068_),
    .X(_02097_));
 sky130_fd_sc_hd__mux2_1 _13676_ (.A0(_02097_),
    .A1(\fifo_bank_register.data_out[14] ),
    .S(_08172_),
    .X(_02098_));
 sky130_fd_sc_hd__clkbuf_1 _13677_ (.A(_02098_),
    .X(_01455_));
 sky130_fd_sc_hd__a22o_1 _13678_ (.A1(\fifo_bank_register.bank[5][15] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][15] ),
    .X(_02099_));
 sky130_fd_sc_hd__a221o_1 _13679_ (.A1(\fifo_bank_register.bank[7][15] ),
    .A2(_08182_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][15] ),
    .C1(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__a22o_1 _13680_ (.A1(\fifo_bank_register.bank[6][15] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][15] ),
    .X(_02101_));
 sky130_fd_sc_hd__a22o_1 _13681_ (.A1(\fifo_bank_register.bank[1][15] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][15] ),
    .X(_02102_));
 sky130_fd_sc_hd__a2111o_1 _13682_ (.A1(\fifo_bank_register.bank[9][15] ),
    .A2(_08190_),
    .B1(_02100_),
    .C1(_02101_),
    .D1(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__mux2_1 _13683_ (.A0(\fifo_bank_register.bank[0][15] ),
    .A1(_02103_),
    .S(_02068_),
    .X(_02104_));
 sky130_fd_sc_hd__mux2_1 _13684_ (.A0(_02104_),
    .A1(\fifo_bank_register.data_out[15] ),
    .S(_08172_),
    .X(_02105_));
 sky130_fd_sc_hd__clkbuf_1 _13685_ (.A(_02105_),
    .X(_01456_));
 sky130_fd_sc_hd__a22o_1 _13686_ (.A1(\fifo_bank_register.bank[5][16] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][16] ),
    .X(_02106_));
 sky130_fd_sc_hd__a221o_1 _13687_ (.A1(\fifo_bank_register.bank[7][16] ),
    .A2(_08182_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][16] ),
    .C1(_02106_),
    .X(_02107_));
 sky130_fd_sc_hd__a22o_1 _13688_ (.A1(\fifo_bank_register.bank[6][16] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][16] ),
    .X(_02108_));
 sky130_fd_sc_hd__a22o_1 _13689_ (.A1(\fifo_bank_register.bank[1][16] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][16] ),
    .X(_02109_));
 sky130_fd_sc_hd__a2111o_1 _13690_ (.A1(\fifo_bank_register.bank[9][16] ),
    .A2(_08190_),
    .B1(_02107_),
    .C1(_02108_),
    .D1(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__mux2_1 _13691_ (.A0(\fifo_bank_register.bank[0][16] ),
    .A1(_02110_),
    .S(_02068_),
    .X(_02111_));
 sky130_fd_sc_hd__mux2_1 _13692_ (.A0(_02111_),
    .A1(\fifo_bank_register.data_out[16] ),
    .S(_08172_),
    .X(_02112_));
 sky130_fd_sc_hd__clkbuf_1 _13693_ (.A(_02112_),
    .X(_01457_));
 sky130_fd_sc_hd__a22o_1 _13694_ (.A1(\fifo_bank_register.bank[5][17] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][17] ),
    .X(_02113_));
 sky130_fd_sc_hd__a221o_1 _13695_ (.A1(\fifo_bank_register.bank[7][17] ),
    .A2(_08182_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][17] ),
    .C1(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__a22o_1 _13696_ (.A1(\fifo_bank_register.bank[6][17] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][17] ),
    .X(_02115_));
 sky130_fd_sc_hd__a22o_1 _13697_ (.A1(\fifo_bank_register.bank[1][17] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][17] ),
    .X(_02116_));
 sky130_fd_sc_hd__a2111o_1 _13698_ (.A1(\fifo_bank_register.bank[9][17] ),
    .A2(_08190_),
    .B1(_02114_),
    .C1(_02115_),
    .D1(_02116_),
    .X(_02117_));
 sky130_fd_sc_hd__mux2_1 _13699_ (.A0(\fifo_bank_register.bank[0][17] ),
    .A1(_02117_),
    .S(_02068_),
    .X(_02118_));
 sky130_fd_sc_hd__clkbuf_8 _13700_ (.A(_08068_),
    .X(_02119_));
 sky130_fd_sc_hd__mux2_1 _13701_ (.A0(_02118_),
    .A1(\fifo_bank_register.data_out[17] ),
    .S(_02119_),
    .X(_02120_));
 sky130_fd_sc_hd__clkbuf_1 _13702_ (.A(_02120_),
    .X(_01458_));
 sky130_fd_sc_hd__a22o_1 _13703_ (.A1(\fifo_bank_register.bank[5][18] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][18] ),
    .X(_02121_));
 sky130_fd_sc_hd__a221o_1 _13704_ (.A1(\fifo_bank_register.bank[7][18] ),
    .A2(_08182_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][18] ),
    .C1(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__a22o_1 _13705_ (.A1(\fifo_bank_register.bank[6][18] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][18] ),
    .X(_02123_));
 sky130_fd_sc_hd__a22o_1 _13706_ (.A1(\fifo_bank_register.bank[1][18] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][18] ),
    .X(_02124_));
 sky130_fd_sc_hd__a2111o_1 _13707_ (.A1(\fifo_bank_register.bank[9][18] ),
    .A2(_08190_),
    .B1(_02122_),
    .C1(_02123_),
    .D1(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__mux2_1 _13708_ (.A0(\fifo_bank_register.bank[0][18] ),
    .A1(_02125_),
    .S(_02068_),
    .X(_02126_));
 sky130_fd_sc_hd__mux2_1 _13709_ (.A0(_02126_),
    .A1(\fifo_bank_register.data_out[18] ),
    .S(_02119_),
    .X(_02127_));
 sky130_fd_sc_hd__clkbuf_1 _13710_ (.A(_02127_),
    .X(_01459_));
 sky130_fd_sc_hd__clkbuf_4 _13711_ (.A(_08181_),
    .X(_02128_));
 sky130_fd_sc_hd__a22o_1 _13712_ (.A1(\fifo_bank_register.bank[5][19] ),
    .A2(_08192_),
    .B1(_08193_),
    .B2(\fifo_bank_register.bank[3][19] ),
    .X(_02129_));
 sky130_fd_sc_hd__a221o_1 _13713_ (.A1(\fifo_bank_register.bank[7][19] ),
    .A2(_02128_),
    .B1(_08191_),
    .B2(\fifo_bank_register.bank[2][19] ),
    .C1(_02129_),
    .X(_02130_));
 sky130_fd_sc_hd__a22o_1 _13714_ (.A1(\fifo_bank_register.bank[6][19] ),
    .A2(_08196_),
    .B1(_08197_),
    .B2(\fifo_bank_register.bank[4][19] ),
    .X(_02131_));
 sky130_fd_sc_hd__a22o_1 _13715_ (.A1(\fifo_bank_register.bank[1][19] ),
    .A2(_08199_),
    .B1(_08200_),
    .B2(\fifo_bank_register.bank[8][19] ),
    .X(_02132_));
 sky130_fd_sc_hd__a2111o_1 _13716_ (.A1(\fifo_bank_register.bank[9][19] ),
    .A2(_08190_),
    .B1(_02130_),
    .C1(_02131_),
    .D1(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__mux2_1 _13717_ (.A0(\fifo_bank_register.bank[0][19] ),
    .A1(_02133_),
    .S(_02068_),
    .X(_02134_));
 sky130_fd_sc_hd__mux2_1 _13718_ (.A0(_02134_),
    .A1(\fifo_bank_register.data_out[19] ),
    .S(_02119_),
    .X(_02135_));
 sky130_fd_sc_hd__clkbuf_1 _13719_ (.A(_02135_),
    .X(_01460_));
 sky130_fd_sc_hd__clkbuf_8 _13720_ (.A(_08088_),
    .X(_02136_));
 sky130_fd_sc_hd__buf_4 _13721_ (.A(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__buf_6 _13722_ (.A(_08091_),
    .X(_02138_));
 sky130_fd_sc_hd__clkbuf_4 _13723_ (.A(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__buf_6 _13724_ (.A(_08095_),
    .X(_02140_));
 sky130_fd_sc_hd__clkbuf_4 _13725_ (.A(_02140_),
    .X(_02141_));
 sky130_fd_sc_hd__buf_6 _13726_ (.A(_08098_),
    .X(_02142_));
 sky130_fd_sc_hd__clkbuf_4 _13727_ (.A(_02142_),
    .X(_02143_));
 sky130_fd_sc_hd__a22o_1 _13728_ (.A1(\fifo_bank_register.bank[5][20] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][20] ),
    .X(_02144_));
 sky130_fd_sc_hd__a221o_1 _13729_ (.A1(\fifo_bank_register.bank[7][20] ),
    .A2(_02128_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][20] ),
    .C1(_02144_),
    .X(_02145_));
 sky130_fd_sc_hd__buf_6 _13730_ (.A(_08103_),
    .X(_02146_));
 sky130_fd_sc_hd__clkbuf_4 _13731_ (.A(_02146_),
    .X(_02147_));
 sky130_fd_sc_hd__buf_6 _13732_ (.A(_08106_),
    .X(_02148_));
 sky130_fd_sc_hd__clkbuf_4 _13733_ (.A(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__a22o_1 _13734_ (.A1(\fifo_bank_register.bank[6][20] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][20] ),
    .X(_02150_));
 sky130_fd_sc_hd__buf_6 _13735_ (.A(_08110_),
    .X(_02151_));
 sky130_fd_sc_hd__clkbuf_4 _13736_ (.A(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__buf_6 _13737_ (.A(_08113_),
    .X(_02153_));
 sky130_fd_sc_hd__clkbuf_4 _13738_ (.A(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__a22o_1 _13739_ (.A1(\fifo_bank_register.bank[1][20] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][20] ),
    .X(_02155_));
 sky130_fd_sc_hd__a2111o_1 _13740_ (.A1(\fifo_bank_register.bank[9][20] ),
    .A2(_02137_),
    .B1(_02145_),
    .C1(_02150_),
    .D1(_02155_),
    .X(_02156_));
 sky130_fd_sc_hd__clkbuf_8 _13741_ (.A(_08119_),
    .X(_02157_));
 sky130_fd_sc_hd__buf_4 _13742_ (.A(_02157_),
    .X(_02158_));
 sky130_fd_sc_hd__mux2_1 _13743_ (.A0(\fifo_bank_register.bank[0][20] ),
    .A1(_02156_),
    .S(_02158_),
    .X(_02159_));
 sky130_fd_sc_hd__mux2_1 _13744_ (.A0(_02159_),
    .A1(\fifo_bank_register.data_out[20] ),
    .S(_02119_),
    .X(_02160_));
 sky130_fd_sc_hd__clkbuf_1 _13745_ (.A(_02160_),
    .X(_01461_));
 sky130_fd_sc_hd__a22o_1 _13746_ (.A1(\fifo_bank_register.bank[5][21] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][21] ),
    .X(_02161_));
 sky130_fd_sc_hd__a221o_1 _13747_ (.A1(\fifo_bank_register.bank[7][21] ),
    .A2(_02128_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][21] ),
    .C1(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__a22o_1 _13748_ (.A1(\fifo_bank_register.bank[6][21] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][21] ),
    .X(_02163_));
 sky130_fd_sc_hd__a22o_1 _13749_ (.A1(\fifo_bank_register.bank[1][21] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][21] ),
    .X(_02164_));
 sky130_fd_sc_hd__a2111o_1 _13750_ (.A1(\fifo_bank_register.bank[9][21] ),
    .A2(_02137_),
    .B1(_02162_),
    .C1(_02163_),
    .D1(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__mux2_1 _13751_ (.A0(\fifo_bank_register.bank[0][21] ),
    .A1(_02165_),
    .S(_02158_),
    .X(_02166_));
 sky130_fd_sc_hd__mux2_1 _13752_ (.A0(_02166_),
    .A1(\fifo_bank_register.data_out[21] ),
    .S(_02119_),
    .X(_02167_));
 sky130_fd_sc_hd__clkbuf_1 _13753_ (.A(_02167_),
    .X(_01462_));
 sky130_fd_sc_hd__a22o_1 _13754_ (.A1(\fifo_bank_register.bank[5][22] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][22] ),
    .X(_02168_));
 sky130_fd_sc_hd__a221o_1 _13755_ (.A1(\fifo_bank_register.bank[7][22] ),
    .A2(_02128_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][22] ),
    .C1(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _13756_ (.A1(\fifo_bank_register.bank[6][22] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][22] ),
    .X(_02170_));
 sky130_fd_sc_hd__a22o_1 _13757_ (.A1(\fifo_bank_register.bank[1][22] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][22] ),
    .X(_02171_));
 sky130_fd_sc_hd__a2111o_1 _13758_ (.A1(\fifo_bank_register.bank[9][22] ),
    .A2(_02137_),
    .B1(_02169_),
    .C1(_02170_),
    .D1(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__mux2_1 _13759_ (.A0(\fifo_bank_register.bank[0][22] ),
    .A1(_02172_),
    .S(_02158_),
    .X(_02173_));
 sky130_fd_sc_hd__mux2_1 _13760_ (.A0(_02173_),
    .A1(\fifo_bank_register.data_out[22] ),
    .S(_02119_),
    .X(_02174_));
 sky130_fd_sc_hd__clkbuf_1 _13761_ (.A(_02174_),
    .X(_01463_));
 sky130_fd_sc_hd__a22o_1 _13762_ (.A1(\fifo_bank_register.bank[5][23] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][23] ),
    .X(_02175_));
 sky130_fd_sc_hd__a221o_1 _13763_ (.A1(\fifo_bank_register.bank[7][23] ),
    .A2(_02128_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][23] ),
    .C1(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__a22o_1 _13764_ (.A1(\fifo_bank_register.bank[6][23] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][23] ),
    .X(_02177_));
 sky130_fd_sc_hd__a22o_1 _13765_ (.A1(\fifo_bank_register.bank[1][23] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][23] ),
    .X(_02178_));
 sky130_fd_sc_hd__a2111o_1 _13766_ (.A1(\fifo_bank_register.bank[9][23] ),
    .A2(_02137_),
    .B1(_02176_),
    .C1(_02177_),
    .D1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__mux2_1 _13767_ (.A0(\fifo_bank_register.bank[0][23] ),
    .A1(_02179_),
    .S(_02158_),
    .X(_02180_));
 sky130_fd_sc_hd__mux2_1 _13768_ (.A0(_02180_),
    .A1(\fifo_bank_register.data_out[23] ),
    .S(_02119_),
    .X(_02181_));
 sky130_fd_sc_hd__clkbuf_1 _13769_ (.A(_02181_),
    .X(_01464_));
 sky130_fd_sc_hd__a22o_1 _13770_ (.A1(\fifo_bank_register.bank[5][24] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][24] ),
    .X(_02182_));
 sky130_fd_sc_hd__a221o_1 _13771_ (.A1(\fifo_bank_register.bank[7][24] ),
    .A2(_02128_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][24] ),
    .C1(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__a22o_1 _13772_ (.A1(\fifo_bank_register.bank[6][24] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][24] ),
    .X(_02184_));
 sky130_fd_sc_hd__a22o_1 _13773_ (.A1(\fifo_bank_register.bank[1][24] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][24] ),
    .X(_02185_));
 sky130_fd_sc_hd__a2111o_1 _13774_ (.A1(\fifo_bank_register.bank[9][24] ),
    .A2(_02137_),
    .B1(_02183_),
    .C1(_02184_),
    .D1(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__mux2_1 _13775_ (.A0(\fifo_bank_register.bank[0][24] ),
    .A1(_02186_),
    .S(_02158_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _13776_ (.A0(_02187_),
    .A1(\fifo_bank_register.data_out[24] ),
    .S(_02119_),
    .X(_02188_));
 sky130_fd_sc_hd__clkbuf_1 _13777_ (.A(_02188_),
    .X(_01465_));
 sky130_fd_sc_hd__a22o_1 _13778_ (.A1(\fifo_bank_register.bank[5][25] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][25] ),
    .X(_02189_));
 sky130_fd_sc_hd__a221o_1 _13779_ (.A1(\fifo_bank_register.bank[7][25] ),
    .A2(_02128_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][25] ),
    .C1(_02189_),
    .X(_02190_));
 sky130_fd_sc_hd__a22o_1 _13780_ (.A1(\fifo_bank_register.bank[6][25] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][25] ),
    .X(_02191_));
 sky130_fd_sc_hd__a22o_1 _13781_ (.A1(\fifo_bank_register.bank[1][25] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][25] ),
    .X(_02192_));
 sky130_fd_sc_hd__a2111o_1 _13782_ (.A1(\fifo_bank_register.bank[9][25] ),
    .A2(_02137_),
    .B1(_02190_),
    .C1(_02191_),
    .D1(_02192_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _13783_ (.A0(\fifo_bank_register.bank[0][25] ),
    .A1(_02193_),
    .S(_02158_),
    .X(_02194_));
 sky130_fd_sc_hd__mux2_1 _13784_ (.A0(_02194_),
    .A1(\fifo_bank_register.data_out[25] ),
    .S(_02119_),
    .X(_02195_));
 sky130_fd_sc_hd__clkbuf_1 _13785_ (.A(_02195_),
    .X(_01466_));
 sky130_fd_sc_hd__a22o_1 _13786_ (.A1(\fifo_bank_register.bank[5][26] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][26] ),
    .X(_02196_));
 sky130_fd_sc_hd__a221o_1 _13787_ (.A1(\fifo_bank_register.bank[7][26] ),
    .A2(_02128_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][26] ),
    .C1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__a22o_1 _13788_ (.A1(\fifo_bank_register.bank[6][26] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][26] ),
    .X(_02198_));
 sky130_fd_sc_hd__a22o_1 _13789_ (.A1(\fifo_bank_register.bank[1][26] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][26] ),
    .X(_02199_));
 sky130_fd_sc_hd__a2111o_1 _13790_ (.A1(\fifo_bank_register.bank[9][26] ),
    .A2(_02137_),
    .B1(_02197_),
    .C1(_02198_),
    .D1(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _13791_ (.A0(\fifo_bank_register.bank[0][26] ),
    .A1(_02200_),
    .S(_02158_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _13792_ (.A0(_02201_),
    .A1(\fifo_bank_register.data_out[26] ),
    .S(_02119_),
    .X(_02202_));
 sky130_fd_sc_hd__clkbuf_1 _13793_ (.A(_02202_),
    .X(_01467_));
 sky130_fd_sc_hd__a22o_1 _13794_ (.A1(\fifo_bank_register.bank[5][27] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][27] ),
    .X(_02203_));
 sky130_fd_sc_hd__a221o_1 _13795_ (.A1(\fifo_bank_register.bank[7][27] ),
    .A2(_02128_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][27] ),
    .C1(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__a22o_1 _13796_ (.A1(\fifo_bank_register.bank[6][27] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][27] ),
    .X(_02205_));
 sky130_fd_sc_hd__a22o_1 _13797_ (.A1(\fifo_bank_register.bank[1][27] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][27] ),
    .X(_02206_));
 sky130_fd_sc_hd__a2111o_1 _13798_ (.A1(\fifo_bank_register.bank[9][27] ),
    .A2(_02137_),
    .B1(_02204_),
    .C1(_02205_),
    .D1(_02206_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _13799_ (.A0(\fifo_bank_register.bank[0][27] ),
    .A1(_02207_),
    .S(_02158_),
    .X(_02208_));
 sky130_fd_sc_hd__buf_4 _13800_ (.A(_08068_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _13801_ (.A0(_02208_),
    .A1(\fifo_bank_register.data_out[27] ),
    .S(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__clkbuf_1 _13802_ (.A(_02210_),
    .X(_01468_));
 sky130_fd_sc_hd__a22o_1 _13803_ (.A1(\fifo_bank_register.bank[5][28] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][28] ),
    .X(_02211_));
 sky130_fd_sc_hd__a221o_1 _13804_ (.A1(\fifo_bank_register.bank[7][28] ),
    .A2(_02128_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][28] ),
    .C1(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__a22o_1 _13805_ (.A1(\fifo_bank_register.bank[6][28] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][28] ),
    .X(_02213_));
 sky130_fd_sc_hd__a22o_1 _13806_ (.A1(\fifo_bank_register.bank[1][28] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][28] ),
    .X(_02214_));
 sky130_fd_sc_hd__a2111o_1 _13807_ (.A1(\fifo_bank_register.bank[9][28] ),
    .A2(_02137_),
    .B1(_02212_),
    .C1(_02213_),
    .D1(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_1 _13808_ (.A0(\fifo_bank_register.bank[0][28] ),
    .A1(_02215_),
    .S(_02158_),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _13809_ (.A0(_02216_),
    .A1(\fifo_bank_register.data_out[28] ),
    .S(_02209_),
    .X(_02217_));
 sky130_fd_sc_hd__clkbuf_1 _13810_ (.A(_02217_),
    .X(_01469_));
 sky130_fd_sc_hd__buf_4 _13811_ (.A(_08181_),
    .X(_02218_));
 sky130_fd_sc_hd__a22o_1 _13812_ (.A1(\fifo_bank_register.bank[5][29] ),
    .A2(_02141_),
    .B1(_02143_),
    .B2(\fifo_bank_register.bank[3][29] ),
    .X(_02219_));
 sky130_fd_sc_hd__a221o_1 _13813_ (.A1(\fifo_bank_register.bank[7][29] ),
    .A2(_02218_),
    .B1(_02139_),
    .B2(\fifo_bank_register.bank[2][29] ),
    .C1(_02219_),
    .X(_02220_));
 sky130_fd_sc_hd__a22o_1 _13814_ (.A1(\fifo_bank_register.bank[6][29] ),
    .A2(_02147_),
    .B1(_02149_),
    .B2(\fifo_bank_register.bank[4][29] ),
    .X(_02221_));
 sky130_fd_sc_hd__a22o_1 _13815_ (.A1(\fifo_bank_register.bank[1][29] ),
    .A2(_02152_),
    .B1(_02154_),
    .B2(\fifo_bank_register.bank[8][29] ),
    .X(_02222_));
 sky130_fd_sc_hd__a2111o_1 _13816_ (.A1(\fifo_bank_register.bank[9][29] ),
    .A2(_02137_),
    .B1(_02220_),
    .C1(_02221_),
    .D1(_02222_),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _13817_ (.A0(\fifo_bank_register.bank[0][29] ),
    .A1(_02223_),
    .S(_02158_),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _13818_ (.A0(_02224_),
    .A1(\fifo_bank_register.data_out[29] ),
    .S(_02209_),
    .X(_02225_));
 sky130_fd_sc_hd__clkbuf_1 _13819_ (.A(_02225_),
    .X(_01470_));
 sky130_fd_sc_hd__clkbuf_4 _13820_ (.A(_02136_),
    .X(_02226_));
 sky130_fd_sc_hd__clkbuf_4 _13821_ (.A(_02138_),
    .X(_02227_));
 sky130_fd_sc_hd__clkbuf_4 _13822_ (.A(_02140_),
    .X(_02228_));
 sky130_fd_sc_hd__clkbuf_4 _13823_ (.A(_02142_),
    .X(_02229_));
 sky130_fd_sc_hd__a22o_1 _13824_ (.A1(\fifo_bank_register.bank[5][30] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][30] ),
    .X(_02230_));
 sky130_fd_sc_hd__a221o_1 _13825_ (.A1(\fifo_bank_register.bank[7][30] ),
    .A2(_02218_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][30] ),
    .C1(_02230_),
    .X(_02231_));
 sky130_fd_sc_hd__clkbuf_4 _13826_ (.A(_02146_),
    .X(_02232_));
 sky130_fd_sc_hd__clkbuf_4 _13827_ (.A(_02148_),
    .X(_02233_));
 sky130_fd_sc_hd__a22o_1 _13828_ (.A1(\fifo_bank_register.bank[6][30] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][30] ),
    .X(_02234_));
 sky130_fd_sc_hd__clkbuf_4 _13829_ (.A(_02151_),
    .X(_02235_));
 sky130_fd_sc_hd__clkbuf_4 _13830_ (.A(_02153_),
    .X(_02236_));
 sky130_fd_sc_hd__a22o_1 _13831_ (.A1(\fifo_bank_register.bank[1][30] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][30] ),
    .X(_02237_));
 sky130_fd_sc_hd__a2111o_1 _13832_ (.A1(\fifo_bank_register.bank[9][30] ),
    .A2(_02226_),
    .B1(_02231_),
    .C1(_02234_),
    .D1(_02237_),
    .X(_02238_));
 sky130_fd_sc_hd__buf_4 _13833_ (.A(_02157_),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _13834_ (.A0(\fifo_bank_register.bank[0][30] ),
    .A1(_02238_),
    .S(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_1 _13835_ (.A0(_02240_),
    .A1(\fifo_bank_register.data_out[30] ),
    .S(_02209_),
    .X(_02241_));
 sky130_fd_sc_hd__clkbuf_1 _13836_ (.A(_02241_),
    .X(_01471_));
 sky130_fd_sc_hd__a22o_1 _13837_ (.A1(\fifo_bank_register.bank[5][31] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][31] ),
    .X(_02242_));
 sky130_fd_sc_hd__a221o_1 _13838_ (.A1(\fifo_bank_register.bank[7][31] ),
    .A2(_02218_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][31] ),
    .C1(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__a22o_1 _13839_ (.A1(\fifo_bank_register.bank[6][31] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][31] ),
    .X(_02244_));
 sky130_fd_sc_hd__a22o_1 _13840_ (.A1(\fifo_bank_register.bank[1][31] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][31] ),
    .X(_02245_));
 sky130_fd_sc_hd__a2111o_1 _13841_ (.A1(\fifo_bank_register.bank[9][31] ),
    .A2(_02226_),
    .B1(_02243_),
    .C1(_02244_),
    .D1(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _13842_ (.A0(\fifo_bank_register.bank[0][31] ),
    .A1(_02246_),
    .S(_02239_),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _13843_ (.A0(_02247_),
    .A1(\fifo_bank_register.data_out[31] ),
    .S(_02209_),
    .X(_02248_));
 sky130_fd_sc_hd__clkbuf_1 _13844_ (.A(_02248_),
    .X(_01472_));
 sky130_fd_sc_hd__a22o_1 _13845_ (.A1(\fifo_bank_register.bank[5][32] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][32] ),
    .X(_02249_));
 sky130_fd_sc_hd__a221o_1 _13846_ (.A1(\fifo_bank_register.bank[7][32] ),
    .A2(_02218_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][32] ),
    .C1(_02249_),
    .X(_02250_));
 sky130_fd_sc_hd__a22o_1 _13847_ (.A1(\fifo_bank_register.bank[6][32] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][32] ),
    .X(_02251_));
 sky130_fd_sc_hd__a22o_1 _13848_ (.A1(\fifo_bank_register.bank[1][32] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][32] ),
    .X(_02252_));
 sky130_fd_sc_hd__a2111o_1 _13849_ (.A1(\fifo_bank_register.bank[9][32] ),
    .A2(_02226_),
    .B1(_02250_),
    .C1(_02251_),
    .D1(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _13850_ (.A0(\fifo_bank_register.bank[0][32] ),
    .A1(_02253_),
    .S(_02239_),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _13851_ (.A0(_02254_),
    .A1(\fifo_bank_register.data_out[32] ),
    .S(_02209_),
    .X(_02255_));
 sky130_fd_sc_hd__clkbuf_1 _13852_ (.A(_02255_),
    .X(_01473_));
 sky130_fd_sc_hd__a22o_1 _13853_ (.A1(\fifo_bank_register.bank[5][33] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][33] ),
    .X(_02256_));
 sky130_fd_sc_hd__a221o_1 _13854_ (.A1(\fifo_bank_register.bank[7][33] ),
    .A2(_02218_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][33] ),
    .C1(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__a22o_1 _13855_ (.A1(\fifo_bank_register.bank[6][33] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][33] ),
    .X(_02258_));
 sky130_fd_sc_hd__a22o_1 _13856_ (.A1(\fifo_bank_register.bank[1][33] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][33] ),
    .X(_02259_));
 sky130_fd_sc_hd__a2111o_1 _13857_ (.A1(\fifo_bank_register.bank[9][33] ),
    .A2(_02226_),
    .B1(_02257_),
    .C1(_02258_),
    .D1(_02259_),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _13858_ (.A0(\fifo_bank_register.bank[0][33] ),
    .A1(_02260_),
    .S(_02239_),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _13859_ (.A0(_02261_),
    .A1(\fifo_bank_register.data_out[33] ),
    .S(_02209_),
    .X(_02262_));
 sky130_fd_sc_hd__clkbuf_1 _13860_ (.A(_02262_),
    .X(_01474_));
 sky130_fd_sc_hd__a22o_1 _13861_ (.A1(\fifo_bank_register.bank[5][34] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][34] ),
    .X(_02263_));
 sky130_fd_sc_hd__a221o_1 _13862_ (.A1(\fifo_bank_register.bank[7][34] ),
    .A2(_02218_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][34] ),
    .C1(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__a22o_1 _13863_ (.A1(\fifo_bank_register.bank[6][34] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][34] ),
    .X(_02265_));
 sky130_fd_sc_hd__a22o_1 _13864_ (.A1(\fifo_bank_register.bank[1][34] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][34] ),
    .X(_02266_));
 sky130_fd_sc_hd__a2111o_1 _13865_ (.A1(\fifo_bank_register.bank[9][34] ),
    .A2(_02226_),
    .B1(_02264_),
    .C1(_02265_),
    .D1(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _13866_ (.A0(\fifo_bank_register.bank[0][34] ),
    .A1(_02267_),
    .S(_02239_),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _13867_ (.A0(_02268_),
    .A1(\fifo_bank_register.data_out[34] ),
    .S(_02209_),
    .X(_02269_));
 sky130_fd_sc_hd__clkbuf_1 _13868_ (.A(_02269_),
    .X(_01475_));
 sky130_fd_sc_hd__a22o_1 _13869_ (.A1(\fifo_bank_register.bank[5][35] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][35] ),
    .X(_02270_));
 sky130_fd_sc_hd__a221o_1 _13870_ (.A1(\fifo_bank_register.bank[7][35] ),
    .A2(_02218_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][35] ),
    .C1(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__a22o_1 _13871_ (.A1(\fifo_bank_register.bank[6][35] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][35] ),
    .X(_02272_));
 sky130_fd_sc_hd__a22o_1 _13872_ (.A1(\fifo_bank_register.bank[1][35] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][35] ),
    .X(_02273_));
 sky130_fd_sc_hd__a2111o_1 _13873_ (.A1(\fifo_bank_register.bank[9][35] ),
    .A2(_02226_),
    .B1(_02271_),
    .C1(_02272_),
    .D1(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _13874_ (.A0(\fifo_bank_register.bank[0][35] ),
    .A1(_02274_),
    .S(_02239_),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _13875_ (.A0(_02275_),
    .A1(\fifo_bank_register.data_out[35] ),
    .S(_02209_),
    .X(_02276_));
 sky130_fd_sc_hd__clkbuf_1 _13876_ (.A(_02276_),
    .X(_01476_));
 sky130_fd_sc_hd__a22o_1 _13877_ (.A1(\fifo_bank_register.bank[5][36] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][36] ),
    .X(_02277_));
 sky130_fd_sc_hd__a221o_1 _13878_ (.A1(\fifo_bank_register.bank[7][36] ),
    .A2(_02218_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][36] ),
    .C1(_02277_),
    .X(_02278_));
 sky130_fd_sc_hd__a22o_1 _13879_ (.A1(\fifo_bank_register.bank[6][36] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][36] ),
    .X(_02279_));
 sky130_fd_sc_hd__a22o_1 _13880_ (.A1(\fifo_bank_register.bank[1][36] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][36] ),
    .X(_02280_));
 sky130_fd_sc_hd__a2111o_1 _13881_ (.A1(\fifo_bank_register.bank[9][36] ),
    .A2(_02226_),
    .B1(_02278_),
    .C1(_02279_),
    .D1(_02280_),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _13882_ (.A0(\fifo_bank_register.bank[0][36] ),
    .A1(_02281_),
    .S(_02239_),
    .X(_02282_));
 sky130_fd_sc_hd__mux2_1 _13883_ (.A0(_02282_),
    .A1(\fifo_bank_register.data_out[36] ),
    .S(_02209_),
    .X(_02283_));
 sky130_fd_sc_hd__clkbuf_1 _13884_ (.A(_02283_),
    .X(_01477_));
 sky130_fd_sc_hd__a22o_1 _13885_ (.A1(\fifo_bank_register.bank[5][37] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][37] ),
    .X(_02284_));
 sky130_fd_sc_hd__a221o_1 _13886_ (.A1(\fifo_bank_register.bank[7][37] ),
    .A2(_02218_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][37] ),
    .C1(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__a22o_1 _13887_ (.A1(\fifo_bank_register.bank[6][37] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][37] ),
    .X(_02286_));
 sky130_fd_sc_hd__a22o_1 _13888_ (.A1(\fifo_bank_register.bank[1][37] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][37] ),
    .X(_02287_));
 sky130_fd_sc_hd__a2111o_1 _13889_ (.A1(\fifo_bank_register.bank[9][37] ),
    .A2(_02226_),
    .B1(_02285_),
    .C1(_02286_),
    .D1(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _13890_ (.A0(\fifo_bank_register.bank[0][37] ),
    .A1(_02288_),
    .S(_02239_),
    .X(_02289_));
 sky130_fd_sc_hd__buf_4 _13891_ (.A(_08068_),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _13892_ (.A0(_02289_),
    .A1(\fifo_bank_register.data_out[37] ),
    .S(_02290_),
    .X(_02291_));
 sky130_fd_sc_hd__clkbuf_1 _13893_ (.A(_02291_),
    .X(_01478_));
 sky130_fd_sc_hd__a22o_1 _13894_ (.A1(\fifo_bank_register.bank[5][38] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][38] ),
    .X(_02292_));
 sky130_fd_sc_hd__a221o_1 _13895_ (.A1(\fifo_bank_register.bank[7][38] ),
    .A2(_02218_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][38] ),
    .C1(_02292_),
    .X(_02293_));
 sky130_fd_sc_hd__a22o_1 _13896_ (.A1(\fifo_bank_register.bank[6][38] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][38] ),
    .X(_02294_));
 sky130_fd_sc_hd__a22o_1 _13897_ (.A1(\fifo_bank_register.bank[1][38] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][38] ),
    .X(_02295_));
 sky130_fd_sc_hd__a2111o_1 _13898_ (.A1(\fifo_bank_register.bank[9][38] ),
    .A2(_02226_),
    .B1(_02293_),
    .C1(_02294_),
    .D1(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__mux2_1 _13899_ (.A0(\fifo_bank_register.bank[0][38] ),
    .A1(_02296_),
    .S(_02239_),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _13900_ (.A0(_02297_),
    .A1(\fifo_bank_register.data_out[38] ),
    .S(_02290_),
    .X(_02298_));
 sky130_fd_sc_hd__clkbuf_1 _13901_ (.A(_02298_),
    .X(_01479_));
 sky130_fd_sc_hd__clkbuf_4 _13902_ (.A(_08181_),
    .X(_02299_));
 sky130_fd_sc_hd__a22o_1 _13903_ (.A1(\fifo_bank_register.bank[5][39] ),
    .A2(_02228_),
    .B1(_02229_),
    .B2(\fifo_bank_register.bank[3][39] ),
    .X(_02300_));
 sky130_fd_sc_hd__a221o_1 _13904_ (.A1(\fifo_bank_register.bank[7][39] ),
    .A2(_02299_),
    .B1(_02227_),
    .B2(\fifo_bank_register.bank[2][39] ),
    .C1(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__a22o_1 _13905_ (.A1(\fifo_bank_register.bank[6][39] ),
    .A2(_02232_),
    .B1(_02233_),
    .B2(\fifo_bank_register.bank[4][39] ),
    .X(_02302_));
 sky130_fd_sc_hd__a22o_1 _13906_ (.A1(\fifo_bank_register.bank[1][39] ),
    .A2(_02235_),
    .B1(_02236_),
    .B2(\fifo_bank_register.bank[8][39] ),
    .X(_02303_));
 sky130_fd_sc_hd__a2111o_1 _13907_ (.A1(\fifo_bank_register.bank[9][39] ),
    .A2(_02226_),
    .B1(_02301_),
    .C1(_02302_),
    .D1(_02303_),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _13908_ (.A0(\fifo_bank_register.bank[0][39] ),
    .A1(_02304_),
    .S(_02239_),
    .X(_02305_));
 sky130_fd_sc_hd__mux2_1 _13909_ (.A0(_02305_),
    .A1(\fifo_bank_register.data_out[39] ),
    .S(_02290_),
    .X(_02306_));
 sky130_fd_sc_hd__clkbuf_1 _13910_ (.A(_02306_),
    .X(_01480_));
 sky130_fd_sc_hd__clkbuf_4 _13911_ (.A(_02136_),
    .X(_02307_));
 sky130_fd_sc_hd__clkbuf_4 _13912_ (.A(_02138_),
    .X(_02308_));
 sky130_fd_sc_hd__clkbuf_4 _13913_ (.A(_02140_),
    .X(_02309_));
 sky130_fd_sc_hd__clkbuf_4 _13914_ (.A(_02142_),
    .X(_02310_));
 sky130_fd_sc_hd__a22o_1 _13915_ (.A1(\fifo_bank_register.bank[5][40] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][40] ),
    .X(_02311_));
 sky130_fd_sc_hd__a221o_1 _13916_ (.A1(\fifo_bank_register.bank[7][40] ),
    .A2(_02299_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][40] ),
    .C1(_02311_),
    .X(_02312_));
 sky130_fd_sc_hd__clkbuf_4 _13917_ (.A(_02146_),
    .X(_02313_));
 sky130_fd_sc_hd__clkbuf_4 _13918_ (.A(_02148_),
    .X(_02314_));
 sky130_fd_sc_hd__a22o_1 _13919_ (.A1(\fifo_bank_register.bank[6][40] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][40] ),
    .X(_02315_));
 sky130_fd_sc_hd__clkbuf_4 _13920_ (.A(_02151_),
    .X(_02316_));
 sky130_fd_sc_hd__clkbuf_4 _13921_ (.A(_02153_),
    .X(_02317_));
 sky130_fd_sc_hd__a22o_1 _13922_ (.A1(\fifo_bank_register.bank[1][40] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][40] ),
    .X(_02318_));
 sky130_fd_sc_hd__a2111o_1 _13923_ (.A1(\fifo_bank_register.bank[9][40] ),
    .A2(_02307_),
    .B1(_02312_),
    .C1(_02315_),
    .D1(_02318_),
    .X(_02319_));
 sky130_fd_sc_hd__buf_4 _13924_ (.A(_02157_),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _13925_ (.A0(\fifo_bank_register.bank[0][40] ),
    .A1(_02319_),
    .S(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__mux2_1 _13926_ (.A0(_02321_),
    .A1(\fifo_bank_register.data_out[40] ),
    .S(_02290_),
    .X(_02322_));
 sky130_fd_sc_hd__clkbuf_1 _13927_ (.A(_02322_),
    .X(_01481_));
 sky130_fd_sc_hd__a22o_1 _13928_ (.A1(\fifo_bank_register.bank[5][41] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][41] ),
    .X(_02323_));
 sky130_fd_sc_hd__a221o_1 _13929_ (.A1(\fifo_bank_register.bank[7][41] ),
    .A2(_02299_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][41] ),
    .C1(_02323_),
    .X(_02324_));
 sky130_fd_sc_hd__a22o_1 _13930_ (.A1(\fifo_bank_register.bank[6][41] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][41] ),
    .X(_02325_));
 sky130_fd_sc_hd__a22o_1 _13931_ (.A1(\fifo_bank_register.bank[1][41] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][41] ),
    .X(_02326_));
 sky130_fd_sc_hd__a2111o_1 _13932_ (.A1(\fifo_bank_register.bank[9][41] ),
    .A2(_02307_),
    .B1(_02324_),
    .C1(_02325_),
    .D1(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__mux2_1 _13933_ (.A0(\fifo_bank_register.bank[0][41] ),
    .A1(_02327_),
    .S(_02320_),
    .X(_02328_));
 sky130_fd_sc_hd__mux2_1 _13934_ (.A0(_02328_),
    .A1(\fifo_bank_register.data_out[41] ),
    .S(_02290_),
    .X(_02329_));
 sky130_fd_sc_hd__clkbuf_1 _13935_ (.A(_02329_),
    .X(_01482_));
 sky130_fd_sc_hd__a22o_1 _13936_ (.A1(\fifo_bank_register.bank[5][42] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][42] ),
    .X(_02330_));
 sky130_fd_sc_hd__a221o_1 _13937_ (.A1(\fifo_bank_register.bank[7][42] ),
    .A2(_02299_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][42] ),
    .C1(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__a22o_1 _13938_ (.A1(\fifo_bank_register.bank[6][42] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][42] ),
    .X(_02332_));
 sky130_fd_sc_hd__a22o_1 _13939_ (.A1(\fifo_bank_register.bank[1][42] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][42] ),
    .X(_02333_));
 sky130_fd_sc_hd__a2111o_1 _13940_ (.A1(\fifo_bank_register.bank[9][42] ),
    .A2(_02307_),
    .B1(_02331_),
    .C1(_02332_),
    .D1(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__mux2_1 _13941_ (.A0(\fifo_bank_register.bank[0][42] ),
    .A1(_02334_),
    .S(_02320_),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _13942_ (.A0(_02335_),
    .A1(\fifo_bank_register.data_out[42] ),
    .S(_02290_),
    .X(_02336_));
 sky130_fd_sc_hd__clkbuf_1 _13943_ (.A(_02336_),
    .X(_01483_));
 sky130_fd_sc_hd__a22o_1 _13944_ (.A1(\fifo_bank_register.bank[5][43] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][43] ),
    .X(_02337_));
 sky130_fd_sc_hd__a221o_1 _13945_ (.A1(\fifo_bank_register.bank[7][43] ),
    .A2(_02299_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][43] ),
    .C1(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__a22o_1 _13946_ (.A1(\fifo_bank_register.bank[6][43] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][43] ),
    .X(_02339_));
 sky130_fd_sc_hd__a22o_1 _13947_ (.A1(\fifo_bank_register.bank[1][43] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][43] ),
    .X(_02340_));
 sky130_fd_sc_hd__a2111o_1 _13948_ (.A1(\fifo_bank_register.bank[9][43] ),
    .A2(_02307_),
    .B1(_02338_),
    .C1(_02339_),
    .D1(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _13949_ (.A0(\fifo_bank_register.bank[0][43] ),
    .A1(_02341_),
    .S(_02320_),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _13950_ (.A0(_02342_),
    .A1(\fifo_bank_register.data_out[43] ),
    .S(_02290_),
    .X(_02343_));
 sky130_fd_sc_hd__clkbuf_1 _13951_ (.A(_02343_),
    .X(_01484_));
 sky130_fd_sc_hd__a22o_1 _13952_ (.A1(\fifo_bank_register.bank[5][44] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][44] ),
    .X(_02344_));
 sky130_fd_sc_hd__a221o_1 _13953_ (.A1(\fifo_bank_register.bank[7][44] ),
    .A2(_02299_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][44] ),
    .C1(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__a22o_1 _13954_ (.A1(\fifo_bank_register.bank[6][44] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][44] ),
    .X(_02346_));
 sky130_fd_sc_hd__a22o_1 _13955_ (.A1(\fifo_bank_register.bank[1][44] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][44] ),
    .X(_02347_));
 sky130_fd_sc_hd__a2111o_1 _13956_ (.A1(\fifo_bank_register.bank[9][44] ),
    .A2(_02307_),
    .B1(_02345_),
    .C1(_02346_),
    .D1(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__mux2_1 _13957_ (.A0(\fifo_bank_register.bank[0][44] ),
    .A1(_02348_),
    .S(_02320_),
    .X(_02349_));
 sky130_fd_sc_hd__mux2_1 _13958_ (.A0(_02349_),
    .A1(\fifo_bank_register.data_out[44] ),
    .S(_02290_),
    .X(_02350_));
 sky130_fd_sc_hd__clkbuf_1 _13959_ (.A(_02350_),
    .X(_01485_));
 sky130_fd_sc_hd__a22o_1 _13960_ (.A1(\fifo_bank_register.bank[5][45] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][45] ),
    .X(_02351_));
 sky130_fd_sc_hd__a221o_1 _13961_ (.A1(\fifo_bank_register.bank[7][45] ),
    .A2(_02299_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][45] ),
    .C1(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__a22o_1 _13962_ (.A1(\fifo_bank_register.bank[6][45] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][45] ),
    .X(_02353_));
 sky130_fd_sc_hd__a22o_1 _13963_ (.A1(\fifo_bank_register.bank[1][45] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][45] ),
    .X(_02354_));
 sky130_fd_sc_hd__a2111o_1 _13964_ (.A1(\fifo_bank_register.bank[9][45] ),
    .A2(_02307_),
    .B1(_02352_),
    .C1(_02353_),
    .D1(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__mux2_1 _13965_ (.A0(\fifo_bank_register.bank[0][45] ),
    .A1(_02355_),
    .S(_02320_),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _13966_ (.A0(_02356_),
    .A1(\fifo_bank_register.data_out[45] ),
    .S(_02290_),
    .X(_02357_));
 sky130_fd_sc_hd__clkbuf_1 _13967_ (.A(_02357_),
    .X(_01486_));
 sky130_fd_sc_hd__a22o_1 _13968_ (.A1(\fifo_bank_register.bank[5][46] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][46] ),
    .X(_02358_));
 sky130_fd_sc_hd__a221o_1 _13969_ (.A1(\fifo_bank_register.bank[7][46] ),
    .A2(_02299_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][46] ),
    .C1(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__a22o_1 _13970_ (.A1(\fifo_bank_register.bank[6][46] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][46] ),
    .X(_02360_));
 sky130_fd_sc_hd__a22o_1 _13971_ (.A1(\fifo_bank_register.bank[1][46] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][46] ),
    .X(_02361_));
 sky130_fd_sc_hd__a2111o_1 _13972_ (.A1(\fifo_bank_register.bank[9][46] ),
    .A2(_02307_),
    .B1(_02359_),
    .C1(_02360_),
    .D1(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _13973_ (.A0(\fifo_bank_register.bank[0][46] ),
    .A1(_02362_),
    .S(_02320_),
    .X(_02363_));
 sky130_fd_sc_hd__mux2_1 _13974_ (.A0(_02363_),
    .A1(\fifo_bank_register.data_out[46] ),
    .S(_02290_),
    .X(_02364_));
 sky130_fd_sc_hd__clkbuf_1 _13975_ (.A(_02364_),
    .X(_01487_));
 sky130_fd_sc_hd__a22o_1 _13976_ (.A1(\fifo_bank_register.bank[5][47] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][47] ),
    .X(_02365_));
 sky130_fd_sc_hd__a221o_1 _13977_ (.A1(\fifo_bank_register.bank[7][47] ),
    .A2(_02299_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][47] ),
    .C1(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__a22o_1 _13978_ (.A1(\fifo_bank_register.bank[6][47] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][47] ),
    .X(_02367_));
 sky130_fd_sc_hd__a22o_1 _13979_ (.A1(\fifo_bank_register.bank[1][47] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][47] ),
    .X(_02368_));
 sky130_fd_sc_hd__a2111o_1 _13980_ (.A1(\fifo_bank_register.bank[9][47] ),
    .A2(_02307_),
    .B1(_02366_),
    .C1(_02367_),
    .D1(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__mux2_1 _13981_ (.A0(\fifo_bank_register.bank[0][47] ),
    .A1(_02369_),
    .S(_02320_),
    .X(_02370_));
 sky130_fd_sc_hd__buf_8 _13982_ (.A(_08068_),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _13983_ (.A0(_02370_),
    .A1(\fifo_bank_register.data_out[47] ),
    .S(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__clkbuf_1 _13984_ (.A(_02372_),
    .X(_01488_));
 sky130_fd_sc_hd__a22o_1 _13985_ (.A1(\fifo_bank_register.bank[5][48] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][48] ),
    .X(_02373_));
 sky130_fd_sc_hd__a221o_1 _13986_ (.A1(\fifo_bank_register.bank[7][48] ),
    .A2(_02299_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][48] ),
    .C1(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__a22o_1 _13987_ (.A1(\fifo_bank_register.bank[6][48] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][48] ),
    .X(_02375_));
 sky130_fd_sc_hd__a22o_1 _13988_ (.A1(\fifo_bank_register.bank[1][48] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][48] ),
    .X(_02376_));
 sky130_fd_sc_hd__a2111o_1 _13989_ (.A1(\fifo_bank_register.bank[9][48] ),
    .A2(_02307_),
    .B1(_02374_),
    .C1(_02375_),
    .D1(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _13990_ (.A0(\fifo_bank_register.bank[0][48] ),
    .A1(_02377_),
    .S(_02320_),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _13991_ (.A0(_02378_),
    .A1(\fifo_bank_register.data_out[48] ),
    .S(_02371_),
    .X(_02379_));
 sky130_fd_sc_hd__clkbuf_1 _13992_ (.A(_02379_),
    .X(_01489_));
 sky130_fd_sc_hd__clkbuf_8 _13993_ (.A(_08181_),
    .X(_02380_));
 sky130_fd_sc_hd__a22o_1 _13994_ (.A1(\fifo_bank_register.bank[5][49] ),
    .A2(_02309_),
    .B1(_02310_),
    .B2(\fifo_bank_register.bank[3][49] ),
    .X(_02381_));
 sky130_fd_sc_hd__a221o_1 _13995_ (.A1(\fifo_bank_register.bank[7][49] ),
    .A2(_02380_),
    .B1(_02308_),
    .B2(\fifo_bank_register.bank[2][49] ),
    .C1(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__a22o_1 _13996_ (.A1(\fifo_bank_register.bank[6][49] ),
    .A2(_02313_),
    .B1(_02314_),
    .B2(\fifo_bank_register.bank[4][49] ),
    .X(_02383_));
 sky130_fd_sc_hd__a22o_1 _13997_ (.A1(\fifo_bank_register.bank[1][49] ),
    .A2(_02316_),
    .B1(_02317_),
    .B2(\fifo_bank_register.bank[8][49] ),
    .X(_02384_));
 sky130_fd_sc_hd__a2111o_1 _13998_ (.A1(\fifo_bank_register.bank[9][49] ),
    .A2(_02307_),
    .B1(_02382_),
    .C1(_02383_),
    .D1(_02384_),
    .X(_02385_));
 sky130_fd_sc_hd__mux2_1 _13999_ (.A0(\fifo_bank_register.bank[0][49] ),
    .A1(_02385_),
    .S(_02320_),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _14000_ (.A0(_02386_),
    .A1(\fifo_bank_register.data_out[49] ),
    .S(_02371_),
    .X(_02387_));
 sky130_fd_sc_hd__clkbuf_1 _14001_ (.A(_02387_),
    .X(_01490_));
 sky130_fd_sc_hd__clkbuf_4 _14002_ (.A(_02136_),
    .X(_02388_));
 sky130_fd_sc_hd__clkbuf_4 _14003_ (.A(_02138_),
    .X(_02389_));
 sky130_fd_sc_hd__clkbuf_4 _14004_ (.A(_02140_),
    .X(_02390_));
 sky130_fd_sc_hd__clkbuf_4 _14005_ (.A(_02142_),
    .X(_02391_));
 sky130_fd_sc_hd__a22o_1 _14006_ (.A1(\fifo_bank_register.bank[5][50] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][50] ),
    .X(_02392_));
 sky130_fd_sc_hd__a221o_1 _14007_ (.A1(\fifo_bank_register.bank[7][50] ),
    .A2(_02380_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][50] ),
    .C1(_02392_),
    .X(_02393_));
 sky130_fd_sc_hd__buf_4 _14008_ (.A(_02146_),
    .X(_02394_));
 sky130_fd_sc_hd__buf_4 _14009_ (.A(_02148_),
    .X(_02395_));
 sky130_fd_sc_hd__a22o_1 _14010_ (.A1(\fifo_bank_register.bank[6][50] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][50] ),
    .X(_02396_));
 sky130_fd_sc_hd__clkbuf_4 _14011_ (.A(_02151_),
    .X(_02397_));
 sky130_fd_sc_hd__clkbuf_4 _14012_ (.A(_02153_),
    .X(_02398_));
 sky130_fd_sc_hd__a22o_1 _14013_ (.A1(\fifo_bank_register.bank[1][50] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][50] ),
    .X(_02399_));
 sky130_fd_sc_hd__a2111o_1 _14014_ (.A1(\fifo_bank_register.bank[9][50] ),
    .A2(_02388_),
    .B1(_02393_),
    .C1(_02396_),
    .D1(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__buf_4 _14015_ (.A(_02157_),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _14016_ (.A0(\fifo_bank_register.bank[0][50] ),
    .A1(_02400_),
    .S(_02401_),
    .X(_02402_));
 sky130_fd_sc_hd__mux2_1 _14017_ (.A0(_02402_),
    .A1(\fifo_bank_register.data_out[50] ),
    .S(_02371_),
    .X(_02403_));
 sky130_fd_sc_hd__clkbuf_1 _14018_ (.A(_02403_),
    .X(_01491_));
 sky130_fd_sc_hd__a22o_1 _14019_ (.A1(\fifo_bank_register.bank[5][51] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][51] ),
    .X(_02404_));
 sky130_fd_sc_hd__a221o_1 _14020_ (.A1(\fifo_bank_register.bank[7][51] ),
    .A2(_02380_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][51] ),
    .C1(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__a22o_1 _14021_ (.A1(\fifo_bank_register.bank[6][51] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][51] ),
    .X(_02406_));
 sky130_fd_sc_hd__a22o_1 _14022_ (.A1(\fifo_bank_register.bank[1][51] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][51] ),
    .X(_02407_));
 sky130_fd_sc_hd__a2111o_1 _14023_ (.A1(\fifo_bank_register.bank[9][51] ),
    .A2(_02388_),
    .B1(_02405_),
    .C1(_02406_),
    .D1(_02407_),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _14024_ (.A0(\fifo_bank_register.bank[0][51] ),
    .A1(_02408_),
    .S(_02401_),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _14025_ (.A0(_02409_),
    .A1(\fifo_bank_register.data_out[51] ),
    .S(_02371_),
    .X(_02410_));
 sky130_fd_sc_hd__clkbuf_1 _14026_ (.A(_02410_),
    .X(_01492_));
 sky130_fd_sc_hd__a22o_1 _14027_ (.A1(\fifo_bank_register.bank[5][52] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][52] ),
    .X(_02411_));
 sky130_fd_sc_hd__a221o_1 _14028_ (.A1(\fifo_bank_register.bank[7][52] ),
    .A2(_02380_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][52] ),
    .C1(_02411_),
    .X(_02412_));
 sky130_fd_sc_hd__a22o_1 _14029_ (.A1(\fifo_bank_register.bank[6][52] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][52] ),
    .X(_02413_));
 sky130_fd_sc_hd__a22o_1 _14030_ (.A1(\fifo_bank_register.bank[1][52] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][52] ),
    .X(_02414_));
 sky130_fd_sc_hd__a2111o_1 _14031_ (.A1(\fifo_bank_register.bank[9][52] ),
    .A2(_02388_),
    .B1(_02412_),
    .C1(_02413_),
    .D1(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _14032_ (.A0(\fifo_bank_register.bank[0][52] ),
    .A1(_02415_),
    .S(_02401_),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _14033_ (.A0(_02416_),
    .A1(\fifo_bank_register.data_out[52] ),
    .S(_02371_),
    .X(_02417_));
 sky130_fd_sc_hd__clkbuf_1 _14034_ (.A(_02417_),
    .X(_01493_));
 sky130_fd_sc_hd__a22o_1 _14035_ (.A1(\fifo_bank_register.bank[5][53] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][53] ),
    .X(_02418_));
 sky130_fd_sc_hd__a221o_1 _14036_ (.A1(\fifo_bank_register.bank[7][53] ),
    .A2(_02380_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][53] ),
    .C1(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__a22o_1 _14037_ (.A1(\fifo_bank_register.bank[6][53] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][53] ),
    .X(_02420_));
 sky130_fd_sc_hd__a22o_1 _14038_ (.A1(\fifo_bank_register.bank[1][53] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][53] ),
    .X(_02421_));
 sky130_fd_sc_hd__a2111o_1 _14039_ (.A1(\fifo_bank_register.bank[9][53] ),
    .A2(_02388_),
    .B1(_02419_),
    .C1(_02420_),
    .D1(_02421_),
    .X(_02422_));
 sky130_fd_sc_hd__mux2_1 _14040_ (.A0(\fifo_bank_register.bank[0][53] ),
    .A1(_02422_),
    .S(_02401_),
    .X(_02423_));
 sky130_fd_sc_hd__mux2_1 _14041_ (.A0(_02423_),
    .A1(\fifo_bank_register.data_out[53] ),
    .S(_02371_),
    .X(_02424_));
 sky130_fd_sc_hd__clkbuf_1 _14042_ (.A(_02424_),
    .X(_01494_));
 sky130_fd_sc_hd__a22o_1 _14043_ (.A1(\fifo_bank_register.bank[5][54] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][54] ),
    .X(_02425_));
 sky130_fd_sc_hd__a221o_1 _14044_ (.A1(\fifo_bank_register.bank[7][54] ),
    .A2(_02380_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][54] ),
    .C1(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__a22o_1 _14045_ (.A1(\fifo_bank_register.bank[6][54] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][54] ),
    .X(_02427_));
 sky130_fd_sc_hd__a22o_1 _14046_ (.A1(\fifo_bank_register.bank[1][54] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][54] ),
    .X(_02428_));
 sky130_fd_sc_hd__a2111o_1 _14047_ (.A1(\fifo_bank_register.bank[9][54] ),
    .A2(_02388_),
    .B1(_02426_),
    .C1(_02427_),
    .D1(_02428_),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _14048_ (.A0(\fifo_bank_register.bank[0][54] ),
    .A1(_02429_),
    .S(_02401_),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _14049_ (.A0(_02430_),
    .A1(\fifo_bank_register.data_out[54] ),
    .S(_02371_),
    .X(_02431_));
 sky130_fd_sc_hd__clkbuf_1 _14050_ (.A(_02431_),
    .X(_01495_));
 sky130_fd_sc_hd__a22o_1 _14051_ (.A1(\fifo_bank_register.bank[5][55] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][55] ),
    .X(_02432_));
 sky130_fd_sc_hd__a221o_1 _14052_ (.A1(\fifo_bank_register.bank[7][55] ),
    .A2(_02380_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][55] ),
    .C1(_02432_),
    .X(_02433_));
 sky130_fd_sc_hd__a22o_1 _14053_ (.A1(\fifo_bank_register.bank[6][55] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][55] ),
    .X(_02434_));
 sky130_fd_sc_hd__a22o_1 _14054_ (.A1(\fifo_bank_register.bank[1][55] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][55] ),
    .X(_02435_));
 sky130_fd_sc_hd__a2111o_1 _14055_ (.A1(\fifo_bank_register.bank[9][55] ),
    .A2(_02388_),
    .B1(_02433_),
    .C1(_02434_),
    .D1(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__mux2_1 _14056_ (.A0(\fifo_bank_register.bank[0][55] ),
    .A1(_02436_),
    .S(_02401_),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _14057_ (.A0(_02437_),
    .A1(\fifo_bank_register.data_out[55] ),
    .S(_02371_),
    .X(_02438_));
 sky130_fd_sc_hd__clkbuf_1 _14058_ (.A(_02438_),
    .X(_01496_));
 sky130_fd_sc_hd__a22o_1 _14059_ (.A1(\fifo_bank_register.bank[5][56] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][56] ),
    .X(_02439_));
 sky130_fd_sc_hd__a221o_1 _14060_ (.A1(\fifo_bank_register.bank[7][56] ),
    .A2(_02380_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][56] ),
    .C1(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__a22o_1 _14061_ (.A1(\fifo_bank_register.bank[6][56] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][56] ),
    .X(_02441_));
 sky130_fd_sc_hd__a22o_1 _14062_ (.A1(\fifo_bank_register.bank[1][56] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][56] ),
    .X(_02442_));
 sky130_fd_sc_hd__a2111o_1 _14063_ (.A1(\fifo_bank_register.bank[9][56] ),
    .A2(_02388_),
    .B1(_02440_),
    .C1(_02441_),
    .D1(_02442_),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _14064_ (.A0(\fifo_bank_register.bank[0][56] ),
    .A1(_02443_),
    .S(_02401_),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _14065_ (.A0(_02444_),
    .A1(\fifo_bank_register.data_out[56] ),
    .S(_02371_),
    .X(_02445_));
 sky130_fd_sc_hd__clkbuf_1 _14066_ (.A(_02445_),
    .X(_01497_));
 sky130_fd_sc_hd__a22o_1 _14067_ (.A1(\fifo_bank_register.bank[5][57] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][57] ),
    .X(_02446_));
 sky130_fd_sc_hd__a221o_1 _14068_ (.A1(\fifo_bank_register.bank[7][57] ),
    .A2(_02380_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][57] ),
    .C1(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__a22o_1 _14069_ (.A1(\fifo_bank_register.bank[6][57] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][57] ),
    .X(_02448_));
 sky130_fd_sc_hd__a22o_1 _14070_ (.A1(\fifo_bank_register.bank[1][57] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][57] ),
    .X(_02449_));
 sky130_fd_sc_hd__a2111o_1 _14071_ (.A1(\fifo_bank_register.bank[9][57] ),
    .A2(_02388_),
    .B1(_02447_),
    .C1(_02448_),
    .D1(_02449_),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _14072_ (.A0(\fifo_bank_register.bank[0][57] ),
    .A1(_02450_),
    .S(_02401_),
    .X(_02451_));
 sky130_fd_sc_hd__clkbuf_8 _14073_ (.A(_08068_),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _14074_ (.A0(_02451_),
    .A1(\fifo_bank_register.data_out[57] ),
    .S(_02452_),
    .X(_02453_));
 sky130_fd_sc_hd__clkbuf_1 _14075_ (.A(_02453_),
    .X(_01498_));
 sky130_fd_sc_hd__a22o_1 _14076_ (.A1(\fifo_bank_register.bank[5][58] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][58] ),
    .X(_02454_));
 sky130_fd_sc_hd__a221o_1 _14077_ (.A1(\fifo_bank_register.bank[7][58] ),
    .A2(_02380_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][58] ),
    .C1(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__a22o_1 _14078_ (.A1(\fifo_bank_register.bank[6][58] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][58] ),
    .X(_02456_));
 sky130_fd_sc_hd__a22o_1 _14079_ (.A1(\fifo_bank_register.bank[1][58] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][58] ),
    .X(_02457_));
 sky130_fd_sc_hd__a2111o_1 _14080_ (.A1(\fifo_bank_register.bank[9][58] ),
    .A2(_02388_),
    .B1(_02455_),
    .C1(_02456_),
    .D1(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _14081_ (.A0(\fifo_bank_register.bank[0][58] ),
    .A1(_02458_),
    .S(_02401_),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _14082_ (.A0(_02459_),
    .A1(\fifo_bank_register.data_out[58] ),
    .S(_02452_),
    .X(_02460_));
 sky130_fd_sc_hd__clkbuf_1 _14083_ (.A(_02460_),
    .X(_01499_));
 sky130_fd_sc_hd__buf_4 _14084_ (.A(_08181_),
    .X(_02461_));
 sky130_fd_sc_hd__a22o_1 _14085_ (.A1(\fifo_bank_register.bank[5][59] ),
    .A2(_02390_),
    .B1(_02391_),
    .B2(\fifo_bank_register.bank[3][59] ),
    .X(_02462_));
 sky130_fd_sc_hd__a221o_1 _14086_ (.A1(\fifo_bank_register.bank[7][59] ),
    .A2(_02461_),
    .B1(_02389_),
    .B2(\fifo_bank_register.bank[2][59] ),
    .C1(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__a22o_1 _14087_ (.A1(\fifo_bank_register.bank[6][59] ),
    .A2(_02394_),
    .B1(_02395_),
    .B2(\fifo_bank_register.bank[4][59] ),
    .X(_02464_));
 sky130_fd_sc_hd__a22o_1 _14088_ (.A1(\fifo_bank_register.bank[1][59] ),
    .A2(_02397_),
    .B1(_02398_),
    .B2(\fifo_bank_register.bank[8][59] ),
    .X(_02465_));
 sky130_fd_sc_hd__a2111o_1 _14089_ (.A1(\fifo_bank_register.bank[9][59] ),
    .A2(_02388_),
    .B1(_02463_),
    .C1(_02464_),
    .D1(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _14090_ (.A0(\fifo_bank_register.bank[0][59] ),
    .A1(_02466_),
    .S(_02401_),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _14091_ (.A0(_02467_),
    .A1(\fifo_bank_register.data_out[59] ),
    .S(_02452_),
    .X(_02468_));
 sky130_fd_sc_hd__clkbuf_1 _14092_ (.A(_02468_),
    .X(_01500_));
 sky130_fd_sc_hd__clkbuf_4 _14093_ (.A(_02136_),
    .X(_02469_));
 sky130_fd_sc_hd__clkbuf_4 _14094_ (.A(_02138_),
    .X(_02470_));
 sky130_fd_sc_hd__clkbuf_4 _14095_ (.A(_02140_),
    .X(_02471_));
 sky130_fd_sc_hd__clkbuf_4 _14096_ (.A(_02142_),
    .X(_02472_));
 sky130_fd_sc_hd__a22o_1 _14097_ (.A1(\fifo_bank_register.bank[5][60] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][60] ),
    .X(_02473_));
 sky130_fd_sc_hd__a221o_1 _14098_ (.A1(\fifo_bank_register.bank[7][60] ),
    .A2(_02461_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][60] ),
    .C1(_02473_),
    .X(_02474_));
 sky130_fd_sc_hd__clkbuf_4 _14099_ (.A(_02146_),
    .X(_02475_));
 sky130_fd_sc_hd__clkbuf_4 _14100_ (.A(_02148_),
    .X(_02476_));
 sky130_fd_sc_hd__a22o_1 _14101_ (.A1(\fifo_bank_register.bank[6][60] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][60] ),
    .X(_02477_));
 sky130_fd_sc_hd__buf_4 _14102_ (.A(_02151_),
    .X(_02478_));
 sky130_fd_sc_hd__buf_4 _14103_ (.A(_02153_),
    .X(_02479_));
 sky130_fd_sc_hd__a22o_1 _14104_ (.A1(\fifo_bank_register.bank[1][60] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][60] ),
    .X(_02480_));
 sky130_fd_sc_hd__a2111o_1 _14105_ (.A1(\fifo_bank_register.bank[9][60] ),
    .A2(_02469_),
    .B1(_02474_),
    .C1(_02477_),
    .D1(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__buf_4 _14106_ (.A(_02157_),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _14107_ (.A0(\fifo_bank_register.bank[0][60] ),
    .A1(_02481_),
    .S(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _14108_ (.A0(_02483_),
    .A1(\fifo_bank_register.data_out[60] ),
    .S(_02452_),
    .X(_02484_));
 sky130_fd_sc_hd__clkbuf_1 _14109_ (.A(_02484_),
    .X(_01501_));
 sky130_fd_sc_hd__a22o_1 _14110_ (.A1(\fifo_bank_register.bank[5][61] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][61] ),
    .X(_02485_));
 sky130_fd_sc_hd__a221o_1 _14111_ (.A1(\fifo_bank_register.bank[7][61] ),
    .A2(_02461_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][61] ),
    .C1(_02485_),
    .X(_02486_));
 sky130_fd_sc_hd__a22o_1 _14112_ (.A1(\fifo_bank_register.bank[6][61] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][61] ),
    .X(_02487_));
 sky130_fd_sc_hd__a22o_1 _14113_ (.A1(\fifo_bank_register.bank[1][61] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][61] ),
    .X(_02488_));
 sky130_fd_sc_hd__a2111o_1 _14114_ (.A1(\fifo_bank_register.bank[9][61] ),
    .A2(_02469_),
    .B1(_02486_),
    .C1(_02487_),
    .D1(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _14115_ (.A0(\fifo_bank_register.bank[0][61] ),
    .A1(_02489_),
    .S(_02482_),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _14116_ (.A0(_02490_),
    .A1(\fifo_bank_register.data_out[61] ),
    .S(_02452_),
    .X(_02491_));
 sky130_fd_sc_hd__clkbuf_1 _14117_ (.A(_02491_),
    .X(_01502_));
 sky130_fd_sc_hd__a22o_1 _14118_ (.A1(\fifo_bank_register.bank[5][62] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][62] ),
    .X(_02492_));
 sky130_fd_sc_hd__a221o_1 _14119_ (.A1(\fifo_bank_register.bank[7][62] ),
    .A2(_02461_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][62] ),
    .C1(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__a22o_1 _14120_ (.A1(\fifo_bank_register.bank[6][62] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][62] ),
    .X(_02494_));
 sky130_fd_sc_hd__a22o_1 _14121_ (.A1(\fifo_bank_register.bank[1][62] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][62] ),
    .X(_02495_));
 sky130_fd_sc_hd__a2111o_1 _14122_ (.A1(\fifo_bank_register.bank[9][62] ),
    .A2(_02469_),
    .B1(_02493_),
    .C1(_02494_),
    .D1(_02495_),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _14123_ (.A0(\fifo_bank_register.bank[0][62] ),
    .A1(_02496_),
    .S(_02482_),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _14124_ (.A0(_02497_),
    .A1(\fifo_bank_register.data_out[62] ),
    .S(_02452_),
    .X(_02498_));
 sky130_fd_sc_hd__clkbuf_1 _14125_ (.A(_02498_),
    .X(_01503_));
 sky130_fd_sc_hd__a22o_1 _14126_ (.A1(\fifo_bank_register.bank[5][63] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][63] ),
    .X(_02499_));
 sky130_fd_sc_hd__a221o_1 _14127_ (.A1(\fifo_bank_register.bank[7][63] ),
    .A2(_02461_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][63] ),
    .C1(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__a22o_1 _14128_ (.A1(\fifo_bank_register.bank[6][63] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][63] ),
    .X(_02501_));
 sky130_fd_sc_hd__a22o_1 _14129_ (.A1(\fifo_bank_register.bank[1][63] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][63] ),
    .X(_02502_));
 sky130_fd_sc_hd__a2111o_1 _14130_ (.A1(\fifo_bank_register.bank[9][63] ),
    .A2(_02469_),
    .B1(_02500_),
    .C1(_02501_),
    .D1(_02502_),
    .X(_02503_));
 sky130_fd_sc_hd__mux2_2 _14131_ (.A0(\fifo_bank_register.bank[0][63] ),
    .A1(_02503_),
    .S(_02482_),
    .X(_02504_));
 sky130_fd_sc_hd__mux2_1 _14132_ (.A0(_02504_),
    .A1(\fifo_bank_register.data_out[63] ),
    .S(_02452_),
    .X(_02505_));
 sky130_fd_sc_hd__clkbuf_1 _14133_ (.A(_02505_),
    .X(_01504_));
 sky130_fd_sc_hd__a22o_1 _14134_ (.A1(\fifo_bank_register.bank[5][64] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][64] ),
    .X(_02506_));
 sky130_fd_sc_hd__a221o_1 _14135_ (.A1(\fifo_bank_register.bank[7][64] ),
    .A2(_02461_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][64] ),
    .C1(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__a22o_1 _14136_ (.A1(\fifo_bank_register.bank[6][64] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][64] ),
    .X(_02508_));
 sky130_fd_sc_hd__a22o_1 _14137_ (.A1(\fifo_bank_register.bank[1][64] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][64] ),
    .X(_02509_));
 sky130_fd_sc_hd__a2111o_1 _14138_ (.A1(\fifo_bank_register.bank[9][64] ),
    .A2(_02469_),
    .B1(_02507_),
    .C1(_02508_),
    .D1(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _14139_ (.A0(\fifo_bank_register.bank[0][64] ),
    .A1(_02510_),
    .S(_02482_),
    .X(_02511_));
 sky130_fd_sc_hd__mux2_1 _14140_ (.A0(_02511_),
    .A1(\fifo_bank_register.data_out[64] ),
    .S(_02452_),
    .X(_02512_));
 sky130_fd_sc_hd__clkbuf_1 _14141_ (.A(_02512_),
    .X(_01505_));
 sky130_fd_sc_hd__a22o_1 _14142_ (.A1(\fifo_bank_register.bank[5][65] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][65] ),
    .X(_02513_));
 sky130_fd_sc_hd__a221o_1 _14143_ (.A1(\fifo_bank_register.bank[7][65] ),
    .A2(_02461_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][65] ),
    .C1(_02513_),
    .X(_02514_));
 sky130_fd_sc_hd__a22o_1 _14144_ (.A1(\fifo_bank_register.bank[6][65] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][65] ),
    .X(_02515_));
 sky130_fd_sc_hd__a22o_1 _14145_ (.A1(\fifo_bank_register.bank[1][65] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][65] ),
    .X(_02516_));
 sky130_fd_sc_hd__a2111o_1 _14146_ (.A1(\fifo_bank_register.bank[9][65] ),
    .A2(_02469_),
    .B1(_02514_),
    .C1(_02515_),
    .D1(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__mux2_1 _14147_ (.A0(\fifo_bank_register.bank[0][65] ),
    .A1(_02517_),
    .S(_02482_),
    .X(_02518_));
 sky130_fd_sc_hd__mux2_1 _14148_ (.A0(_02518_),
    .A1(\fifo_bank_register.data_out[65] ),
    .S(_02452_),
    .X(_02519_));
 sky130_fd_sc_hd__clkbuf_1 _14149_ (.A(_02519_),
    .X(_01506_));
 sky130_fd_sc_hd__a22o_1 _14150_ (.A1(\fifo_bank_register.bank[5][66] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][66] ),
    .X(_02520_));
 sky130_fd_sc_hd__a221o_1 _14151_ (.A1(\fifo_bank_register.bank[7][66] ),
    .A2(_02461_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][66] ),
    .C1(_02520_),
    .X(_02521_));
 sky130_fd_sc_hd__a22o_1 _14152_ (.A1(\fifo_bank_register.bank[6][66] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][66] ),
    .X(_02522_));
 sky130_fd_sc_hd__a22o_1 _14153_ (.A1(\fifo_bank_register.bank[1][66] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][66] ),
    .X(_02523_));
 sky130_fd_sc_hd__a2111o_1 _14154_ (.A1(\fifo_bank_register.bank[9][66] ),
    .A2(_02469_),
    .B1(_02521_),
    .C1(_02522_),
    .D1(_02523_),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _14155_ (.A0(\fifo_bank_register.bank[0][66] ),
    .A1(_02524_),
    .S(_02482_),
    .X(_02525_));
 sky130_fd_sc_hd__mux2_1 _14156_ (.A0(_02525_),
    .A1(\fifo_bank_register.data_out[66] ),
    .S(_02452_),
    .X(_02526_));
 sky130_fd_sc_hd__clkbuf_1 _14157_ (.A(_02526_),
    .X(_01507_));
 sky130_fd_sc_hd__a22o_1 _14158_ (.A1(\fifo_bank_register.bank[5][67] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][67] ),
    .X(_02527_));
 sky130_fd_sc_hd__a221o_1 _14159_ (.A1(\fifo_bank_register.bank[7][67] ),
    .A2(_02461_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][67] ),
    .C1(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__a22o_1 _14160_ (.A1(\fifo_bank_register.bank[6][67] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][67] ),
    .X(_02529_));
 sky130_fd_sc_hd__a22o_1 _14161_ (.A1(\fifo_bank_register.bank[1][67] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][67] ),
    .X(_02530_));
 sky130_fd_sc_hd__a2111o_1 _14162_ (.A1(\fifo_bank_register.bank[9][67] ),
    .A2(_02469_),
    .B1(_02528_),
    .C1(_02529_),
    .D1(_02530_),
    .X(_02531_));
 sky130_fd_sc_hd__mux2_1 _14163_ (.A0(\fifo_bank_register.bank[0][67] ),
    .A1(_02531_),
    .S(_02482_),
    .X(_02532_));
 sky130_fd_sc_hd__clkbuf_8 _14164_ (.A(_08068_),
    .X(_02533_));
 sky130_fd_sc_hd__mux2_1 _14165_ (.A0(_02532_),
    .A1(\fifo_bank_register.data_out[67] ),
    .S(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__clkbuf_1 _14166_ (.A(_02534_),
    .X(_01508_));
 sky130_fd_sc_hd__a22o_1 _14167_ (.A1(\fifo_bank_register.bank[5][68] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][68] ),
    .X(_02535_));
 sky130_fd_sc_hd__a221o_1 _14168_ (.A1(\fifo_bank_register.bank[7][68] ),
    .A2(_02461_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][68] ),
    .C1(_02535_),
    .X(_02536_));
 sky130_fd_sc_hd__a22o_1 _14169_ (.A1(\fifo_bank_register.bank[6][68] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][68] ),
    .X(_02537_));
 sky130_fd_sc_hd__a22o_1 _14170_ (.A1(\fifo_bank_register.bank[1][68] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][68] ),
    .X(_02538_));
 sky130_fd_sc_hd__a2111o_1 _14171_ (.A1(\fifo_bank_register.bank[9][68] ),
    .A2(_02469_),
    .B1(_02536_),
    .C1(_02537_),
    .D1(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__mux2_1 _14172_ (.A0(\fifo_bank_register.bank[0][68] ),
    .A1(_02539_),
    .S(_02482_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _14173_ (.A0(_02540_),
    .A1(\fifo_bank_register.data_out[68] ),
    .S(_02533_),
    .X(_02541_));
 sky130_fd_sc_hd__clkbuf_1 _14174_ (.A(_02541_),
    .X(_01509_));
 sky130_fd_sc_hd__clkbuf_4 _14175_ (.A(_08181_),
    .X(_02542_));
 sky130_fd_sc_hd__a22o_1 _14176_ (.A1(\fifo_bank_register.bank[5][69] ),
    .A2(_02471_),
    .B1(_02472_),
    .B2(\fifo_bank_register.bank[3][69] ),
    .X(_02543_));
 sky130_fd_sc_hd__a221o_1 _14177_ (.A1(\fifo_bank_register.bank[7][69] ),
    .A2(_02542_),
    .B1(_02470_),
    .B2(\fifo_bank_register.bank[2][69] ),
    .C1(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__a22o_1 _14178_ (.A1(\fifo_bank_register.bank[6][69] ),
    .A2(_02475_),
    .B1(_02476_),
    .B2(\fifo_bank_register.bank[4][69] ),
    .X(_02545_));
 sky130_fd_sc_hd__a22o_1 _14179_ (.A1(\fifo_bank_register.bank[1][69] ),
    .A2(_02478_),
    .B1(_02479_),
    .B2(\fifo_bank_register.bank[8][69] ),
    .X(_02546_));
 sky130_fd_sc_hd__a2111o_1 _14180_ (.A1(\fifo_bank_register.bank[9][69] ),
    .A2(_02469_),
    .B1(_02544_),
    .C1(_02545_),
    .D1(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__mux2_1 _14181_ (.A0(\fifo_bank_register.bank[0][69] ),
    .A1(_02547_),
    .S(_02482_),
    .X(_02548_));
 sky130_fd_sc_hd__mux2_1 _14182_ (.A0(_02548_),
    .A1(\fifo_bank_register.data_out[69] ),
    .S(_02533_),
    .X(_02549_));
 sky130_fd_sc_hd__clkbuf_1 _14183_ (.A(_02549_),
    .X(_01510_));
 sky130_fd_sc_hd__clkbuf_4 _14184_ (.A(_02136_),
    .X(_02550_));
 sky130_fd_sc_hd__clkbuf_4 _14185_ (.A(_02138_),
    .X(_02551_));
 sky130_fd_sc_hd__clkbuf_4 _14186_ (.A(_02140_),
    .X(_02552_));
 sky130_fd_sc_hd__clkbuf_4 _14187_ (.A(_02142_),
    .X(_02553_));
 sky130_fd_sc_hd__a22o_1 _14188_ (.A1(\fifo_bank_register.bank[5][70] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][70] ),
    .X(_02554_));
 sky130_fd_sc_hd__a221o_1 _14189_ (.A1(\fifo_bank_register.bank[7][70] ),
    .A2(_02542_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][70] ),
    .C1(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__clkbuf_4 _14190_ (.A(_02146_),
    .X(_02556_));
 sky130_fd_sc_hd__clkbuf_4 _14191_ (.A(_02148_),
    .X(_02557_));
 sky130_fd_sc_hd__a22o_1 _14192_ (.A1(\fifo_bank_register.bank[6][70] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][70] ),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_4 _14193_ (.A(_02151_),
    .X(_02559_));
 sky130_fd_sc_hd__clkbuf_4 _14194_ (.A(_02153_),
    .X(_02560_));
 sky130_fd_sc_hd__a22o_1 _14195_ (.A1(\fifo_bank_register.bank[1][70] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][70] ),
    .X(_02561_));
 sky130_fd_sc_hd__a2111o_1 _14196_ (.A1(\fifo_bank_register.bank[9][70] ),
    .A2(_02550_),
    .B1(_02555_),
    .C1(_02558_),
    .D1(_02561_),
    .X(_02562_));
 sky130_fd_sc_hd__buf_4 _14197_ (.A(_02157_),
    .X(_02563_));
 sky130_fd_sc_hd__mux2_1 _14198_ (.A0(\fifo_bank_register.bank[0][70] ),
    .A1(_02562_),
    .S(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_1 _14199_ (.A0(_02564_),
    .A1(\fifo_bank_register.data_out[70] ),
    .S(_02533_),
    .X(_02565_));
 sky130_fd_sc_hd__clkbuf_1 _14200_ (.A(_02565_),
    .X(_01511_));
 sky130_fd_sc_hd__a22o_1 _14201_ (.A1(\fifo_bank_register.bank[5][71] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][71] ),
    .X(_02566_));
 sky130_fd_sc_hd__a221o_1 _14202_ (.A1(\fifo_bank_register.bank[7][71] ),
    .A2(_02542_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][71] ),
    .C1(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__a22o_1 _14203_ (.A1(\fifo_bank_register.bank[6][71] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][71] ),
    .X(_02568_));
 sky130_fd_sc_hd__a22o_1 _14204_ (.A1(\fifo_bank_register.bank[1][71] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][71] ),
    .X(_02569_));
 sky130_fd_sc_hd__a2111o_1 _14205_ (.A1(\fifo_bank_register.bank[9][71] ),
    .A2(_02550_),
    .B1(_02567_),
    .C1(_02568_),
    .D1(_02569_),
    .X(_02570_));
 sky130_fd_sc_hd__mux2_1 _14206_ (.A0(\fifo_bank_register.bank[0][71] ),
    .A1(_02570_),
    .S(_02563_),
    .X(_02571_));
 sky130_fd_sc_hd__mux2_1 _14207_ (.A0(_02571_),
    .A1(\fifo_bank_register.data_out[71] ),
    .S(_02533_),
    .X(_02572_));
 sky130_fd_sc_hd__clkbuf_1 _14208_ (.A(_02572_),
    .X(_01512_));
 sky130_fd_sc_hd__a22o_1 _14209_ (.A1(\fifo_bank_register.bank[5][72] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][72] ),
    .X(_02573_));
 sky130_fd_sc_hd__a221o_1 _14210_ (.A1(\fifo_bank_register.bank[7][72] ),
    .A2(_02542_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][72] ),
    .C1(_02573_),
    .X(_02574_));
 sky130_fd_sc_hd__a22o_1 _14211_ (.A1(\fifo_bank_register.bank[6][72] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][72] ),
    .X(_02575_));
 sky130_fd_sc_hd__a22o_1 _14212_ (.A1(\fifo_bank_register.bank[1][72] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][72] ),
    .X(_02576_));
 sky130_fd_sc_hd__a2111o_1 _14213_ (.A1(\fifo_bank_register.bank[9][72] ),
    .A2(_02550_),
    .B1(_02574_),
    .C1(_02575_),
    .D1(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__mux2_1 _14214_ (.A0(\fifo_bank_register.bank[0][72] ),
    .A1(_02577_),
    .S(_02563_),
    .X(_02578_));
 sky130_fd_sc_hd__mux2_1 _14215_ (.A0(_02578_),
    .A1(\fifo_bank_register.data_out[72] ),
    .S(_02533_),
    .X(_02579_));
 sky130_fd_sc_hd__clkbuf_1 _14216_ (.A(_02579_),
    .X(_01513_));
 sky130_fd_sc_hd__a22o_1 _14217_ (.A1(\fifo_bank_register.bank[5][73] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][73] ),
    .X(_02580_));
 sky130_fd_sc_hd__a221o_1 _14218_ (.A1(\fifo_bank_register.bank[7][73] ),
    .A2(_02542_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][73] ),
    .C1(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__a22o_1 _14219_ (.A1(\fifo_bank_register.bank[6][73] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][73] ),
    .X(_02582_));
 sky130_fd_sc_hd__a22o_1 _14220_ (.A1(\fifo_bank_register.bank[1][73] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][73] ),
    .X(_02583_));
 sky130_fd_sc_hd__a2111o_1 _14221_ (.A1(\fifo_bank_register.bank[9][73] ),
    .A2(_02550_),
    .B1(_02581_),
    .C1(_02582_),
    .D1(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _14222_ (.A0(\fifo_bank_register.bank[0][73] ),
    .A1(_02584_),
    .S(_02563_),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _14223_ (.A0(_02585_),
    .A1(\fifo_bank_register.data_out[73] ),
    .S(_02533_),
    .X(_02586_));
 sky130_fd_sc_hd__clkbuf_1 _14224_ (.A(_02586_),
    .X(_01514_));
 sky130_fd_sc_hd__a22o_1 _14225_ (.A1(\fifo_bank_register.bank[5][74] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][74] ),
    .X(_02587_));
 sky130_fd_sc_hd__a221o_1 _14226_ (.A1(\fifo_bank_register.bank[7][74] ),
    .A2(_02542_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][74] ),
    .C1(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__a22o_1 _14227_ (.A1(\fifo_bank_register.bank[6][74] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][74] ),
    .X(_02589_));
 sky130_fd_sc_hd__a22o_1 _14228_ (.A1(\fifo_bank_register.bank[1][74] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][74] ),
    .X(_02590_));
 sky130_fd_sc_hd__a2111o_1 _14229_ (.A1(\fifo_bank_register.bank[9][74] ),
    .A2(_02550_),
    .B1(_02588_),
    .C1(_02589_),
    .D1(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__mux2_1 _14230_ (.A0(\fifo_bank_register.bank[0][74] ),
    .A1(_02591_),
    .S(_02563_),
    .X(_02592_));
 sky130_fd_sc_hd__mux2_1 _14231_ (.A0(_02592_),
    .A1(\fifo_bank_register.data_out[74] ),
    .S(_02533_),
    .X(_02593_));
 sky130_fd_sc_hd__clkbuf_1 _14232_ (.A(_02593_),
    .X(_01515_));
 sky130_fd_sc_hd__a22o_1 _14233_ (.A1(\fifo_bank_register.bank[5][75] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][75] ),
    .X(_02594_));
 sky130_fd_sc_hd__a221o_1 _14234_ (.A1(\fifo_bank_register.bank[7][75] ),
    .A2(_02542_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][75] ),
    .C1(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__a22o_1 _14235_ (.A1(\fifo_bank_register.bank[6][75] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][75] ),
    .X(_02596_));
 sky130_fd_sc_hd__a22o_1 _14236_ (.A1(\fifo_bank_register.bank[1][75] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][75] ),
    .X(_02597_));
 sky130_fd_sc_hd__a2111o_1 _14237_ (.A1(\fifo_bank_register.bank[9][75] ),
    .A2(_02550_),
    .B1(_02595_),
    .C1(_02596_),
    .D1(_02597_),
    .X(_02598_));
 sky130_fd_sc_hd__mux2_1 _14238_ (.A0(\fifo_bank_register.bank[0][75] ),
    .A1(_02598_),
    .S(_02563_),
    .X(_02599_));
 sky130_fd_sc_hd__mux2_1 _14239_ (.A0(_02599_),
    .A1(\fifo_bank_register.data_out[75] ),
    .S(_02533_),
    .X(_02600_));
 sky130_fd_sc_hd__clkbuf_1 _14240_ (.A(_02600_),
    .X(_01516_));
 sky130_fd_sc_hd__a22o_1 _14241_ (.A1(\fifo_bank_register.bank[5][76] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][76] ),
    .X(_02601_));
 sky130_fd_sc_hd__a221o_1 _14242_ (.A1(\fifo_bank_register.bank[7][76] ),
    .A2(_02542_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][76] ),
    .C1(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__a22o_1 _14243_ (.A1(\fifo_bank_register.bank[6][76] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][76] ),
    .X(_02603_));
 sky130_fd_sc_hd__a22o_1 _14244_ (.A1(\fifo_bank_register.bank[1][76] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][76] ),
    .X(_02604_));
 sky130_fd_sc_hd__a2111o_1 _14245_ (.A1(\fifo_bank_register.bank[9][76] ),
    .A2(_02550_),
    .B1(_02602_),
    .C1(_02603_),
    .D1(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__mux2_1 _14246_ (.A0(\fifo_bank_register.bank[0][76] ),
    .A1(_02605_),
    .S(_02563_),
    .X(_02606_));
 sky130_fd_sc_hd__mux2_1 _14247_ (.A0(_02606_),
    .A1(\fifo_bank_register.data_out[76] ),
    .S(_02533_),
    .X(_02607_));
 sky130_fd_sc_hd__clkbuf_1 _14248_ (.A(_02607_),
    .X(_01517_));
 sky130_fd_sc_hd__a22o_1 _14249_ (.A1(\fifo_bank_register.bank[5][77] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][77] ),
    .X(_02608_));
 sky130_fd_sc_hd__a221o_1 _14250_ (.A1(\fifo_bank_register.bank[7][77] ),
    .A2(_02542_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][77] ),
    .C1(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__a22o_1 _14251_ (.A1(\fifo_bank_register.bank[6][77] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][77] ),
    .X(_02610_));
 sky130_fd_sc_hd__a22o_1 _14252_ (.A1(\fifo_bank_register.bank[1][77] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][77] ),
    .X(_02611_));
 sky130_fd_sc_hd__a2111o_1 _14253_ (.A1(\fifo_bank_register.bank[9][77] ),
    .A2(_02550_),
    .B1(_02609_),
    .C1(_02610_),
    .D1(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__mux2_1 _14254_ (.A0(\fifo_bank_register.bank[0][77] ),
    .A1(_02612_),
    .S(_02563_),
    .X(_02613_));
 sky130_fd_sc_hd__clkbuf_8 _14255_ (.A(_08068_),
    .X(_02614_));
 sky130_fd_sc_hd__mux2_1 _14256_ (.A0(_02613_),
    .A1(\fifo_bank_register.data_out[77] ),
    .S(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__clkbuf_1 _14257_ (.A(_02615_),
    .X(_01518_));
 sky130_fd_sc_hd__a22o_1 _14258_ (.A1(\fifo_bank_register.bank[5][78] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][78] ),
    .X(_02616_));
 sky130_fd_sc_hd__a221o_1 _14259_ (.A1(\fifo_bank_register.bank[7][78] ),
    .A2(_02542_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][78] ),
    .C1(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__a22o_1 _14260_ (.A1(\fifo_bank_register.bank[6][78] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][78] ),
    .X(_02618_));
 sky130_fd_sc_hd__a22o_1 _14261_ (.A1(\fifo_bank_register.bank[1][78] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][78] ),
    .X(_02619_));
 sky130_fd_sc_hd__a2111o_1 _14262_ (.A1(\fifo_bank_register.bank[9][78] ),
    .A2(_02550_),
    .B1(_02617_),
    .C1(_02618_),
    .D1(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__mux2_1 _14263_ (.A0(\fifo_bank_register.bank[0][78] ),
    .A1(_02620_),
    .S(_02563_),
    .X(_02621_));
 sky130_fd_sc_hd__mux2_1 _14264_ (.A0(_02621_),
    .A1(\fifo_bank_register.data_out[78] ),
    .S(_02614_),
    .X(_02622_));
 sky130_fd_sc_hd__clkbuf_1 _14265_ (.A(_02622_),
    .X(_01519_));
 sky130_fd_sc_hd__clkbuf_4 _14266_ (.A(_08181_),
    .X(_02623_));
 sky130_fd_sc_hd__a22o_1 _14267_ (.A1(\fifo_bank_register.bank[5][79] ),
    .A2(_02552_),
    .B1(_02553_),
    .B2(\fifo_bank_register.bank[3][79] ),
    .X(_02624_));
 sky130_fd_sc_hd__a221o_1 _14268_ (.A1(\fifo_bank_register.bank[7][79] ),
    .A2(_02623_),
    .B1(_02551_),
    .B2(\fifo_bank_register.bank[2][79] ),
    .C1(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__a22o_1 _14269_ (.A1(\fifo_bank_register.bank[6][79] ),
    .A2(_02556_),
    .B1(_02557_),
    .B2(\fifo_bank_register.bank[4][79] ),
    .X(_02626_));
 sky130_fd_sc_hd__a22o_1 _14270_ (.A1(\fifo_bank_register.bank[1][79] ),
    .A2(_02559_),
    .B1(_02560_),
    .B2(\fifo_bank_register.bank[8][79] ),
    .X(_02627_));
 sky130_fd_sc_hd__a2111o_1 _14271_ (.A1(\fifo_bank_register.bank[9][79] ),
    .A2(_02550_),
    .B1(_02625_),
    .C1(_02626_),
    .D1(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__mux2_1 _14272_ (.A0(\fifo_bank_register.bank[0][79] ),
    .A1(_02628_),
    .S(_02563_),
    .X(_02629_));
 sky130_fd_sc_hd__mux2_1 _14273_ (.A0(_02629_),
    .A1(\fifo_bank_register.data_out[79] ),
    .S(_02614_),
    .X(_02630_));
 sky130_fd_sc_hd__clkbuf_1 _14274_ (.A(_02630_),
    .X(_01520_));
 sky130_fd_sc_hd__clkbuf_4 _14275_ (.A(_02136_),
    .X(_02631_));
 sky130_fd_sc_hd__clkbuf_4 _14276_ (.A(_02138_),
    .X(_02632_));
 sky130_fd_sc_hd__clkbuf_4 _14277_ (.A(_02140_),
    .X(_02633_));
 sky130_fd_sc_hd__clkbuf_4 _14278_ (.A(_02142_),
    .X(_02634_));
 sky130_fd_sc_hd__a22o_1 _14279_ (.A1(\fifo_bank_register.bank[5][80] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][80] ),
    .X(_02635_));
 sky130_fd_sc_hd__a221o_1 _14280_ (.A1(\fifo_bank_register.bank[7][80] ),
    .A2(_02623_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][80] ),
    .C1(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__clkbuf_4 _14281_ (.A(_02146_),
    .X(_02637_));
 sky130_fd_sc_hd__clkbuf_4 _14282_ (.A(_02148_),
    .X(_02638_));
 sky130_fd_sc_hd__a22o_1 _14283_ (.A1(\fifo_bank_register.bank[6][80] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][80] ),
    .X(_02639_));
 sky130_fd_sc_hd__clkbuf_4 _14284_ (.A(_02151_),
    .X(_02640_));
 sky130_fd_sc_hd__clkbuf_4 _14285_ (.A(_02153_),
    .X(_02641_));
 sky130_fd_sc_hd__a22o_1 _14286_ (.A1(\fifo_bank_register.bank[1][80] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][80] ),
    .X(_02642_));
 sky130_fd_sc_hd__a2111o_1 _14287_ (.A1(\fifo_bank_register.bank[9][80] ),
    .A2(_02631_),
    .B1(_02636_),
    .C1(_02639_),
    .D1(_02642_),
    .X(_02643_));
 sky130_fd_sc_hd__buf_4 _14288_ (.A(_02157_),
    .X(_02644_));
 sky130_fd_sc_hd__mux2_1 _14289_ (.A0(\fifo_bank_register.bank[0][80] ),
    .A1(_02643_),
    .S(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__mux2_1 _14290_ (.A0(_02645_),
    .A1(\fifo_bank_register.data_out[80] ),
    .S(_02614_),
    .X(_02646_));
 sky130_fd_sc_hd__clkbuf_1 _14291_ (.A(_02646_),
    .X(_01521_));
 sky130_fd_sc_hd__a22o_1 _14292_ (.A1(\fifo_bank_register.bank[5][81] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][81] ),
    .X(_02647_));
 sky130_fd_sc_hd__a221o_1 _14293_ (.A1(\fifo_bank_register.bank[7][81] ),
    .A2(_02623_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][81] ),
    .C1(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__a22o_1 _14294_ (.A1(\fifo_bank_register.bank[6][81] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][81] ),
    .X(_02649_));
 sky130_fd_sc_hd__a22o_1 _14295_ (.A1(\fifo_bank_register.bank[1][81] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][81] ),
    .X(_02650_));
 sky130_fd_sc_hd__a2111o_1 _14296_ (.A1(\fifo_bank_register.bank[9][81] ),
    .A2(_02631_),
    .B1(_02648_),
    .C1(_02649_),
    .D1(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__mux2_1 _14297_ (.A0(\fifo_bank_register.bank[0][81] ),
    .A1(_02651_),
    .S(_02644_),
    .X(_02652_));
 sky130_fd_sc_hd__mux2_1 _14298_ (.A0(_02652_),
    .A1(\fifo_bank_register.data_out[81] ),
    .S(_02614_),
    .X(_02653_));
 sky130_fd_sc_hd__clkbuf_1 _14299_ (.A(_02653_),
    .X(_01522_));
 sky130_fd_sc_hd__a22o_1 _14300_ (.A1(\fifo_bank_register.bank[5][82] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][82] ),
    .X(_02654_));
 sky130_fd_sc_hd__a221o_1 _14301_ (.A1(\fifo_bank_register.bank[7][82] ),
    .A2(_02623_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][82] ),
    .C1(_02654_),
    .X(_02655_));
 sky130_fd_sc_hd__a22o_1 _14302_ (.A1(\fifo_bank_register.bank[6][82] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][82] ),
    .X(_02656_));
 sky130_fd_sc_hd__a22o_1 _14303_ (.A1(\fifo_bank_register.bank[1][82] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][82] ),
    .X(_02657_));
 sky130_fd_sc_hd__a2111o_1 _14304_ (.A1(\fifo_bank_register.bank[9][82] ),
    .A2(_02631_),
    .B1(_02655_),
    .C1(_02656_),
    .D1(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _14305_ (.A0(\fifo_bank_register.bank[0][82] ),
    .A1(_02658_),
    .S(_02644_),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _14306_ (.A0(_02659_),
    .A1(\fifo_bank_register.data_out[82] ),
    .S(_02614_),
    .X(_02660_));
 sky130_fd_sc_hd__clkbuf_1 _14307_ (.A(_02660_),
    .X(_01523_));
 sky130_fd_sc_hd__a22o_1 _14308_ (.A1(\fifo_bank_register.bank[5][83] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][83] ),
    .X(_02661_));
 sky130_fd_sc_hd__a221o_1 _14309_ (.A1(\fifo_bank_register.bank[7][83] ),
    .A2(_02623_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][83] ),
    .C1(_02661_),
    .X(_02662_));
 sky130_fd_sc_hd__a22o_1 _14310_ (.A1(\fifo_bank_register.bank[6][83] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][83] ),
    .X(_02663_));
 sky130_fd_sc_hd__a22o_1 _14311_ (.A1(\fifo_bank_register.bank[1][83] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][83] ),
    .X(_02664_));
 sky130_fd_sc_hd__a2111o_1 _14312_ (.A1(\fifo_bank_register.bank[9][83] ),
    .A2(_02631_),
    .B1(_02662_),
    .C1(_02663_),
    .D1(_02664_),
    .X(_02665_));
 sky130_fd_sc_hd__mux2_1 _14313_ (.A0(\fifo_bank_register.bank[0][83] ),
    .A1(_02665_),
    .S(_02644_),
    .X(_02666_));
 sky130_fd_sc_hd__mux2_1 _14314_ (.A0(_02666_),
    .A1(\fifo_bank_register.data_out[83] ),
    .S(_02614_),
    .X(_02667_));
 sky130_fd_sc_hd__clkbuf_1 _14315_ (.A(_02667_),
    .X(_01524_));
 sky130_fd_sc_hd__a22o_1 _14316_ (.A1(\fifo_bank_register.bank[5][84] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][84] ),
    .X(_02668_));
 sky130_fd_sc_hd__a221o_1 _14317_ (.A1(\fifo_bank_register.bank[7][84] ),
    .A2(_02623_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][84] ),
    .C1(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__a22o_1 _14318_ (.A1(\fifo_bank_register.bank[6][84] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][84] ),
    .X(_02670_));
 sky130_fd_sc_hd__a22o_1 _14319_ (.A1(\fifo_bank_register.bank[1][84] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][84] ),
    .X(_02671_));
 sky130_fd_sc_hd__a2111o_1 _14320_ (.A1(\fifo_bank_register.bank[9][84] ),
    .A2(_02631_),
    .B1(_02669_),
    .C1(_02670_),
    .D1(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__mux2_1 _14321_ (.A0(\fifo_bank_register.bank[0][84] ),
    .A1(_02672_),
    .S(_02644_),
    .X(_02673_));
 sky130_fd_sc_hd__mux2_1 _14322_ (.A0(_02673_),
    .A1(\fifo_bank_register.data_out[84] ),
    .S(_02614_),
    .X(_02674_));
 sky130_fd_sc_hd__clkbuf_1 _14323_ (.A(_02674_),
    .X(_01525_));
 sky130_fd_sc_hd__a22o_1 _14324_ (.A1(\fifo_bank_register.bank[5][85] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][85] ),
    .X(_02675_));
 sky130_fd_sc_hd__a221o_1 _14325_ (.A1(\fifo_bank_register.bank[7][85] ),
    .A2(_02623_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][85] ),
    .C1(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__a22o_1 _14326_ (.A1(\fifo_bank_register.bank[6][85] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][85] ),
    .X(_02677_));
 sky130_fd_sc_hd__a22o_1 _14327_ (.A1(\fifo_bank_register.bank[1][85] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][85] ),
    .X(_02678_));
 sky130_fd_sc_hd__a2111o_1 _14328_ (.A1(\fifo_bank_register.bank[9][85] ),
    .A2(_02631_),
    .B1(_02676_),
    .C1(_02677_),
    .D1(_02678_),
    .X(_02679_));
 sky130_fd_sc_hd__mux2_1 _14329_ (.A0(\fifo_bank_register.bank[0][85] ),
    .A1(_02679_),
    .S(_02644_),
    .X(_02680_));
 sky130_fd_sc_hd__mux2_1 _14330_ (.A0(_02680_),
    .A1(\fifo_bank_register.data_out[85] ),
    .S(_02614_),
    .X(_02681_));
 sky130_fd_sc_hd__clkbuf_1 _14331_ (.A(_02681_),
    .X(_01526_));
 sky130_fd_sc_hd__a22o_1 _14332_ (.A1(\fifo_bank_register.bank[5][86] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][86] ),
    .X(_02682_));
 sky130_fd_sc_hd__a221o_1 _14333_ (.A1(\fifo_bank_register.bank[7][86] ),
    .A2(_02623_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][86] ),
    .C1(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__a22o_1 _14334_ (.A1(\fifo_bank_register.bank[6][86] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][86] ),
    .X(_02684_));
 sky130_fd_sc_hd__a22o_1 _14335_ (.A1(\fifo_bank_register.bank[1][86] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][86] ),
    .X(_02685_));
 sky130_fd_sc_hd__a2111o_1 _14336_ (.A1(\fifo_bank_register.bank[9][86] ),
    .A2(_02631_),
    .B1(_02683_),
    .C1(_02684_),
    .D1(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__mux2_1 _14337_ (.A0(\fifo_bank_register.bank[0][86] ),
    .A1(_02686_),
    .S(_02644_),
    .X(_02687_));
 sky130_fd_sc_hd__mux2_1 _14338_ (.A0(_02687_),
    .A1(\fifo_bank_register.data_out[86] ),
    .S(_02614_),
    .X(_02688_));
 sky130_fd_sc_hd__clkbuf_1 _14339_ (.A(_02688_),
    .X(_01527_));
 sky130_fd_sc_hd__a22o_1 _14340_ (.A1(\fifo_bank_register.bank[5][87] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][87] ),
    .X(_02689_));
 sky130_fd_sc_hd__a221o_1 _14341_ (.A1(\fifo_bank_register.bank[7][87] ),
    .A2(_02623_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][87] ),
    .C1(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__a22o_1 _14342_ (.A1(\fifo_bank_register.bank[6][87] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][87] ),
    .X(_02691_));
 sky130_fd_sc_hd__a22o_1 _14343_ (.A1(\fifo_bank_register.bank[1][87] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][87] ),
    .X(_02692_));
 sky130_fd_sc_hd__a2111o_1 _14344_ (.A1(\fifo_bank_register.bank[9][87] ),
    .A2(_02631_),
    .B1(_02690_),
    .C1(_02691_),
    .D1(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__mux2_1 _14345_ (.A0(\fifo_bank_register.bank[0][87] ),
    .A1(_02693_),
    .S(_02644_),
    .X(_02694_));
 sky130_fd_sc_hd__buf_6 _14346_ (.A(_08063_),
    .X(_02695_));
 sky130_fd_sc_hd__mux2_1 _14347_ (.A0(_02694_),
    .A1(\fifo_bank_register.data_out[87] ),
    .S(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__clkbuf_1 _14348_ (.A(_02696_),
    .X(_01528_));
 sky130_fd_sc_hd__a22o_1 _14349_ (.A1(\fifo_bank_register.bank[5][88] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][88] ),
    .X(_02697_));
 sky130_fd_sc_hd__a221o_1 _14350_ (.A1(\fifo_bank_register.bank[7][88] ),
    .A2(_02623_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][88] ),
    .C1(_02697_),
    .X(_02698_));
 sky130_fd_sc_hd__a22o_1 _14351_ (.A1(\fifo_bank_register.bank[6][88] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][88] ),
    .X(_02699_));
 sky130_fd_sc_hd__a22o_1 _14352_ (.A1(\fifo_bank_register.bank[1][88] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][88] ),
    .X(_02700_));
 sky130_fd_sc_hd__a2111o_1 _14353_ (.A1(\fifo_bank_register.bank[9][88] ),
    .A2(_02631_),
    .B1(_02698_),
    .C1(_02699_),
    .D1(_02700_),
    .X(_02701_));
 sky130_fd_sc_hd__mux2_1 _14354_ (.A0(\fifo_bank_register.bank[0][88] ),
    .A1(_02701_),
    .S(_02644_),
    .X(_02702_));
 sky130_fd_sc_hd__mux2_1 _14355_ (.A0(_02702_),
    .A1(\fifo_bank_register.data_out[88] ),
    .S(_02695_),
    .X(_02703_));
 sky130_fd_sc_hd__clkbuf_1 _14356_ (.A(_02703_),
    .X(_01529_));
 sky130_fd_sc_hd__clkbuf_8 _14357_ (.A(_08181_),
    .X(_02704_));
 sky130_fd_sc_hd__a22o_1 _14358_ (.A1(\fifo_bank_register.bank[5][89] ),
    .A2(_02633_),
    .B1(_02634_),
    .B2(\fifo_bank_register.bank[3][89] ),
    .X(_02705_));
 sky130_fd_sc_hd__a221o_1 _14359_ (.A1(\fifo_bank_register.bank[7][89] ),
    .A2(_02704_),
    .B1(_02632_),
    .B2(\fifo_bank_register.bank[2][89] ),
    .C1(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__a22o_1 _14360_ (.A1(\fifo_bank_register.bank[6][89] ),
    .A2(_02637_),
    .B1(_02638_),
    .B2(\fifo_bank_register.bank[4][89] ),
    .X(_02707_));
 sky130_fd_sc_hd__a22o_1 _14361_ (.A1(\fifo_bank_register.bank[1][89] ),
    .A2(_02640_),
    .B1(_02641_),
    .B2(\fifo_bank_register.bank[8][89] ),
    .X(_02708_));
 sky130_fd_sc_hd__a2111o_1 _14362_ (.A1(\fifo_bank_register.bank[9][89] ),
    .A2(_02631_),
    .B1(_02706_),
    .C1(_02707_),
    .D1(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__mux2_2 _14363_ (.A0(\fifo_bank_register.bank[0][89] ),
    .A1(_02709_),
    .S(_02644_),
    .X(_02710_));
 sky130_fd_sc_hd__mux2_1 _14364_ (.A0(_02710_),
    .A1(\fifo_bank_register.data_out[89] ),
    .S(_02695_),
    .X(_02711_));
 sky130_fd_sc_hd__clkbuf_1 _14365_ (.A(_02711_),
    .X(_01530_));
 sky130_fd_sc_hd__clkbuf_4 _14366_ (.A(_02136_),
    .X(_02712_));
 sky130_fd_sc_hd__clkbuf_4 _14367_ (.A(_02138_),
    .X(_02713_));
 sky130_fd_sc_hd__clkbuf_4 _14368_ (.A(_02140_),
    .X(_02714_));
 sky130_fd_sc_hd__clkbuf_4 _14369_ (.A(_02142_),
    .X(_02715_));
 sky130_fd_sc_hd__a22o_1 _14370_ (.A1(\fifo_bank_register.bank[5][90] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][90] ),
    .X(_02716_));
 sky130_fd_sc_hd__a221o_1 _14371_ (.A1(\fifo_bank_register.bank[7][90] ),
    .A2(_02704_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][90] ),
    .C1(_02716_),
    .X(_02717_));
 sky130_fd_sc_hd__clkbuf_4 _14372_ (.A(_02146_),
    .X(_02718_));
 sky130_fd_sc_hd__clkbuf_4 _14373_ (.A(_02148_),
    .X(_02719_));
 sky130_fd_sc_hd__a22o_1 _14374_ (.A1(\fifo_bank_register.bank[6][90] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][90] ),
    .X(_02720_));
 sky130_fd_sc_hd__clkbuf_4 _14375_ (.A(_02151_),
    .X(_02721_));
 sky130_fd_sc_hd__clkbuf_4 _14376_ (.A(_02153_),
    .X(_02722_));
 sky130_fd_sc_hd__a22o_1 _14377_ (.A1(\fifo_bank_register.bank[1][90] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][90] ),
    .X(_02723_));
 sky130_fd_sc_hd__a2111o_1 _14378_ (.A1(\fifo_bank_register.bank[9][90] ),
    .A2(_02712_),
    .B1(_02717_),
    .C1(_02720_),
    .D1(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__buf_4 _14379_ (.A(_02157_),
    .X(_02725_));
 sky130_fd_sc_hd__mux2_1 _14380_ (.A0(\fifo_bank_register.bank[0][90] ),
    .A1(_02724_),
    .S(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__mux2_1 _14381_ (.A0(_02726_),
    .A1(\fifo_bank_register.data_out[90] ),
    .S(_02695_),
    .X(_02727_));
 sky130_fd_sc_hd__clkbuf_1 _14382_ (.A(_02727_),
    .X(_01531_));
 sky130_fd_sc_hd__a22o_1 _14383_ (.A1(\fifo_bank_register.bank[5][91] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][91] ),
    .X(_02728_));
 sky130_fd_sc_hd__a221o_1 _14384_ (.A1(\fifo_bank_register.bank[7][91] ),
    .A2(_02704_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][91] ),
    .C1(_02728_),
    .X(_02729_));
 sky130_fd_sc_hd__a22o_1 _14385_ (.A1(\fifo_bank_register.bank[6][91] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][91] ),
    .X(_02730_));
 sky130_fd_sc_hd__a22o_1 _14386_ (.A1(\fifo_bank_register.bank[1][91] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][91] ),
    .X(_02731_));
 sky130_fd_sc_hd__a2111o_1 _14387_ (.A1(\fifo_bank_register.bank[9][91] ),
    .A2(_02712_),
    .B1(_02729_),
    .C1(_02730_),
    .D1(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__mux2_2 _14388_ (.A0(\fifo_bank_register.bank[0][91] ),
    .A1(_02732_),
    .S(_02725_),
    .X(_02733_));
 sky130_fd_sc_hd__mux2_1 _14389_ (.A0(_02733_),
    .A1(\fifo_bank_register.data_out[91] ),
    .S(_02695_),
    .X(_02734_));
 sky130_fd_sc_hd__clkbuf_1 _14390_ (.A(_02734_),
    .X(_01532_));
 sky130_fd_sc_hd__a22o_1 _14391_ (.A1(\fifo_bank_register.bank[5][92] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][92] ),
    .X(_02735_));
 sky130_fd_sc_hd__a221o_1 _14392_ (.A1(\fifo_bank_register.bank[7][92] ),
    .A2(_02704_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][92] ),
    .C1(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__a22o_1 _14393_ (.A1(\fifo_bank_register.bank[6][92] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][92] ),
    .X(_02737_));
 sky130_fd_sc_hd__a22o_1 _14394_ (.A1(\fifo_bank_register.bank[1][92] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][92] ),
    .X(_02738_));
 sky130_fd_sc_hd__a2111o_1 _14395_ (.A1(\fifo_bank_register.bank[9][92] ),
    .A2(_02712_),
    .B1(_02736_),
    .C1(_02737_),
    .D1(_02738_),
    .X(_02739_));
 sky130_fd_sc_hd__mux2_1 _14396_ (.A0(\fifo_bank_register.bank[0][92] ),
    .A1(_02739_),
    .S(_02725_),
    .X(_02740_));
 sky130_fd_sc_hd__mux2_1 _14397_ (.A0(_02740_),
    .A1(\fifo_bank_register.data_out[92] ),
    .S(_02695_),
    .X(_02741_));
 sky130_fd_sc_hd__clkbuf_1 _14398_ (.A(_02741_),
    .X(_01533_));
 sky130_fd_sc_hd__a22o_1 _14399_ (.A1(\fifo_bank_register.bank[5][93] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][93] ),
    .X(_02742_));
 sky130_fd_sc_hd__a221o_1 _14400_ (.A1(\fifo_bank_register.bank[7][93] ),
    .A2(_02704_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][93] ),
    .C1(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__a22o_1 _14401_ (.A1(\fifo_bank_register.bank[6][93] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][93] ),
    .X(_02744_));
 sky130_fd_sc_hd__a22o_1 _14402_ (.A1(\fifo_bank_register.bank[1][93] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][93] ),
    .X(_02745_));
 sky130_fd_sc_hd__a2111o_1 _14403_ (.A1(\fifo_bank_register.bank[9][93] ),
    .A2(_02712_),
    .B1(_02743_),
    .C1(_02744_),
    .D1(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__mux2_1 _14404_ (.A0(\fifo_bank_register.bank[0][93] ),
    .A1(_02746_),
    .S(_02725_),
    .X(_02747_));
 sky130_fd_sc_hd__mux2_1 _14405_ (.A0(_02747_),
    .A1(\fifo_bank_register.data_out[93] ),
    .S(_02695_),
    .X(_02748_));
 sky130_fd_sc_hd__clkbuf_1 _14406_ (.A(_02748_),
    .X(_01534_));
 sky130_fd_sc_hd__a22o_1 _14407_ (.A1(\fifo_bank_register.bank[5][94] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][94] ),
    .X(_02749_));
 sky130_fd_sc_hd__a221o_1 _14408_ (.A1(\fifo_bank_register.bank[7][94] ),
    .A2(_02704_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][94] ),
    .C1(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__a22o_1 _14409_ (.A1(\fifo_bank_register.bank[6][94] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][94] ),
    .X(_02751_));
 sky130_fd_sc_hd__a22o_1 _14410_ (.A1(\fifo_bank_register.bank[1][94] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][94] ),
    .X(_02752_));
 sky130_fd_sc_hd__a2111o_1 _14411_ (.A1(\fifo_bank_register.bank[9][94] ),
    .A2(_02712_),
    .B1(_02750_),
    .C1(_02751_),
    .D1(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_1 _14412_ (.A0(\fifo_bank_register.bank[0][94] ),
    .A1(_02753_),
    .S(_02725_),
    .X(_02754_));
 sky130_fd_sc_hd__mux2_1 _14413_ (.A0(_02754_),
    .A1(\fifo_bank_register.data_out[94] ),
    .S(_02695_),
    .X(_02755_));
 sky130_fd_sc_hd__clkbuf_1 _14414_ (.A(_02755_),
    .X(_01535_));
 sky130_fd_sc_hd__a22o_1 _14415_ (.A1(\fifo_bank_register.bank[5][95] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][95] ),
    .X(_02756_));
 sky130_fd_sc_hd__a221o_1 _14416_ (.A1(\fifo_bank_register.bank[7][95] ),
    .A2(_02704_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][95] ),
    .C1(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__a22o_1 _14417_ (.A1(\fifo_bank_register.bank[6][95] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][95] ),
    .X(_02758_));
 sky130_fd_sc_hd__a22o_1 _14418_ (.A1(\fifo_bank_register.bank[1][95] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][95] ),
    .X(_02759_));
 sky130_fd_sc_hd__a2111o_1 _14419_ (.A1(\fifo_bank_register.bank[9][95] ),
    .A2(_02712_),
    .B1(_02757_),
    .C1(_02758_),
    .D1(_02759_),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _14420_ (.A0(\fifo_bank_register.bank[0][95] ),
    .A1(_02760_),
    .S(_02725_),
    .X(_02761_));
 sky130_fd_sc_hd__mux2_1 _14421_ (.A0(_02761_),
    .A1(\fifo_bank_register.data_out[95] ),
    .S(_02695_),
    .X(_02762_));
 sky130_fd_sc_hd__clkbuf_1 _14422_ (.A(_02762_),
    .X(_01536_));
 sky130_fd_sc_hd__a22o_1 _14423_ (.A1(\fifo_bank_register.bank[5][96] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][96] ),
    .X(_02763_));
 sky130_fd_sc_hd__a221o_1 _14424_ (.A1(\fifo_bank_register.bank[7][96] ),
    .A2(_02704_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][96] ),
    .C1(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__a22o_1 _14425_ (.A1(\fifo_bank_register.bank[6][96] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][96] ),
    .X(_02765_));
 sky130_fd_sc_hd__a22o_1 _14426_ (.A1(\fifo_bank_register.bank[1][96] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][96] ),
    .X(_02766_));
 sky130_fd_sc_hd__a2111o_1 _14427_ (.A1(\fifo_bank_register.bank[9][96] ),
    .A2(_02712_),
    .B1(_02764_),
    .C1(_02765_),
    .D1(_02766_),
    .X(_02767_));
 sky130_fd_sc_hd__mux2_1 _14428_ (.A0(\fifo_bank_register.bank[0][96] ),
    .A1(_02767_),
    .S(_02725_),
    .X(_02768_));
 sky130_fd_sc_hd__mux2_1 _14429_ (.A0(_02768_),
    .A1(\fifo_bank_register.data_out[96] ),
    .S(_02695_),
    .X(_02769_));
 sky130_fd_sc_hd__clkbuf_1 _14430_ (.A(_02769_),
    .X(_01537_));
 sky130_fd_sc_hd__a22o_1 _14431_ (.A1(\fifo_bank_register.bank[5][97] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][97] ),
    .X(_02770_));
 sky130_fd_sc_hd__a221o_1 _14432_ (.A1(\fifo_bank_register.bank[7][97] ),
    .A2(_02704_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][97] ),
    .C1(_02770_),
    .X(_02771_));
 sky130_fd_sc_hd__a22o_1 _14433_ (.A1(\fifo_bank_register.bank[6][97] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][97] ),
    .X(_02772_));
 sky130_fd_sc_hd__a22o_1 _14434_ (.A1(\fifo_bank_register.bank[1][97] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][97] ),
    .X(_02773_));
 sky130_fd_sc_hd__a2111o_1 _14435_ (.A1(\fifo_bank_register.bank[9][97] ),
    .A2(_02712_),
    .B1(_02771_),
    .C1(_02772_),
    .D1(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _14436_ (.A0(\fifo_bank_register.bank[0][97] ),
    .A1(_02774_),
    .S(_02725_),
    .X(_02775_));
 sky130_fd_sc_hd__buf_4 _14437_ (.A(_08063_),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_1 _14438_ (.A0(_02775_),
    .A1(\fifo_bank_register.data_out[97] ),
    .S(_02776_),
    .X(_02777_));
 sky130_fd_sc_hd__clkbuf_1 _14439_ (.A(_02777_),
    .X(_01538_));
 sky130_fd_sc_hd__a22o_1 _14440_ (.A1(\fifo_bank_register.bank[5][98] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][98] ),
    .X(_02778_));
 sky130_fd_sc_hd__a221o_1 _14441_ (.A1(\fifo_bank_register.bank[7][98] ),
    .A2(_02704_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][98] ),
    .C1(_02778_),
    .X(_02779_));
 sky130_fd_sc_hd__a22o_1 _14442_ (.A1(\fifo_bank_register.bank[6][98] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][98] ),
    .X(_02780_));
 sky130_fd_sc_hd__a22o_1 _14443_ (.A1(\fifo_bank_register.bank[1][98] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][98] ),
    .X(_02781_));
 sky130_fd_sc_hd__a2111o_1 _14444_ (.A1(\fifo_bank_register.bank[9][98] ),
    .A2(_02712_),
    .B1(_02779_),
    .C1(_02780_),
    .D1(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _14445_ (.A0(\fifo_bank_register.bank[0][98] ),
    .A1(_02782_),
    .S(_02725_),
    .X(_02783_));
 sky130_fd_sc_hd__mux2_1 _14446_ (.A0(_02783_),
    .A1(\fifo_bank_register.data_out[98] ),
    .S(_02776_),
    .X(_02784_));
 sky130_fd_sc_hd__clkbuf_1 _14447_ (.A(_02784_),
    .X(_01539_));
 sky130_fd_sc_hd__clkbuf_4 _14448_ (.A(_08181_),
    .X(_02785_));
 sky130_fd_sc_hd__a22o_1 _14449_ (.A1(\fifo_bank_register.bank[5][99] ),
    .A2(_02714_),
    .B1(_02715_),
    .B2(\fifo_bank_register.bank[3][99] ),
    .X(_02786_));
 sky130_fd_sc_hd__a221o_1 _14450_ (.A1(\fifo_bank_register.bank[7][99] ),
    .A2(_02785_),
    .B1(_02713_),
    .B2(\fifo_bank_register.bank[2][99] ),
    .C1(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__a22o_1 _14451_ (.A1(\fifo_bank_register.bank[6][99] ),
    .A2(_02718_),
    .B1(_02719_),
    .B2(\fifo_bank_register.bank[4][99] ),
    .X(_02788_));
 sky130_fd_sc_hd__a22o_1 _14452_ (.A1(\fifo_bank_register.bank[1][99] ),
    .A2(_02721_),
    .B1(_02722_),
    .B2(\fifo_bank_register.bank[8][99] ),
    .X(_02789_));
 sky130_fd_sc_hd__a2111o_1 _14453_ (.A1(\fifo_bank_register.bank[9][99] ),
    .A2(_02712_),
    .B1(_02787_),
    .C1(_02788_),
    .D1(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__mux2_1 _14454_ (.A0(\fifo_bank_register.bank[0][99] ),
    .A1(_02790_),
    .S(_02725_),
    .X(_02791_));
 sky130_fd_sc_hd__mux2_1 _14455_ (.A0(_02791_),
    .A1(\fifo_bank_register.data_out[99] ),
    .S(_02776_),
    .X(_02792_));
 sky130_fd_sc_hd__clkbuf_1 _14456_ (.A(_02792_),
    .X(_01540_));
 sky130_fd_sc_hd__clkbuf_4 _14457_ (.A(_02136_),
    .X(_02793_));
 sky130_fd_sc_hd__clkbuf_4 _14458_ (.A(_02138_),
    .X(_02794_));
 sky130_fd_sc_hd__clkbuf_4 _14459_ (.A(_02140_),
    .X(_02795_));
 sky130_fd_sc_hd__clkbuf_4 _14460_ (.A(_02142_),
    .X(_02796_));
 sky130_fd_sc_hd__a22o_1 _14461_ (.A1(\fifo_bank_register.bank[5][100] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][100] ),
    .X(_02797_));
 sky130_fd_sc_hd__a221o_1 _14462_ (.A1(\fifo_bank_register.bank[7][100] ),
    .A2(_02785_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][100] ),
    .C1(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_4 _14463_ (.A(_02146_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_4 _14464_ (.A(_02148_),
    .X(_02800_));
 sky130_fd_sc_hd__a22o_1 _14465_ (.A1(\fifo_bank_register.bank[6][100] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][100] ),
    .X(_02801_));
 sky130_fd_sc_hd__clkbuf_4 _14466_ (.A(_02151_),
    .X(_02802_));
 sky130_fd_sc_hd__clkbuf_4 _14467_ (.A(_02153_),
    .X(_02803_));
 sky130_fd_sc_hd__a22o_1 _14468_ (.A1(\fifo_bank_register.bank[1][100] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][100] ),
    .X(_02804_));
 sky130_fd_sc_hd__a2111o_1 _14469_ (.A1(\fifo_bank_register.bank[9][100] ),
    .A2(_02793_),
    .B1(_02798_),
    .C1(_02801_),
    .D1(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__buf_4 _14470_ (.A(_02157_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _14471_ (.A0(\fifo_bank_register.bank[0][100] ),
    .A1(_02805_),
    .S(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _14472_ (.A0(_02807_),
    .A1(\fifo_bank_register.data_out[100] ),
    .S(_02776_),
    .X(_02808_));
 sky130_fd_sc_hd__clkbuf_1 _14473_ (.A(_02808_),
    .X(_01541_));
 sky130_fd_sc_hd__a22o_1 _14474_ (.A1(\fifo_bank_register.bank[5][101] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][101] ),
    .X(_02809_));
 sky130_fd_sc_hd__a221o_1 _14475_ (.A1(\fifo_bank_register.bank[7][101] ),
    .A2(_02785_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][101] ),
    .C1(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__a22o_1 _14476_ (.A1(\fifo_bank_register.bank[6][101] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][101] ),
    .X(_02811_));
 sky130_fd_sc_hd__a22o_1 _14477_ (.A1(\fifo_bank_register.bank[1][101] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][101] ),
    .X(_02812_));
 sky130_fd_sc_hd__a2111o_1 _14478_ (.A1(\fifo_bank_register.bank[9][101] ),
    .A2(_02793_),
    .B1(_02810_),
    .C1(_02811_),
    .D1(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _14479_ (.A0(\fifo_bank_register.bank[0][101] ),
    .A1(_02813_),
    .S(_02806_),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_1 _14480_ (.A0(_02814_),
    .A1(\fifo_bank_register.data_out[101] ),
    .S(_02776_),
    .X(_02815_));
 sky130_fd_sc_hd__clkbuf_1 _14481_ (.A(_02815_),
    .X(_01542_));
 sky130_fd_sc_hd__a22o_1 _14482_ (.A1(\fifo_bank_register.bank[5][102] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][102] ),
    .X(_02816_));
 sky130_fd_sc_hd__a221o_1 _14483_ (.A1(\fifo_bank_register.bank[7][102] ),
    .A2(_02785_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][102] ),
    .C1(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__a22o_1 _14484_ (.A1(\fifo_bank_register.bank[6][102] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][102] ),
    .X(_02818_));
 sky130_fd_sc_hd__a22o_1 _14485_ (.A1(\fifo_bank_register.bank[1][102] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][102] ),
    .X(_02819_));
 sky130_fd_sc_hd__a2111o_1 _14486_ (.A1(\fifo_bank_register.bank[9][102] ),
    .A2(_02793_),
    .B1(_02817_),
    .C1(_02818_),
    .D1(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__mux2_1 _14487_ (.A0(\fifo_bank_register.bank[0][102] ),
    .A1(_02820_),
    .S(_02806_),
    .X(_02821_));
 sky130_fd_sc_hd__mux2_1 _14488_ (.A0(_02821_),
    .A1(\fifo_bank_register.data_out[102] ),
    .S(_02776_),
    .X(_02822_));
 sky130_fd_sc_hd__clkbuf_1 _14489_ (.A(_02822_),
    .X(_01543_));
 sky130_fd_sc_hd__a22o_1 _14490_ (.A1(\fifo_bank_register.bank[5][103] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][103] ),
    .X(_02823_));
 sky130_fd_sc_hd__a221o_1 _14491_ (.A1(\fifo_bank_register.bank[7][103] ),
    .A2(_02785_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][103] ),
    .C1(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__a22o_1 _14492_ (.A1(\fifo_bank_register.bank[6][103] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][103] ),
    .X(_02825_));
 sky130_fd_sc_hd__a22o_1 _14493_ (.A1(\fifo_bank_register.bank[1][103] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][103] ),
    .X(_02826_));
 sky130_fd_sc_hd__a2111o_1 _14494_ (.A1(\fifo_bank_register.bank[9][103] ),
    .A2(_02793_),
    .B1(_02824_),
    .C1(_02825_),
    .D1(_02826_),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _14495_ (.A0(\fifo_bank_register.bank[0][103] ),
    .A1(_02827_),
    .S(_02806_),
    .X(_02828_));
 sky130_fd_sc_hd__mux2_1 _14496_ (.A0(_02828_),
    .A1(\fifo_bank_register.data_out[103] ),
    .S(_02776_),
    .X(_02829_));
 sky130_fd_sc_hd__clkbuf_1 _14497_ (.A(_02829_),
    .X(_01544_));
 sky130_fd_sc_hd__a22o_1 _14498_ (.A1(\fifo_bank_register.bank[5][104] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][104] ),
    .X(_02830_));
 sky130_fd_sc_hd__a221o_1 _14499_ (.A1(\fifo_bank_register.bank[7][104] ),
    .A2(_02785_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][104] ),
    .C1(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__a22o_1 _14500_ (.A1(\fifo_bank_register.bank[6][104] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][104] ),
    .X(_02832_));
 sky130_fd_sc_hd__a22o_1 _14501_ (.A1(\fifo_bank_register.bank[1][104] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][104] ),
    .X(_02833_));
 sky130_fd_sc_hd__a2111o_1 _14502_ (.A1(\fifo_bank_register.bank[9][104] ),
    .A2(_02793_),
    .B1(_02831_),
    .C1(_02832_),
    .D1(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_1 _14503_ (.A0(\fifo_bank_register.bank[0][104] ),
    .A1(_02834_),
    .S(_02806_),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _14504_ (.A0(_02835_),
    .A1(\fifo_bank_register.data_out[104] ),
    .S(_02776_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_1 _14505_ (.A(_02836_),
    .X(_01545_));
 sky130_fd_sc_hd__a22o_1 _14506_ (.A1(\fifo_bank_register.bank[5][105] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][105] ),
    .X(_02837_));
 sky130_fd_sc_hd__a221o_1 _14507_ (.A1(\fifo_bank_register.bank[7][105] ),
    .A2(_02785_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][105] ),
    .C1(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__a22o_1 _14508_ (.A1(\fifo_bank_register.bank[6][105] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][105] ),
    .X(_02839_));
 sky130_fd_sc_hd__a22o_1 _14509_ (.A1(\fifo_bank_register.bank[1][105] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][105] ),
    .X(_02840_));
 sky130_fd_sc_hd__a2111o_1 _14510_ (.A1(\fifo_bank_register.bank[9][105] ),
    .A2(_02793_),
    .B1(_02838_),
    .C1(_02839_),
    .D1(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__mux2_1 _14511_ (.A0(\fifo_bank_register.bank[0][105] ),
    .A1(_02841_),
    .S(_02806_),
    .X(_02842_));
 sky130_fd_sc_hd__mux2_1 _14512_ (.A0(_02842_),
    .A1(\fifo_bank_register.data_out[105] ),
    .S(_02776_),
    .X(_02843_));
 sky130_fd_sc_hd__clkbuf_1 _14513_ (.A(_02843_),
    .X(_01546_));
 sky130_fd_sc_hd__a22o_1 _14514_ (.A1(\fifo_bank_register.bank[5][106] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][106] ),
    .X(_02844_));
 sky130_fd_sc_hd__a221o_1 _14515_ (.A1(\fifo_bank_register.bank[7][106] ),
    .A2(_02785_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][106] ),
    .C1(_02844_),
    .X(_02845_));
 sky130_fd_sc_hd__a22o_1 _14516_ (.A1(\fifo_bank_register.bank[6][106] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][106] ),
    .X(_02846_));
 sky130_fd_sc_hd__a22o_1 _14517_ (.A1(\fifo_bank_register.bank[1][106] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][106] ),
    .X(_02847_));
 sky130_fd_sc_hd__a2111o_1 _14518_ (.A1(\fifo_bank_register.bank[9][106] ),
    .A2(_02793_),
    .B1(_02845_),
    .C1(_02846_),
    .D1(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__mux2_1 _14519_ (.A0(\fifo_bank_register.bank[0][106] ),
    .A1(_02848_),
    .S(_02806_),
    .X(_02849_));
 sky130_fd_sc_hd__mux2_1 _14520_ (.A0(_02849_),
    .A1(\fifo_bank_register.data_out[106] ),
    .S(_02776_),
    .X(_02850_));
 sky130_fd_sc_hd__clkbuf_1 _14521_ (.A(_02850_),
    .X(_01547_));
 sky130_fd_sc_hd__a22o_1 _14522_ (.A1(\fifo_bank_register.bank[5][107] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][107] ),
    .X(_02851_));
 sky130_fd_sc_hd__a221o_1 _14523_ (.A1(\fifo_bank_register.bank[7][107] ),
    .A2(_02785_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][107] ),
    .C1(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__a22o_1 _14524_ (.A1(\fifo_bank_register.bank[6][107] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][107] ),
    .X(_02853_));
 sky130_fd_sc_hd__a22o_1 _14525_ (.A1(\fifo_bank_register.bank[1][107] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][107] ),
    .X(_02854_));
 sky130_fd_sc_hd__a2111o_1 _14526_ (.A1(\fifo_bank_register.bank[9][107] ),
    .A2(_02793_),
    .B1(_02852_),
    .C1(_02853_),
    .D1(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__mux2_1 _14527_ (.A0(\fifo_bank_register.bank[0][107] ),
    .A1(_02855_),
    .S(_02806_),
    .X(_02856_));
 sky130_fd_sc_hd__buf_4 _14528_ (.A(_08063_),
    .X(_02857_));
 sky130_fd_sc_hd__mux2_1 _14529_ (.A0(_02856_),
    .A1(\fifo_bank_register.data_out[107] ),
    .S(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__clkbuf_1 _14530_ (.A(_02858_),
    .X(_01548_));
 sky130_fd_sc_hd__a22o_1 _14531_ (.A1(\fifo_bank_register.bank[5][108] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][108] ),
    .X(_02859_));
 sky130_fd_sc_hd__a221o_1 _14532_ (.A1(\fifo_bank_register.bank[7][108] ),
    .A2(_02785_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][108] ),
    .C1(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__a22o_1 _14533_ (.A1(\fifo_bank_register.bank[6][108] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][108] ),
    .X(_02861_));
 sky130_fd_sc_hd__a22o_1 _14534_ (.A1(\fifo_bank_register.bank[1][108] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][108] ),
    .X(_02862_));
 sky130_fd_sc_hd__a2111o_1 _14535_ (.A1(\fifo_bank_register.bank[9][108] ),
    .A2(_02793_),
    .B1(_02860_),
    .C1(_02861_),
    .D1(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__mux2_1 _14536_ (.A0(\fifo_bank_register.bank[0][108] ),
    .A1(_02863_),
    .S(_02806_),
    .X(_02864_));
 sky130_fd_sc_hd__mux2_1 _14537_ (.A0(_02864_),
    .A1(\fifo_bank_register.data_out[108] ),
    .S(_02857_),
    .X(_02865_));
 sky130_fd_sc_hd__clkbuf_1 _14538_ (.A(_02865_),
    .X(_01549_));
 sky130_fd_sc_hd__clkbuf_4 _14539_ (.A(_08076_),
    .X(_02866_));
 sky130_fd_sc_hd__a22o_1 _14540_ (.A1(\fifo_bank_register.bank[5][109] ),
    .A2(_02795_),
    .B1(_02796_),
    .B2(\fifo_bank_register.bank[3][109] ),
    .X(_02867_));
 sky130_fd_sc_hd__a221o_1 _14541_ (.A1(\fifo_bank_register.bank[7][109] ),
    .A2(_02866_),
    .B1(_02794_),
    .B2(\fifo_bank_register.bank[2][109] ),
    .C1(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__a22o_1 _14542_ (.A1(\fifo_bank_register.bank[6][109] ),
    .A2(_02799_),
    .B1(_02800_),
    .B2(\fifo_bank_register.bank[4][109] ),
    .X(_02869_));
 sky130_fd_sc_hd__a22o_1 _14543_ (.A1(\fifo_bank_register.bank[1][109] ),
    .A2(_02802_),
    .B1(_02803_),
    .B2(\fifo_bank_register.bank[8][109] ),
    .X(_02870_));
 sky130_fd_sc_hd__a2111o_1 _14544_ (.A1(\fifo_bank_register.bank[9][109] ),
    .A2(_02793_),
    .B1(_02868_),
    .C1(_02869_),
    .D1(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__mux2_1 _14545_ (.A0(\fifo_bank_register.bank[0][109] ),
    .A1(_02871_),
    .S(_02806_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _14546_ (.A0(_02872_),
    .A1(\fifo_bank_register.data_out[109] ),
    .S(_02857_),
    .X(_02873_));
 sky130_fd_sc_hd__clkbuf_1 _14547_ (.A(_02873_),
    .X(_01550_));
 sky130_fd_sc_hd__clkbuf_4 _14548_ (.A(_02136_),
    .X(_02874_));
 sky130_fd_sc_hd__clkbuf_4 _14549_ (.A(_02138_),
    .X(_02875_));
 sky130_fd_sc_hd__clkbuf_4 _14550_ (.A(_02140_),
    .X(_02876_));
 sky130_fd_sc_hd__clkbuf_4 _14551_ (.A(_02142_),
    .X(_02877_));
 sky130_fd_sc_hd__a22o_1 _14552_ (.A1(\fifo_bank_register.bank[5][110] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][110] ),
    .X(_02878_));
 sky130_fd_sc_hd__a221o_1 _14553_ (.A1(\fifo_bank_register.bank[7][110] ),
    .A2(_02866_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][110] ),
    .C1(_02878_),
    .X(_02879_));
 sky130_fd_sc_hd__clkbuf_4 _14554_ (.A(_02146_),
    .X(_02880_));
 sky130_fd_sc_hd__clkbuf_4 _14555_ (.A(_02148_),
    .X(_02881_));
 sky130_fd_sc_hd__a22o_1 _14556_ (.A1(\fifo_bank_register.bank[6][110] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][110] ),
    .X(_02882_));
 sky130_fd_sc_hd__clkbuf_4 _14557_ (.A(_02151_),
    .X(_02883_));
 sky130_fd_sc_hd__clkbuf_4 _14558_ (.A(_02153_),
    .X(_02884_));
 sky130_fd_sc_hd__a22o_1 _14559_ (.A1(\fifo_bank_register.bank[1][110] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][110] ),
    .X(_02885_));
 sky130_fd_sc_hd__a2111o_1 _14560_ (.A1(\fifo_bank_register.bank[9][110] ),
    .A2(_02874_),
    .B1(_02879_),
    .C1(_02882_),
    .D1(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__buf_4 _14561_ (.A(_02157_),
    .X(_02887_));
 sky130_fd_sc_hd__mux2_1 _14562_ (.A0(\fifo_bank_register.bank[0][110] ),
    .A1(_02886_),
    .S(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__mux2_1 _14563_ (.A0(_02888_),
    .A1(\fifo_bank_register.data_out[110] ),
    .S(_02857_),
    .X(_02889_));
 sky130_fd_sc_hd__clkbuf_1 _14564_ (.A(_02889_),
    .X(_01551_));
 sky130_fd_sc_hd__a22o_1 _14565_ (.A1(\fifo_bank_register.bank[5][111] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][111] ),
    .X(_02890_));
 sky130_fd_sc_hd__a221o_1 _14566_ (.A1(\fifo_bank_register.bank[7][111] ),
    .A2(_02866_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][111] ),
    .C1(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__a22o_1 _14567_ (.A1(\fifo_bank_register.bank[6][111] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][111] ),
    .X(_02892_));
 sky130_fd_sc_hd__a22o_1 _14568_ (.A1(\fifo_bank_register.bank[1][111] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][111] ),
    .X(_02893_));
 sky130_fd_sc_hd__a2111o_1 _14569_ (.A1(\fifo_bank_register.bank[9][111] ),
    .A2(_02874_),
    .B1(_02891_),
    .C1(_02892_),
    .D1(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__mux2_1 _14570_ (.A0(\fifo_bank_register.bank[0][111] ),
    .A1(_02894_),
    .S(_02887_),
    .X(_02895_));
 sky130_fd_sc_hd__mux2_1 _14571_ (.A0(_02895_),
    .A1(\fifo_bank_register.data_out[111] ),
    .S(_02857_),
    .X(_02896_));
 sky130_fd_sc_hd__clkbuf_1 _14572_ (.A(_02896_),
    .X(_01552_));
 sky130_fd_sc_hd__a22o_1 _14573_ (.A1(\fifo_bank_register.bank[5][112] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][112] ),
    .X(_02897_));
 sky130_fd_sc_hd__a221o_1 _14574_ (.A1(\fifo_bank_register.bank[7][112] ),
    .A2(_02866_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][112] ),
    .C1(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__a22o_1 _14575_ (.A1(\fifo_bank_register.bank[6][112] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][112] ),
    .X(_02899_));
 sky130_fd_sc_hd__a22o_1 _14576_ (.A1(\fifo_bank_register.bank[1][112] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][112] ),
    .X(_02900_));
 sky130_fd_sc_hd__a2111o_1 _14577_ (.A1(\fifo_bank_register.bank[9][112] ),
    .A2(_02874_),
    .B1(_02898_),
    .C1(_02899_),
    .D1(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__mux2_1 _14578_ (.A0(\fifo_bank_register.bank[0][112] ),
    .A1(_02901_),
    .S(_02887_),
    .X(_02902_));
 sky130_fd_sc_hd__mux2_1 _14579_ (.A0(_02902_),
    .A1(\fifo_bank_register.data_out[112] ),
    .S(_02857_),
    .X(_02903_));
 sky130_fd_sc_hd__clkbuf_1 _14580_ (.A(_02903_),
    .X(_01553_));
 sky130_fd_sc_hd__a22o_1 _14581_ (.A1(\fifo_bank_register.bank[5][113] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][113] ),
    .X(_02904_));
 sky130_fd_sc_hd__a221o_1 _14582_ (.A1(\fifo_bank_register.bank[7][113] ),
    .A2(_02866_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][113] ),
    .C1(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__a22o_1 _14583_ (.A1(\fifo_bank_register.bank[6][113] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][113] ),
    .X(_02906_));
 sky130_fd_sc_hd__a22o_1 _14584_ (.A1(\fifo_bank_register.bank[1][113] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][113] ),
    .X(_02907_));
 sky130_fd_sc_hd__a2111o_1 _14585_ (.A1(\fifo_bank_register.bank[9][113] ),
    .A2(_02874_),
    .B1(_02905_),
    .C1(_02906_),
    .D1(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__mux2_1 _14586_ (.A0(\fifo_bank_register.bank[0][113] ),
    .A1(_02908_),
    .S(_02887_),
    .X(_02909_));
 sky130_fd_sc_hd__mux2_1 _14587_ (.A0(_02909_),
    .A1(\fifo_bank_register.data_out[113] ),
    .S(_02857_),
    .X(_02910_));
 sky130_fd_sc_hd__clkbuf_1 _14588_ (.A(_02910_),
    .X(_01554_));
 sky130_fd_sc_hd__a22o_1 _14589_ (.A1(\fifo_bank_register.bank[5][114] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][114] ),
    .X(_02911_));
 sky130_fd_sc_hd__a221o_1 _14590_ (.A1(\fifo_bank_register.bank[7][114] ),
    .A2(_02866_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][114] ),
    .C1(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__a22o_1 _14591_ (.A1(\fifo_bank_register.bank[6][114] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][114] ),
    .X(_02913_));
 sky130_fd_sc_hd__a22o_1 _14592_ (.A1(\fifo_bank_register.bank[1][114] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][114] ),
    .X(_02914_));
 sky130_fd_sc_hd__a2111o_1 _14593_ (.A1(\fifo_bank_register.bank[9][114] ),
    .A2(_02874_),
    .B1(_02912_),
    .C1(_02913_),
    .D1(_02914_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _14594_ (.A0(\fifo_bank_register.bank[0][114] ),
    .A1(_02915_),
    .S(_02887_),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _14595_ (.A0(_02916_),
    .A1(\fifo_bank_register.data_out[114] ),
    .S(_02857_),
    .X(_02917_));
 sky130_fd_sc_hd__clkbuf_1 _14596_ (.A(_02917_),
    .X(_01555_));
 sky130_fd_sc_hd__a22o_1 _14597_ (.A1(\fifo_bank_register.bank[5][115] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][115] ),
    .X(_02918_));
 sky130_fd_sc_hd__a221o_1 _14598_ (.A1(\fifo_bank_register.bank[7][115] ),
    .A2(_02866_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][115] ),
    .C1(_02918_),
    .X(_02919_));
 sky130_fd_sc_hd__a22o_1 _14599_ (.A1(\fifo_bank_register.bank[6][115] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][115] ),
    .X(_02920_));
 sky130_fd_sc_hd__a22o_1 _14600_ (.A1(\fifo_bank_register.bank[1][115] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][115] ),
    .X(_02921_));
 sky130_fd_sc_hd__a2111o_1 _14601_ (.A1(\fifo_bank_register.bank[9][115] ),
    .A2(_02874_),
    .B1(_02919_),
    .C1(_02920_),
    .D1(_02921_),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _14602_ (.A0(\fifo_bank_register.bank[0][115] ),
    .A1(_02922_),
    .S(_02887_),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_1 _14603_ (.A0(_02923_),
    .A1(\fifo_bank_register.data_out[115] ),
    .S(_02857_),
    .X(_02924_));
 sky130_fd_sc_hd__clkbuf_1 _14604_ (.A(_02924_),
    .X(_01556_));
 sky130_fd_sc_hd__a22o_1 _14605_ (.A1(\fifo_bank_register.bank[5][116] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][116] ),
    .X(_02925_));
 sky130_fd_sc_hd__a221o_1 _14606_ (.A1(\fifo_bank_register.bank[7][116] ),
    .A2(_02866_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][116] ),
    .C1(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__a22o_1 _14607_ (.A1(\fifo_bank_register.bank[6][116] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][116] ),
    .X(_02927_));
 sky130_fd_sc_hd__a22o_1 _14608_ (.A1(\fifo_bank_register.bank[1][116] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][116] ),
    .X(_02928_));
 sky130_fd_sc_hd__a2111o_1 _14609_ (.A1(\fifo_bank_register.bank[9][116] ),
    .A2(_02874_),
    .B1(_02926_),
    .C1(_02927_),
    .D1(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__mux2_1 _14610_ (.A0(\fifo_bank_register.bank[0][116] ),
    .A1(_02929_),
    .S(_02887_),
    .X(_02930_));
 sky130_fd_sc_hd__mux2_1 _14611_ (.A0(_02930_),
    .A1(\fifo_bank_register.data_out[116] ),
    .S(_02857_),
    .X(_02931_));
 sky130_fd_sc_hd__clkbuf_1 _14612_ (.A(_02931_),
    .X(_01557_));
 sky130_fd_sc_hd__a22o_1 _14613_ (.A1(\fifo_bank_register.bank[5][117] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][117] ),
    .X(_02932_));
 sky130_fd_sc_hd__a221o_1 _14614_ (.A1(\fifo_bank_register.bank[7][117] ),
    .A2(_02866_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][117] ),
    .C1(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__a22o_1 _14615_ (.A1(\fifo_bank_register.bank[6][117] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][117] ),
    .X(_02934_));
 sky130_fd_sc_hd__a22o_1 _14616_ (.A1(\fifo_bank_register.bank[1][117] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][117] ),
    .X(_02935_));
 sky130_fd_sc_hd__a2111o_1 _14617_ (.A1(\fifo_bank_register.bank[9][117] ),
    .A2(_02874_),
    .B1(_02933_),
    .C1(_02934_),
    .D1(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__mux2_1 _14618_ (.A0(\fifo_bank_register.bank[0][117] ),
    .A1(_02936_),
    .S(_02887_),
    .X(_02937_));
 sky130_fd_sc_hd__clkbuf_8 _14619_ (.A(_08063_),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _14620_ (.A0(_02937_),
    .A1(\fifo_bank_register.data_out[117] ),
    .S(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__clkbuf_1 _14621_ (.A(_02939_),
    .X(_01558_));
 sky130_fd_sc_hd__a22o_1 _14622_ (.A1(\fifo_bank_register.bank[5][118] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][118] ),
    .X(_02940_));
 sky130_fd_sc_hd__a221o_1 _14623_ (.A1(\fifo_bank_register.bank[7][118] ),
    .A2(_02866_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][118] ),
    .C1(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__a22o_1 _14624_ (.A1(\fifo_bank_register.bank[6][118] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][118] ),
    .X(_02942_));
 sky130_fd_sc_hd__a22o_1 _14625_ (.A1(\fifo_bank_register.bank[1][118] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][118] ),
    .X(_02943_));
 sky130_fd_sc_hd__a2111o_1 _14626_ (.A1(\fifo_bank_register.bank[9][118] ),
    .A2(_02874_),
    .B1(_02941_),
    .C1(_02942_),
    .D1(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__mux2_1 _14627_ (.A0(\fifo_bank_register.bank[0][118] ),
    .A1(_02944_),
    .S(_02887_),
    .X(_02945_));
 sky130_fd_sc_hd__mux2_1 _14628_ (.A0(_02945_),
    .A1(\fifo_bank_register.data_out[118] ),
    .S(_02938_),
    .X(_02946_));
 sky130_fd_sc_hd__clkbuf_1 _14629_ (.A(_02946_),
    .X(_01559_));
 sky130_fd_sc_hd__a22o_1 _14630_ (.A1(\fifo_bank_register.bank[5][119] ),
    .A2(_02876_),
    .B1(_02877_),
    .B2(\fifo_bank_register.bank[3][119] ),
    .X(_02947_));
 sky130_fd_sc_hd__a221o_1 _14631_ (.A1(\fifo_bank_register.bank[7][119] ),
    .A2(_08077_),
    .B1(_02875_),
    .B2(\fifo_bank_register.bank[2][119] ),
    .C1(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__a22o_1 _14632_ (.A1(\fifo_bank_register.bank[6][119] ),
    .A2(_02880_),
    .B1(_02881_),
    .B2(\fifo_bank_register.bank[4][119] ),
    .X(_02949_));
 sky130_fd_sc_hd__a22o_1 _14633_ (.A1(\fifo_bank_register.bank[1][119] ),
    .A2(_02883_),
    .B1(_02884_),
    .B2(\fifo_bank_register.bank[8][119] ),
    .X(_02950_));
 sky130_fd_sc_hd__a2111o_1 _14634_ (.A1(\fifo_bank_register.bank[9][119] ),
    .A2(_02874_),
    .B1(_02948_),
    .C1(_02949_),
    .D1(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__mux2_1 _14635_ (.A0(\fifo_bank_register.bank[0][119] ),
    .A1(_02951_),
    .S(_02887_),
    .X(_02952_));
 sky130_fd_sc_hd__mux2_1 _14636_ (.A0(_02952_),
    .A1(\fifo_bank_register.data_out[119] ),
    .S(_02938_),
    .X(_02953_));
 sky130_fd_sc_hd__clkbuf_1 _14637_ (.A(_02953_),
    .X(_01560_));
 sky130_fd_sc_hd__a22o_1 _14638_ (.A1(\fifo_bank_register.bank[5][120] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(\fifo_bank_register.bank[3][120] ),
    .X(_02954_));
 sky130_fd_sc_hd__a221o_1 _14639_ (.A1(\fifo_bank_register.bank[7][120] ),
    .A2(_08077_),
    .B1(_08092_),
    .B2(\fifo_bank_register.bank[2][120] ),
    .C1(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__a22o_1 _14640_ (.A1(\fifo_bank_register.bank[6][120] ),
    .A2(_08104_),
    .B1(_08107_),
    .B2(\fifo_bank_register.bank[4][120] ),
    .X(_02956_));
 sky130_fd_sc_hd__a22o_1 _14641_ (.A1(\fifo_bank_register.bank[1][120] ),
    .A2(_08111_),
    .B1(_08114_),
    .B2(\fifo_bank_register.bank[8][120] ),
    .X(_02957_));
 sky130_fd_sc_hd__a2111o_1 _14642_ (.A1(\fifo_bank_register.bank[9][120] ),
    .A2(_08089_),
    .B1(_02955_),
    .C1(_02956_),
    .D1(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__mux2_1 _14643_ (.A0(\fifo_bank_register.bank[0][120] ),
    .A1(_02958_),
    .S(_08120_),
    .X(_02959_));
 sky130_fd_sc_hd__mux2_1 _14644_ (.A0(_02959_),
    .A1(\fifo_bank_register.data_out[120] ),
    .S(_02938_),
    .X(_02960_));
 sky130_fd_sc_hd__clkbuf_1 _14645_ (.A(_02960_),
    .X(_01561_));
 sky130_fd_sc_hd__a22o_1 _14646_ (.A1(\fifo_bank_register.bank[5][121] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(\fifo_bank_register.bank[3][121] ),
    .X(_02961_));
 sky130_fd_sc_hd__a221o_1 _14647_ (.A1(\fifo_bank_register.bank[7][121] ),
    .A2(_08077_),
    .B1(_08092_),
    .B2(\fifo_bank_register.bank[2][121] ),
    .C1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__a22o_1 _14648_ (.A1(\fifo_bank_register.bank[6][121] ),
    .A2(_08104_),
    .B1(_08107_),
    .B2(\fifo_bank_register.bank[4][121] ),
    .X(_02963_));
 sky130_fd_sc_hd__a22o_1 _14649_ (.A1(\fifo_bank_register.bank[1][121] ),
    .A2(_08111_),
    .B1(_08114_),
    .B2(\fifo_bank_register.bank[8][121] ),
    .X(_02964_));
 sky130_fd_sc_hd__a2111o_1 _14650_ (.A1(\fifo_bank_register.bank[9][121] ),
    .A2(_08089_),
    .B1(_02962_),
    .C1(_02963_),
    .D1(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _14651_ (.A0(\fifo_bank_register.bank[0][121] ),
    .A1(_02965_),
    .S(_08120_),
    .X(_02966_));
 sky130_fd_sc_hd__mux2_1 _14652_ (.A0(_02966_),
    .A1(\fifo_bank_register.data_out[121] ),
    .S(_02938_),
    .X(_02967_));
 sky130_fd_sc_hd__clkbuf_1 _14653_ (.A(_02967_),
    .X(_01562_));
 sky130_fd_sc_hd__a22o_1 _14654_ (.A1(\fifo_bank_register.bank[5][122] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(\fifo_bank_register.bank[3][122] ),
    .X(_02968_));
 sky130_fd_sc_hd__a221o_1 _14655_ (.A1(\fifo_bank_register.bank[7][122] ),
    .A2(_08077_),
    .B1(_08092_),
    .B2(\fifo_bank_register.bank[2][122] ),
    .C1(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__a22o_1 _14656_ (.A1(\fifo_bank_register.bank[6][122] ),
    .A2(_08104_),
    .B1(_08107_),
    .B2(\fifo_bank_register.bank[4][122] ),
    .X(_02970_));
 sky130_fd_sc_hd__a22o_1 _14657_ (.A1(\fifo_bank_register.bank[1][122] ),
    .A2(_08111_),
    .B1(_08114_),
    .B2(\fifo_bank_register.bank[8][122] ),
    .X(_02971_));
 sky130_fd_sc_hd__a2111o_1 _14658_ (.A1(\fifo_bank_register.bank[9][122] ),
    .A2(_08089_),
    .B1(_02969_),
    .C1(_02970_),
    .D1(_02971_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _14659_ (.A0(\fifo_bank_register.bank[0][122] ),
    .A1(_02972_),
    .S(_08120_),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_1 _14660_ (.A0(_02973_),
    .A1(\fifo_bank_register.data_out[122] ),
    .S(_02938_),
    .X(_02974_));
 sky130_fd_sc_hd__clkbuf_1 _14661_ (.A(_02974_),
    .X(_01563_));
 sky130_fd_sc_hd__a22o_1 _14662_ (.A1(\fifo_bank_register.bank[5][123] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(\fifo_bank_register.bank[3][123] ),
    .X(_02975_));
 sky130_fd_sc_hd__a221o_1 _14663_ (.A1(\fifo_bank_register.bank[7][123] ),
    .A2(_08077_),
    .B1(_08092_),
    .B2(\fifo_bank_register.bank[2][123] ),
    .C1(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__a22o_1 _14664_ (.A1(\fifo_bank_register.bank[6][123] ),
    .A2(_08104_),
    .B1(_08107_),
    .B2(\fifo_bank_register.bank[4][123] ),
    .X(_02977_));
 sky130_fd_sc_hd__a22o_1 _14665_ (.A1(\fifo_bank_register.bank[1][123] ),
    .A2(_08111_),
    .B1(_08114_),
    .B2(\fifo_bank_register.bank[8][123] ),
    .X(_02978_));
 sky130_fd_sc_hd__a2111o_1 _14666_ (.A1(\fifo_bank_register.bank[9][123] ),
    .A2(_08089_),
    .B1(_02976_),
    .C1(_02977_),
    .D1(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__mux2_1 _14667_ (.A0(\fifo_bank_register.bank[0][123] ),
    .A1(_02979_),
    .S(_08120_),
    .X(_02980_));
 sky130_fd_sc_hd__mux2_1 _14668_ (.A0(_02980_),
    .A1(\fifo_bank_register.data_out[123] ),
    .S(_02938_),
    .X(_02981_));
 sky130_fd_sc_hd__clkbuf_1 _14669_ (.A(_02981_),
    .X(_01564_));
 sky130_fd_sc_hd__a22o_1 _14670_ (.A1(\fifo_bank_register.bank[5][124] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(\fifo_bank_register.bank[3][124] ),
    .X(_02982_));
 sky130_fd_sc_hd__a221o_1 _14671_ (.A1(\fifo_bank_register.bank[7][124] ),
    .A2(_08077_),
    .B1(_08092_),
    .B2(\fifo_bank_register.bank[2][124] ),
    .C1(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__a22o_1 _14672_ (.A1(\fifo_bank_register.bank[6][124] ),
    .A2(_08104_),
    .B1(_08107_),
    .B2(\fifo_bank_register.bank[4][124] ),
    .X(_02984_));
 sky130_fd_sc_hd__a22o_1 _14673_ (.A1(\fifo_bank_register.bank[1][124] ),
    .A2(_08111_),
    .B1(_08114_),
    .B2(\fifo_bank_register.bank[8][124] ),
    .X(_02985_));
 sky130_fd_sc_hd__a2111o_1 _14674_ (.A1(\fifo_bank_register.bank[9][124] ),
    .A2(_08089_),
    .B1(_02983_),
    .C1(_02984_),
    .D1(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__mux2_1 _14675_ (.A0(\fifo_bank_register.bank[0][124] ),
    .A1(_02986_),
    .S(_08120_),
    .X(_02987_));
 sky130_fd_sc_hd__mux2_1 _14676_ (.A0(_02987_),
    .A1(\fifo_bank_register.data_out[124] ),
    .S(_02938_),
    .X(_02988_));
 sky130_fd_sc_hd__clkbuf_1 _14677_ (.A(_02988_),
    .X(_01565_));
 sky130_fd_sc_hd__a22o_1 _14678_ (.A1(\fifo_bank_register.bank[5][125] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(\fifo_bank_register.bank[3][125] ),
    .X(_02989_));
 sky130_fd_sc_hd__a221o_1 _14679_ (.A1(\fifo_bank_register.bank[7][125] ),
    .A2(_08077_),
    .B1(_08092_),
    .B2(\fifo_bank_register.bank[2][125] ),
    .C1(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__a22o_1 _14680_ (.A1(\fifo_bank_register.bank[6][125] ),
    .A2(_08104_),
    .B1(_08107_),
    .B2(\fifo_bank_register.bank[4][125] ),
    .X(_02991_));
 sky130_fd_sc_hd__a22o_1 _14681_ (.A1(\fifo_bank_register.bank[1][125] ),
    .A2(_08111_),
    .B1(_08114_),
    .B2(\fifo_bank_register.bank[8][125] ),
    .X(_02992_));
 sky130_fd_sc_hd__a2111o_1 _14682_ (.A1(\fifo_bank_register.bank[9][125] ),
    .A2(_08089_),
    .B1(_02990_),
    .C1(_02991_),
    .D1(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__mux2_1 _14683_ (.A0(\fifo_bank_register.bank[0][125] ),
    .A1(_02993_),
    .S(_08120_),
    .X(_02994_));
 sky130_fd_sc_hd__mux2_1 _14684_ (.A0(_02994_),
    .A1(\fifo_bank_register.data_out[125] ),
    .S(_02938_),
    .X(_02995_));
 sky130_fd_sc_hd__clkbuf_1 _14685_ (.A(_02995_),
    .X(_01566_));
 sky130_fd_sc_hd__a22o_1 _14686_ (.A1(\fifo_bank_register.bank[5][126] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(\fifo_bank_register.bank[3][126] ),
    .X(_02996_));
 sky130_fd_sc_hd__a221o_1 _14687_ (.A1(\fifo_bank_register.bank[7][126] ),
    .A2(_08077_),
    .B1(_08092_),
    .B2(\fifo_bank_register.bank[2][126] ),
    .C1(_02996_),
    .X(_02997_));
 sky130_fd_sc_hd__a22o_1 _14688_ (.A1(\fifo_bank_register.bank[6][126] ),
    .A2(_08104_),
    .B1(_08107_),
    .B2(\fifo_bank_register.bank[4][126] ),
    .X(_02998_));
 sky130_fd_sc_hd__a22o_1 _14689_ (.A1(\fifo_bank_register.bank[1][126] ),
    .A2(_08111_),
    .B1(_08114_),
    .B2(\fifo_bank_register.bank[8][126] ),
    .X(_02999_));
 sky130_fd_sc_hd__a2111o_1 _14690_ (.A1(\fifo_bank_register.bank[9][126] ),
    .A2(_08089_),
    .B1(_02997_),
    .C1(_02998_),
    .D1(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__mux2_1 _14691_ (.A0(\fifo_bank_register.bank[0][126] ),
    .A1(_03000_),
    .S(_08120_),
    .X(_03001_));
 sky130_fd_sc_hd__mux2_1 _14692_ (.A0(_03001_),
    .A1(\fifo_bank_register.data_out[126] ),
    .S(_02938_),
    .X(_03002_));
 sky130_fd_sc_hd__clkbuf_1 _14693_ (.A(_03002_),
    .X(_01567_));
 sky130_fd_sc_hd__a22o_1 _14694_ (.A1(\fifo_bank_register.bank[5][127] ),
    .A2(_08096_),
    .B1(_08099_),
    .B2(\fifo_bank_register.bank[3][127] ),
    .X(_03003_));
 sky130_fd_sc_hd__a221o_1 _14695_ (.A1(\fifo_bank_register.bank[7][127] ),
    .A2(_08077_),
    .B1(_08092_),
    .B2(\fifo_bank_register.bank[2][127] ),
    .C1(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__a22o_1 _14696_ (.A1(\fifo_bank_register.bank[6][127] ),
    .A2(_08104_),
    .B1(_08107_),
    .B2(\fifo_bank_register.bank[4][127] ),
    .X(_03005_));
 sky130_fd_sc_hd__a22o_1 _14697_ (.A1(\fifo_bank_register.bank[1][127] ),
    .A2(_08111_),
    .B1(_08114_),
    .B2(\fifo_bank_register.bank[8][127] ),
    .X(_03006_));
 sky130_fd_sc_hd__a2111o_1 _14698_ (.A1(\fifo_bank_register.bank[9][127] ),
    .A2(_08089_),
    .B1(_03004_),
    .C1(_03005_),
    .D1(_03006_),
    .X(_03007_));
 sky130_fd_sc_hd__mux2_1 _14699_ (.A0(\fifo_bank_register.bank[0][127] ),
    .A1(_03007_),
    .S(_08120_),
    .X(_03008_));
 sky130_fd_sc_hd__mux2_1 _14700_ (.A0(_03008_),
    .A1(\fifo_bank_register.data_out[127] ),
    .S(_08068_),
    .X(_03009_));
 sky130_fd_sc_hd__clkbuf_1 _14701_ (.A(_03009_),
    .X(_01568_));
 sky130_fd_sc_hd__nor2_4 _14702_ (.A(_04369_),
    .B(_04927_),
    .Y(_03010_));
 sky130_fd_sc_hd__mux2_1 _14703_ (.A0(\sub1.data_o[48] ),
    .A1(\sub1.data_o[112] ),
    .S(_05598_),
    .X(_03011_));
 sky130_fd_sc_hd__a22o_1 _14704_ (.A1(\sub1.data_o[80] ),
    .A2(_03010_),
    .B1(_03011_),
    .B2(\sub1.next_ready_o ),
    .X(_03012_));
 sky130_fd_sc_hd__a31o_1 _14705_ (.A1(_05104_),
    .A2(_04927_),
    .A3(_05548_),
    .B1(_03012_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _14706_ (.A0(\sub1.data_o[49] ),
    .A1(\sub1.data_o[113] ),
    .S(_05598_),
    .X(_03013_));
 sky130_fd_sc_hd__a22o_1 _14707_ (.A1(\sub1.data_o[81] ),
    .A2(_03010_),
    .B1(_03013_),
    .B2(\sub1.next_ready_o ),
    .X(_03014_));
 sky130_fd_sc_hd__a31o_1 _14708_ (.A1(_05104_),
    .A2(_04927_),
    .A3(_05554_),
    .B1(_03014_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _14709_ (.A0(\sub1.data_o[50] ),
    .A1(\sub1.data_o[114] ),
    .S(_05598_),
    .X(_03015_));
 sky130_fd_sc_hd__a22o_1 _14710_ (.A1(\sub1.data_o[82] ),
    .A2(_03010_),
    .B1(_03015_),
    .B2(\sub1.next_ready_o ),
    .X(_03016_));
 sky130_fd_sc_hd__a31o_1 _14711_ (.A1(_05104_),
    .A2(_04927_),
    .A3(_05560_),
    .B1(_03016_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _14712_ (.A0(\sub1.data_o[51] ),
    .A1(\sub1.data_o[115] ),
    .S(_05598_),
    .X(_03017_));
 sky130_fd_sc_hd__a22o_1 _14713_ (.A1(\sub1.data_o[83] ),
    .A2(_03010_),
    .B1(_03017_),
    .B2(\sub1.next_ready_o ),
    .X(_03018_));
 sky130_fd_sc_hd__a31o_1 _14714_ (.A1(_05104_),
    .A2(_04927_),
    .A3(_05196_),
    .B1(_03018_),
    .X(_01572_));
 sky130_fd_sc_hd__clkbuf_4 _14715_ (.A(_05103_),
    .X(_03019_));
 sky130_fd_sc_hd__mux2_1 _14716_ (.A0(\sub1.data_o[52] ),
    .A1(\sub1.data_o[116] ),
    .S(_05598_),
    .X(_03020_));
 sky130_fd_sc_hd__a22o_1 _14717_ (.A1(\sub1.data_o[84] ),
    .A2(_03010_),
    .B1(_03020_),
    .B2(\sub1.next_ready_o ),
    .X(_03021_));
 sky130_fd_sc_hd__a31o_1 _14718_ (.A1(_03019_),
    .A2(_04927_),
    .A3(_05219_),
    .B1(_03021_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _14719_ (.A0(\sub1.data_o[53] ),
    .A1(\sub1.data_o[117] ),
    .S(_05598_),
    .X(_03022_));
 sky130_fd_sc_hd__a22o_1 _14720_ (.A1(\sub1.data_o[85] ),
    .A2(_03010_),
    .B1(_03022_),
    .B2(\sub1.next_ready_o ),
    .X(_03023_));
 sky130_fd_sc_hd__a31o_1 _14721_ (.A1(_03019_),
    .A2(_04927_),
    .A3(_05228_),
    .B1(_03023_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _14722_ (.A0(\sub1.data_o[54] ),
    .A1(\sub1.data_o[118] ),
    .S(_05598_),
    .X(_03024_));
 sky130_fd_sc_hd__a22o_1 _14723_ (.A1(\sub1.data_o[86] ),
    .A2(_03010_),
    .B1(_03024_),
    .B2(\sub1.next_ready_o ),
    .X(_03025_));
 sky130_fd_sc_hd__a31o_1 _14724_ (.A1(_03019_),
    .A2(_04927_),
    .A3(_05236_),
    .B1(_03025_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _14725_ (.A0(\sub1.data_o[55] ),
    .A1(\sub1.data_o[119] ),
    .S(_05598_),
    .X(_03026_));
 sky130_fd_sc_hd__a22o_1 _14726_ (.A1(\sub1.data_o[87] ),
    .A2(_03010_),
    .B1(_03026_),
    .B2(\sub1.next_ready_o ),
    .X(_03027_));
 sky130_fd_sc_hd__a31o_1 _14727_ (.A1(_03019_),
    .A2(_04927_),
    .A3(_05245_),
    .B1(_03027_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _14728_ (.A0(net806),
    .A1(_05547_),
    .S(_04916_),
    .X(_03028_));
 sky130_fd_sc_hd__clkbuf_1 _14729_ (.A(_03028_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _14730_ (.A0(\ks1.col[1] ),
    .A1(_05553_),
    .S(_04916_),
    .X(_03029_));
 sky130_fd_sc_hd__clkbuf_1 _14731_ (.A(_03029_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _14732_ (.A0(\ks1.col[2] ),
    .A1(_05559_),
    .S(_04916_),
    .X(_03030_));
 sky130_fd_sc_hd__clkbuf_1 _14733_ (.A(_03030_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _14734_ (.A0(\ks1.col[3] ),
    .A1(_05172_),
    .S(_04916_),
    .X(_03031_));
 sky130_fd_sc_hd__clkbuf_1 _14735_ (.A(_03031_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _14736_ (.A0(\ks1.col[4] ),
    .A1(_05217_),
    .S(_04916_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_1 _14737_ (.A(_03032_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _14738_ (.A0(\ks1.col[5] ),
    .A1(_05225_),
    .S(_04916_),
    .X(_03033_));
 sky130_fd_sc_hd__clkbuf_1 _14739_ (.A(_03033_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _14740_ (.A0(\ks1.col[6] ),
    .A1(_05235_),
    .S(_04916_),
    .X(_03034_));
 sky130_fd_sc_hd__clkbuf_1 _14741_ (.A(_03034_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _14742_ (.A0(\ks1.col[7] ),
    .A1(_05244_),
    .S(_04916_),
    .X(_03035_));
 sky130_fd_sc_hd__clkbuf_1 _14743_ (.A(_03035_),
    .X(_01584_));
 sky130_fd_sc_hd__mux2_1 _14744_ (.A0(\ks1.col[24] ),
    .A1(_05547_),
    .S(_04911_),
    .X(_03036_));
 sky130_fd_sc_hd__clkbuf_1 _14745_ (.A(_03036_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _14746_ (.A0(\ks1.col[25] ),
    .A1(_05553_),
    .S(_04911_),
    .X(_03037_));
 sky130_fd_sc_hd__clkbuf_1 _14747_ (.A(_03037_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _14748_ (.A0(\ks1.col[26] ),
    .A1(_05559_),
    .S(_04911_),
    .X(_03038_));
 sky130_fd_sc_hd__clkbuf_1 _14749_ (.A(_03038_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _14750_ (.A0(\ks1.col[27] ),
    .A1(_05172_),
    .S(_04911_),
    .X(_03039_));
 sky130_fd_sc_hd__clkbuf_1 _14751_ (.A(_03039_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _14752_ (.A0(\ks1.col[28] ),
    .A1(_05217_),
    .S(_04911_),
    .X(_03040_));
 sky130_fd_sc_hd__clkbuf_1 _14753_ (.A(_03040_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _14754_ (.A0(\ks1.col[29] ),
    .A1(_05225_),
    .S(_04911_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_1 _14755_ (.A(_03041_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _14756_ (.A0(\ks1.col[30] ),
    .A1(_05235_),
    .S(_04911_),
    .X(_03042_));
 sky130_fd_sc_hd__clkbuf_1 _14757_ (.A(_03042_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _14758_ (.A0(\ks1.col[31] ),
    .A1(_05244_),
    .S(_04911_),
    .X(_03043_));
 sky130_fd_sc_hd__clkbuf_1 _14759_ (.A(_03043_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _14760_ (.A0(\ks1.col[16] ),
    .A1(_05547_),
    .S(_00007_),
    .X(_03044_));
 sky130_fd_sc_hd__clkbuf_1 _14761_ (.A(_03044_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _14762_ (.A0(\ks1.col[17] ),
    .A1(_05553_),
    .S(_00007_),
    .X(_03045_));
 sky130_fd_sc_hd__clkbuf_1 _14763_ (.A(_03045_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _14764_ (.A0(\ks1.col[18] ),
    .A1(_05559_),
    .S(_00007_),
    .X(_03046_));
 sky130_fd_sc_hd__clkbuf_1 _14765_ (.A(_03046_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _14766_ (.A0(\ks1.col[19] ),
    .A1(_05172_),
    .S(_00007_),
    .X(_03047_));
 sky130_fd_sc_hd__clkbuf_1 _14767_ (.A(_03047_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _14768_ (.A0(\ks1.col[20] ),
    .A1(_05217_),
    .S(_00007_),
    .X(_03048_));
 sky130_fd_sc_hd__clkbuf_1 _14769_ (.A(_03048_),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _14770_ (.A0(\ks1.col[21] ),
    .A1(_05225_),
    .S(_00007_),
    .X(_03049_));
 sky130_fd_sc_hd__clkbuf_1 _14771_ (.A(_03049_),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _14772_ (.A0(\ks1.col[22] ),
    .A1(_05235_),
    .S(_00007_),
    .X(_03050_));
 sky130_fd_sc_hd__clkbuf_1 _14773_ (.A(_03050_),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _14774_ (.A0(\ks1.col[23] ),
    .A1(_05244_),
    .S(_00007_),
    .X(_03051_));
 sky130_fd_sc_hd__clkbuf_1 _14775_ (.A(_03051_),
    .X(_01600_));
 sky130_fd_sc_hd__a22oi_1 _14776_ (.A1(_04617_),
    .A2(\sub1.ready_o ),
    .B1(_04666_),
    .B2(addroundkey_ready_o),
    .Y(_03052_));
 sky130_fd_sc_hd__a211o_1 _14777_ (.A1(state),
    .A2(_04622_),
    .B1(_03052_),
    .C1(\mix1.state[0] ),
    .X(_03053_));
 sky130_fd_sc_hd__nor2_4 _14778_ (.A(\mix1.state[1] ),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__buf_6 _14779_ (.A(_03054_),
    .X(_03055_));
 sky130_fd_sc_hd__clkbuf_8 _14780_ (.A(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__buf_6 _14781_ (.A(_03056_),
    .X(_03057_));
 sky130_fd_sc_hd__buf_4 _14782_ (.A(_04658_),
    .X(_03058_));
 sky130_fd_sc_hd__buf_4 _14783_ (.A(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__inv_2 _14784_ (.A(\mix1.state[1] ),
    .Y(_03060_));
 sky130_fd_sc_hd__and2_2 _14785_ (.A(\mix1.state[0] ),
    .B(_03060_),
    .X(_03061_));
 sky130_fd_sc_hd__buf_4 _14786_ (.A(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__clkbuf_4 _14787_ (.A(_03062_),
    .X(_03063_));
 sky130_fd_sc_hd__buf_4 _14788_ (.A(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__nor2_2 _14789_ (.A(\mix1.state[0] ),
    .B(_03060_),
    .Y(_03065_));
 sky130_fd_sc_hd__buf_4 _14790_ (.A(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__buf_4 _14791_ (.A(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__buf_4 _14792_ (.A(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__a22o_1 _14793_ (.A1(\sub1.data_o[80] ),
    .A2(_03064_),
    .B1(_03068_),
    .B2(\sub1.data_o[48] ),
    .X(_03069_));
 sky130_fd_sc_hd__a211o_1 _14794_ (.A1(\sub1.data_o[16] ),
    .A2(_04378_),
    .B1(_03059_),
    .C1(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__a21oi_1 _14795_ (.A1(\sub1.data_o[112] ),
    .A2(_03057_),
    .B1(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__buf_4 _14796_ (.A(_03064_),
    .X(_03072_));
 sky130_fd_sc_hd__a22o_1 _14797_ (.A1(\addroundkey_data_o[80] ),
    .A2(_03072_),
    .B1(_03068_),
    .B2(\addroundkey_data_o[48] ),
    .X(_03073_));
 sky130_fd_sc_hd__a211o_1 _14798_ (.A1(\addroundkey_data_o[16] ),
    .A2(_04378_),
    .B1(_05607_),
    .C1(_03073_),
    .X(_03074_));
 sky130_fd_sc_hd__a21oi_2 _14799_ (.A1(\addroundkey_data_o[112] ),
    .A2(_03057_),
    .B1(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__nor2_4 _14800_ (.A(_03071_),
    .B(_03075_),
    .Y(_03076_));
 sky130_fd_sc_hd__buf_6 _14801_ (.A(_03054_),
    .X(_03077_));
 sky130_fd_sc_hd__clkbuf_8 _14802_ (.A(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__buf_4 _14803_ (.A(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__a22o_1 _14804_ (.A1(\sub1.data_o[24] ),
    .A2(_04376_),
    .B1(_03067_),
    .B2(\sub1.data_o[56] ),
    .X(_03080_));
 sky130_fd_sc_hd__buf_4 _14805_ (.A(_03058_),
    .X(_03081_));
 sky130_fd_sc_hd__a211o_1 _14806_ (.A1(\sub1.data_o[88] ),
    .A2(_03072_),
    .B1(_03080_),
    .C1(_03081_),
    .X(_03082_));
 sky130_fd_sc_hd__a21oi_1 _14807_ (.A1(\sub1.data_o[120] ),
    .A2(_03079_),
    .B1(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__buf_4 _14808_ (.A(_03066_),
    .X(_03084_));
 sky130_fd_sc_hd__a22o_1 _14809_ (.A1(\addroundkey_data_o[24] ),
    .A2(_04376_),
    .B1(_03084_),
    .B2(\addroundkey_data_o[56] ),
    .X(_03085_));
 sky130_fd_sc_hd__clkbuf_4 _14810_ (.A(_05606_),
    .X(_03086_));
 sky130_fd_sc_hd__a211o_1 _14811_ (.A1(\addroundkey_data_o[88] ),
    .A2(_03072_),
    .B1(_03085_),
    .C1(_03086_),
    .X(_03087_));
 sky130_fd_sc_hd__a21oi_1 _14812_ (.A1(\addroundkey_data_o[120] ),
    .A2(_03079_),
    .B1(_03087_),
    .Y(_03088_));
 sky130_fd_sc_hd__nor2_4 _14813_ (.A(_03083_),
    .B(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__xnor2_4 _14814_ (.A(_03076_),
    .B(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__buf_4 _14815_ (.A(_03065_),
    .X(_03091_));
 sky130_fd_sc_hd__clkbuf_4 _14816_ (.A(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__a22o_1 _14817_ (.A1(\sub1.data_o[77] ),
    .A2(_03063_),
    .B1(_03092_),
    .B2(\sub1.data_o[45] ),
    .X(_03093_));
 sky130_fd_sc_hd__a211o_1 _14818_ (.A1(\sub1.data_o[13] ),
    .A2(_04376_),
    .B1(_03081_),
    .C1(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__a21oi_2 _14819_ (.A1(\sub1.data_o[109] ),
    .A2(_03078_),
    .B1(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a22o_1 _14820_ (.A1(\addroundkey_data_o[77] ),
    .A2(_03063_),
    .B1(_03092_),
    .B2(\addroundkey_data_o[45] ),
    .X(_03096_));
 sky130_fd_sc_hd__a211o_1 _14821_ (.A1(\addroundkey_data_o[13] ),
    .A2(_04376_),
    .B1(_05606_),
    .C1(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__a21oi_2 _14822_ (.A1(\addroundkey_data_o[109] ),
    .A2(_03078_),
    .B1(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__nor2_8 _14823_ (.A(_03095_),
    .B(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__buf_4 _14824_ (.A(_04375_),
    .X(_03100_));
 sky130_fd_sc_hd__a22o_1 _14825_ (.A1(\sub1.data_o[70] ),
    .A2(_03062_),
    .B1(_03091_),
    .B2(\sub1.data_o[38] ),
    .X(_03101_));
 sky130_fd_sc_hd__a211o_1 _14826_ (.A1(\sub1.data_o[6] ),
    .A2(_03100_),
    .B1(_03058_),
    .C1(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__a21oi_4 _14827_ (.A1(\sub1.data_o[102] ),
    .A2(_03055_),
    .B1(_03102_),
    .Y(_03103_));
 sky130_fd_sc_hd__a22o_1 _14828_ (.A1(\addroundkey_data_o[70] ),
    .A2(_03062_),
    .B1(_03091_),
    .B2(\addroundkey_data_o[38] ),
    .X(_03104_));
 sky130_fd_sc_hd__a211o_1 _14829_ (.A1(\addroundkey_data_o[6] ),
    .A2(_03100_),
    .B1(_05606_),
    .C1(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__a21oi_4 _14830_ (.A1(\addroundkey_data_o[102] ),
    .A2(_03077_),
    .B1(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__nor2_8 _14831_ (.A(_03103_),
    .B(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__buf_4 _14832_ (.A(_03061_),
    .X(_03108_));
 sky130_fd_sc_hd__a22o_1 _14833_ (.A1(\sub1.data_o[85] ),
    .A2(_03108_),
    .B1(_03066_),
    .B2(\sub1.data_o[53] ),
    .X(_03109_));
 sky130_fd_sc_hd__a211o_1 _14834_ (.A1(\sub1.data_o[21] ),
    .A2(_03100_),
    .B1(_03058_),
    .C1(_03109_),
    .X(_03110_));
 sky130_fd_sc_hd__a21oi_1 _14835_ (.A1(\sub1.data_o[117] ),
    .A2(_03055_),
    .B1(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__a22o_1 _14836_ (.A1(\addroundkey_data_o[85] ),
    .A2(_03108_),
    .B1(_03066_),
    .B2(\addroundkey_data_o[53] ),
    .X(_03112_));
 sky130_fd_sc_hd__a211o_1 _14837_ (.A1(\addroundkey_data_o[21] ),
    .A2(_04376_),
    .B1(_05606_),
    .C1(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__a21oi_2 _14838_ (.A1(\addroundkey_data_o[117] ),
    .A2(_03055_),
    .B1(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__nor2_4 _14839_ (.A(_03111_),
    .B(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__xor2_2 _14840_ (.A(_03107_),
    .B(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__xnor2_4 _14841_ (.A(_03099_),
    .B(_03116_),
    .Y(_03117_));
 sky130_fd_sc_hd__a22o_1 _14842_ (.A1(\sub1.data_o[86] ),
    .A2(_03062_),
    .B1(_03091_),
    .B2(\sub1.data_o[54] ),
    .X(_03118_));
 sky130_fd_sc_hd__a211o_1 _14843_ (.A1(\sub1.data_o[22] ),
    .A2(_03100_),
    .B1(_03058_),
    .C1(_03118_),
    .X(_03119_));
 sky130_fd_sc_hd__a21oi_2 _14844_ (.A1(\sub1.data_o[118] ),
    .A2(_03077_),
    .B1(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__a22o_1 _14845_ (.A1(\addroundkey_data_o[86] ),
    .A2(_03062_),
    .B1(_03091_),
    .B2(\addroundkey_data_o[54] ),
    .X(_03121_));
 sky130_fd_sc_hd__a211o_1 _14846_ (.A1(\addroundkey_data_o[22] ),
    .A2(_04375_),
    .B1(_04900_),
    .C1(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__a21oi_2 _14847_ (.A1(\addroundkey_data_o[118] ),
    .A2(_03077_),
    .B1(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__nor2_8 _14848_ (.A(_03120_),
    .B(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__a22o_1 _14849_ (.A1(\sub1.data_o[69] ),
    .A2(_03108_),
    .B1(_03066_),
    .B2(\sub1.data_o[37] ),
    .X(_03125_));
 sky130_fd_sc_hd__a211o_1 _14850_ (.A1(\sub1.data_o[5] ),
    .A2(_03100_),
    .B1(_03058_),
    .C1(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__a21oi_4 _14851_ (.A1(\sub1.data_o[101] ),
    .A2(_03055_),
    .B1(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__a22o_1 _14852_ (.A1(\addroundkey_data_o[69] ),
    .A2(_03108_),
    .B1(_03066_),
    .B2(\addroundkey_data_o[37] ),
    .X(_03128_));
 sky130_fd_sc_hd__a211o_1 _14853_ (.A1(\addroundkey_data_o[5] ),
    .A2(_03100_),
    .B1(_05606_),
    .C1(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__a21oi_4 _14854_ (.A1(\addroundkey_data_o[101] ),
    .A2(_03055_),
    .B1(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__nor2_8 _14855_ (.A(_03127_),
    .B(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__a22o_1 _14856_ (.A1(\sub1.data_o[93] ),
    .A2(_03108_),
    .B1(_03066_),
    .B2(\sub1.data_o[61] ),
    .X(_03132_));
 sky130_fd_sc_hd__a211o_1 _14857_ (.A1(\sub1.data_o[29] ),
    .A2(_03100_),
    .B1(_03058_),
    .C1(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__a21oi_2 _14858_ (.A1(\sub1.data_o[125] ),
    .A2(_03055_),
    .B1(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__a22o_1 _14859_ (.A1(\addroundkey_data_o[93] ),
    .A2(_03108_),
    .B1(_03066_),
    .B2(\addroundkey_data_o[61] ),
    .X(_03135_));
 sky130_fd_sc_hd__a211o_1 _14860_ (.A1(\addroundkey_data_o[29] ),
    .A2(_03100_),
    .B1(_05606_),
    .C1(_03135_),
    .X(_03136_));
 sky130_fd_sc_hd__a21oi_2 _14861_ (.A1(\addroundkey_data_o[125] ),
    .A2(_03055_),
    .B1(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__nor2_8 _14862_ (.A(_03134_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__xnor2_4 _14863_ (.A(_03131_),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__xnor2_4 _14864_ (.A(_03124_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__xor2_4 _14865_ (.A(_03117_),
    .B(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__or2_1 _14866_ (.A(_04617_),
    .B(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__buf_8 _14867_ (.A(_03057_),
    .X(_03143_));
 sky130_fd_sc_hd__buf_6 _14868_ (.A(_03072_),
    .X(_03144_));
 sky130_fd_sc_hd__buf_6 _14869_ (.A(_03068_),
    .X(_03145_));
 sky130_fd_sc_hd__a22o_1 _14870_ (.A1(\sub1.data_o[72] ),
    .A2(_03144_),
    .B1(_03145_),
    .B2(\sub1.data_o[40] ),
    .X(_03146_));
 sky130_fd_sc_hd__a211o_1 _14871_ (.A1(\sub1.data_o[8] ),
    .A2(_04379_),
    .B1(_03059_),
    .C1(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__a21oi_2 _14872_ (.A1(\sub1.data_o[104] ),
    .A2(_03143_),
    .B1(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__a22o_1 _14873_ (.A1(\addroundkey_data_o[72] ),
    .A2(_03144_),
    .B1(_03145_),
    .B2(\addroundkey_data_o[40] ),
    .X(_03149_));
 sky130_fd_sc_hd__a211o_1 _14874_ (.A1(\addroundkey_data_o[8] ),
    .A2(_04379_),
    .B1(_05607_),
    .C1(_03149_),
    .X(_03150_));
 sky130_fd_sc_hd__a21oi_2 _14875_ (.A1(\addroundkey_data_o[104] ),
    .A2(_03143_),
    .B1(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__nor2_8 _14876_ (.A(_03148_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__xnor2_2 _14877_ (.A(_03142_),
    .B(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__a22o_1 _14878_ (.A1(\sub1.data_o[71] ),
    .A2(_03061_),
    .B1(_03065_),
    .B2(\sub1.data_o[39] ),
    .X(_03154_));
 sky130_fd_sc_hd__a211o_1 _14879_ (.A1(\sub1.data_o[7] ),
    .A2(_04374_),
    .B1(_04658_),
    .C1(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__a21oi_2 _14880_ (.A1(\sub1.data_o[103] ),
    .A2(_03054_),
    .B1(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__a22o_1 _14881_ (.A1(\addroundkey_data_o[71] ),
    .A2(_03061_),
    .B1(_03065_),
    .B2(\addroundkey_data_o[39] ),
    .X(_03157_));
 sky130_fd_sc_hd__a211o_1 _14882_ (.A1(\addroundkey_data_o[7] ),
    .A2(_04374_),
    .B1(_04900_),
    .C1(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__a21oi_4 _14883_ (.A1(\addroundkey_data_o[103] ),
    .A2(_03054_),
    .B1(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hd__nor2_8 _14884_ (.A(_03156_),
    .B(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__a22o_1 _14885_ (.A1(\sub1.data_o[95] ),
    .A2(_03061_),
    .B1(_03065_),
    .B2(\sub1.data_o[63] ),
    .X(_03161_));
 sky130_fd_sc_hd__a211o_1 _14886_ (.A1(\sub1.data_o[31] ),
    .A2(_04374_),
    .B1(_04658_),
    .C1(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__a21oi_2 _14887_ (.A1(\sub1.data_o[127] ),
    .A2(_03054_),
    .B1(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__a22o_1 _14888_ (.A1(\addroundkey_data_o[95] ),
    .A2(_03061_),
    .B1(_03065_),
    .B2(\addroundkey_data_o[63] ),
    .X(_03164_));
 sky130_fd_sc_hd__a211o_1 _14889_ (.A1(\addroundkey_data_o[31] ),
    .A2(_04375_),
    .B1(_04900_),
    .C1(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__a21oi_2 _14890_ (.A1(\addroundkey_data_o[127] ),
    .A2(_03054_),
    .B1(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__nor2_8 _14891_ (.A(_03163_),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__xnor2_4 _14892_ (.A(_03160_),
    .B(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__xnor2_1 _14893_ (.A(_03153_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__xnor2_2 _14894_ (.A(_03090_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__buf_4 _14895_ (.A(_03144_),
    .X(_03171_));
 sky130_fd_sc_hd__mux2_1 _14896_ (.A0(\mix1.data_reg[64] ),
    .A1(_03170_),
    .S(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__clkbuf_1 _14897_ (.A(_03172_),
    .X(_01601_));
 sky130_fd_sc_hd__a22o_1 _14898_ (.A1(\sub1.data_o[94] ),
    .A2(_03063_),
    .B1(_03092_),
    .B2(\sub1.data_o[62] ),
    .X(_03173_));
 sky130_fd_sc_hd__a211o_1 _14899_ (.A1(\sub1.data_o[30] ),
    .A2(_04376_),
    .B1(_03081_),
    .C1(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__a21oi_2 _14900_ (.A1(\sub1.data_o[126] ),
    .A2(_03078_),
    .B1(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__a22o_1 _14901_ (.A1(\addroundkey_data_o[94] ),
    .A2(_03063_),
    .B1(_03092_),
    .B2(\addroundkey_data_o[62] ),
    .X(_03176_));
 sky130_fd_sc_hd__a211o_1 _14902_ (.A1(\addroundkey_data_o[30] ),
    .A2(_04377_),
    .B1(_05606_),
    .C1(_03176_),
    .X(_03177_));
 sky130_fd_sc_hd__a21oi_2 _14903_ (.A1(\addroundkey_data_o[126] ),
    .A2(_03078_),
    .B1(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__nor2_8 _14904_ (.A(_03175_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__xnor2_4 _14905_ (.A(_03107_),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__a22o_1 _14906_ (.A1(\sub1.data_o[87] ),
    .A2(_03062_),
    .B1(_03091_),
    .B2(\sub1.data_o[55] ),
    .X(_03181_));
 sky130_fd_sc_hd__a211o_1 _14907_ (.A1(\sub1.data_o[23] ),
    .A2(_04375_),
    .B1(_03058_),
    .C1(_03181_),
    .X(_03182_));
 sky130_fd_sc_hd__a21oi_2 _14908_ (.A1(\sub1.data_o[119] ),
    .A2(_03077_),
    .B1(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__a22o_1 _14909_ (.A1(\addroundkey_data_o[87] ),
    .A2(_03062_),
    .B1(_03091_),
    .B2(\addroundkey_data_o[55] ),
    .X(_03184_));
 sky130_fd_sc_hd__a211o_1 _14910_ (.A1(\addroundkey_data_o[23] ),
    .A2(_04375_),
    .B1(_04900_),
    .C1(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__a21oi_2 _14911_ (.A1(\addroundkey_data_o[119] ),
    .A2(_03077_),
    .B1(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__nor2_8 _14912_ (.A(_03183_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__xnor2_2 _14913_ (.A(_03160_),
    .B(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__a22o_1 _14914_ (.A1(\sub1.data_o[78] ),
    .A2(_03108_),
    .B1(_03066_),
    .B2(\sub1.data_o[46] ),
    .X(_03189_));
 sky130_fd_sc_hd__a211o_1 _14915_ (.A1(\sub1.data_o[14] ),
    .A2(_03100_),
    .B1(_03058_),
    .C1(_03189_),
    .X(_03190_));
 sky130_fd_sc_hd__a21oi_2 _14916_ (.A1(\sub1.data_o[110] ),
    .A2(_03055_),
    .B1(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__a22o_1 _14917_ (.A1(\addroundkey_data_o[78] ),
    .A2(_03108_),
    .B1(_03066_),
    .B2(\addroundkey_data_o[46] ),
    .X(_03192_));
 sky130_fd_sc_hd__a211o_1 _14918_ (.A1(\addroundkey_data_o[14] ),
    .A2(_03100_),
    .B1(_05606_),
    .C1(_03192_),
    .X(_03193_));
 sky130_fd_sc_hd__a21oi_2 _14919_ (.A1(\addroundkey_data_o[110] ),
    .A2(_03055_),
    .B1(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__nor2_8 _14920_ (.A(_03191_),
    .B(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__xnor2_4 _14921_ (.A(_03124_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__xor2_2 _14922_ (.A(_03188_),
    .B(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__xnor2_4 _14923_ (.A(_03180_),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__xnor2_2 _14924_ (.A(_03141_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__nand2_2 _14925_ (.A(_05201_),
    .B(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__a22o_1 _14926_ (.A1(\sub1.data_o[89] ),
    .A2(_03063_),
    .B1(_03092_),
    .B2(\sub1.data_o[57] ),
    .X(_03201_));
 sky130_fd_sc_hd__a211o_1 _14927_ (.A1(\sub1.data_o[25] ),
    .A2(_04377_),
    .B1(_03081_),
    .C1(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__a21oi_2 _14928_ (.A1(\sub1.data_o[121] ),
    .A2(_03056_),
    .B1(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__a22o_1 _14929_ (.A1(\addroundkey_data_o[89] ),
    .A2(_03063_),
    .B1(_03092_),
    .B2(\addroundkey_data_o[57] ),
    .X(_03204_));
 sky130_fd_sc_hd__a211o_1 _14930_ (.A1(\addroundkey_data_o[25] ),
    .A2(_04377_),
    .B1(_03086_),
    .C1(_03204_),
    .X(_03205_));
 sky130_fd_sc_hd__a21oi_2 _14931_ (.A1(\addroundkey_data_o[121] ),
    .A2(_03078_),
    .B1(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__nor2_8 _14932_ (.A(_03203_),
    .B(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__buf_4 _14933_ (.A(_04376_),
    .X(_03208_));
 sky130_fd_sc_hd__buf_4 _14934_ (.A(_03108_),
    .X(_03209_));
 sky130_fd_sc_hd__a22o_1 _14935_ (.A1(\sub1.data_o[64] ),
    .A2(_03209_),
    .B1(_03067_),
    .B2(\sub1.data_o[32] ),
    .X(_03210_));
 sky130_fd_sc_hd__a211o_1 _14936_ (.A1(\sub1.data_o[0] ),
    .A2(_03208_),
    .B1(_03081_),
    .C1(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__a21oi_1 _14937_ (.A1(\sub1.data_o[96] ),
    .A2(_03056_),
    .B1(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__a22o_1 _14938_ (.A1(\addroundkey_data_o[64] ),
    .A2(_03209_),
    .B1(_03067_),
    .B2(\addroundkey_data_o[32] ),
    .X(_03213_));
 sky130_fd_sc_hd__a211o_1 _14939_ (.A1(\addroundkey_data_o[0] ),
    .A2(_03208_),
    .B1(_03086_),
    .C1(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__a21oi_2 _14940_ (.A1(\addroundkey_data_o[96] ),
    .A2(_03056_),
    .B1(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__nor2_4 _14941_ (.A(_03212_),
    .B(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__xnor2_2 _14942_ (.A(_03089_),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__xor2_2 _14943_ (.A(_03168_),
    .B(_03217_),
    .X(_03218_));
 sky130_fd_sc_hd__a22o_1 _14944_ (.A1(\sub1.data_o[73] ),
    .A2(_03063_),
    .B1(_03092_),
    .B2(\sub1.data_o[41] ),
    .X(_03219_));
 sky130_fd_sc_hd__a211o_1 _14945_ (.A1(\sub1.data_o[9] ),
    .A2(_04377_),
    .B1(_03081_),
    .C1(_03219_),
    .X(_03220_));
 sky130_fd_sc_hd__a21oi_2 _14946_ (.A1(\sub1.data_o[105] ),
    .A2(_03078_),
    .B1(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__a22o_1 _14947_ (.A1(\addroundkey_data_o[73] ),
    .A2(_03063_),
    .B1(_03092_),
    .B2(\addroundkey_data_o[41] ),
    .X(_03222_));
 sky130_fd_sc_hd__a211o_1 _14948_ (.A1(\addroundkey_data_o[9] ),
    .A2(_04377_),
    .B1(_03086_),
    .C1(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__a21oi_4 _14949_ (.A1(\addroundkey_data_o[105] ),
    .A2(_03078_),
    .B1(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__nor2_8 _14950_ (.A(_03221_),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hd__a22o_1 _14951_ (.A1(\sub1.data_o[81] ),
    .A2(_03209_),
    .B1(_03067_),
    .B2(\sub1.data_o[49] ),
    .X(_03226_));
 sky130_fd_sc_hd__a211o_1 _14952_ (.A1(\sub1.data_o[17] ),
    .A2(_04377_),
    .B1(_03081_),
    .C1(_03226_),
    .X(_03227_));
 sky130_fd_sc_hd__a21oi_1 _14953_ (.A1(\sub1.data_o[113] ),
    .A2(_03056_),
    .B1(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__a22o_1 _14954_ (.A1(\addroundkey_data_o[81] ),
    .A2(_03209_),
    .B1(_03067_),
    .B2(\addroundkey_data_o[49] ),
    .X(_03229_));
 sky130_fd_sc_hd__a211o_1 _14955_ (.A1(\addroundkey_data_o[17] ),
    .A2(_04377_),
    .B1(_03086_),
    .C1(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__a21oi_2 _14956_ (.A1(\addroundkey_data_o[113] ),
    .A2(_03056_),
    .B1(_03230_),
    .Y(_03231_));
 sky130_fd_sc_hd__nor2_4 _14957_ (.A(_03228_),
    .B(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__xnor2_4 _14958_ (.A(_03225_),
    .B(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__xor2_1 _14959_ (.A(_03218_),
    .B(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__xnor2_1 _14960_ (.A(_03207_),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__xnor2_2 _14961_ (.A(_03200_),
    .B(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__mux2_1 _14962_ (.A0(\mix1.data_reg[65] ),
    .A1(_03236_),
    .S(_03171_),
    .X(_03237_));
 sky130_fd_sc_hd__clkbuf_1 _14963_ (.A(_03237_),
    .X(_01602_));
 sky130_fd_sc_hd__xnor2_1 _14964_ (.A(_03168_),
    .B(_03216_),
    .Y(_03238_));
 sky130_fd_sc_hd__a22o_1 _14965_ (.A1(\sub1.data_o[79] ),
    .A2(_03063_),
    .B1(_03092_),
    .B2(\sub1.data_o[47] ),
    .X(_03239_));
 sky130_fd_sc_hd__a211o_1 _14966_ (.A1(\sub1.data_o[15] ),
    .A2(_04376_),
    .B1(_03058_),
    .C1(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__a21oi_2 _14967_ (.A1(\sub1.data_o[111] ),
    .A2(_03078_),
    .B1(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__a22o_1 _14968_ (.A1(\addroundkey_data_o[79] ),
    .A2(_03108_),
    .B1(_03092_),
    .B2(\addroundkey_data_o[47] ),
    .X(_03242_));
 sky130_fd_sc_hd__a211o_1 _14969_ (.A1(\addroundkey_data_o[15] ),
    .A2(_04376_),
    .B1(_05606_),
    .C1(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__a21oi_2 _14970_ (.A1(\addroundkey_data_o[111] ),
    .A2(_03078_),
    .B1(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__nor2_8 _14971_ (.A(_03241_),
    .B(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__xnor2_4 _14972_ (.A(_03187_),
    .B(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__xor2_4 _14973_ (.A(_03076_),
    .B(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__xnor2_1 _14974_ (.A(_03238_),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__o21ai_1 _14975_ (.A1(_03198_),
    .A2(_03248_),
    .B1(_05201_),
    .Y(_03249_));
 sky130_fd_sc_hd__a21oi_2 _14976_ (.A1(_03198_),
    .A2(_03248_),
    .B1(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__a22o_1 _14977_ (.A1(\sub1.data_o[74] ),
    .A2(_03209_),
    .B1(_03067_),
    .B2(\sub1.data_o[42] ),
    .X(_03251_));
 sky130_fd_sc_hd__a211o_1 _14978_ (.A1(\sub1.data_o[10] ),
    .A2(_04377_),
    .B1(_03081_),
    .C1(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__a21oi_1 _14979_ (.A1(\sub1.data_o[106] ),
    .A2(_03056_),
    .B1(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__a22o_1 _14980_ (.A1(\addroundkey_data_o[74] ),
    .A2(_03209_),
    .B1(_03067_),
    .B2(\addroundkey_data_o[42] ),
    .X(_03254_));
 sky130_fd_sc_hd__a211o_1 _14981_ (.A1(\addroundkey_data_o[10] ),
    .A2(_04377_),
    .B1(_03086_),
    .C1(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__a21oi_1 _14982_ (.A1(\addroundkey_data_o[106] ),
    .A2(_03056_),
    .B1(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__nor2_4 _14983_ (.A(_03253_),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__a22o_1 _14984_ (.A1(\sub1.data_o[90] ),
    .A2(_03061_),
    .B1(_03065_),
    .B2(\sub1.data_o[58] ),
    .X(_03258_));
 sky130_fd_sc_hd__a211o_1 _14985_ (.A1(\sub1.data_o[26] ),
    .A2(_04375_),
    .B1(_04658_),
    .C1(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__a21oi_1 _14986_ (.A1(\sub1.data_o[122] ),
    .A2(_03077_),
    .B1(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__a22o_1 _14987_ (.A1(\addroundkey_data_o[90] ),
    .A2(_03062_),
    .B1(_03091_),
    .B2(\addroundkey_data_o[58] ),
    .X(_03261_));
 sky130_fd_sc_hd__a211o_1 _14988_ (.A1(\addroundkey_data_o[26] ),
    .A2(_04375_),
    .B1(_04900_),
    .C1(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__a21oi_1 _14989_ (.A1(\addroundkey_data_o[122] ),
    .A2(_03077_),
    .B1(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__nor2_4 _14990_ (.A(_03260_),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__xnor2_4 _14991_ (.A(_03257_),
    .B(_03264_),
    .Y(_03265_));
 sky130_fd_sc_hd__xnor2_4 _14992_ (.A(_03250_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__a22o_1 _14993_ (.A1(\sub1.data_o[82] ),
    .A2(_03064_),
    .B1(_03084_),
    .B2(\sub1.data_o[50] ),
    .X(_03267_));
 sky130_fd_sc_hd__a211o_1 _14994_ (.A1(\sub1.data_o[18] ),
    .A2(_03208_),
    .B1(_03059_),
    .C1(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__a21oi_1 _14995_ (.A1(\sub1.data_o[114] ),
    .A2(_03079_),
    .B1(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__a22o_1 _14996_ (.A1(\addroundkey_data_o[82] ),
    .A2(_03064_),
    .B1(_03084_),
    .B2(\addroundkey_data_o[50] ),
    .X(_03270_));
 sky130_fd_sc_hd__a211o_1 _14997_ (.A1(\addroundkey_data_o[18] ),
    .A2(_03208_),
    .B1(_03086_),
    .C1(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__a21oi_2 _14998_ (.A1(\addroundkey_data_o[114] ),
    .A2(_03079_),
    .B1(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__nor2_4 _14999_ (.A(_03269_),
    .B(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__a22o_1 _15000_ (.A1(\sub1.data_o[65] ),
    .A2(_03209_),
    .B1(_03067_),
    .B2(\sub1.data_o[33] ),
    .X(_03274_));
 sky130_fd_sc_hd__a211o_1 _15001_ (.A1(\sub1.data_o[1] ),
    .A2(_03208_),
    .B1(_03081_),
    .C1(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__a21oi_2 _15002_ (.A1(\sub1.data_o[97] ),
    .A2(_03056_),
    .B1(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__a22o_1 _15003_ (.A1(\addroundkey_data_o[65] ),
    .A2(_03209_),
    .B1(_03067_),
    .B2(\addroundkey_data_o[33] ),
    .X(_03277_));
 sky130_fd_sc_hd__a211o_1 _15004_ (.A1(\addroundkey_data_o[1] ),
    .A2(_03208_),
    .B1(_03086_),
    .C1(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__a21oi_2 _15005_ (.A1(\addroundkey_data_o[97] ),
    .A2(_03056_),
    .B1(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__nor2_8 _15006_ (.A(_03276_),
    .B(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__xnor2_4 _15007_ (.A(_03207_),
    .B(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__xor2_4 _15008_ (.A(_03273_),
    .B(_03281_),
    .X(_03282_));
 sky130_fd_sc_hd__xnor2_4 _15009_ (.A(_03266_),
    .B(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__mux2_1 _15010_ (.A0(\mix1.data_reg[66] ),
    .A1(_03283_),
    .S(_03171_),
    .X(_03284_));
 sky130_fd_sc_hd__clkbuf_1 _15011_ (.A(_03284_),
    .X(_01603_));
 sky130_fd_sc_hd__xnor2_4 _15012_ (.A(_03232_),
    .B(_03280_),
    .Y(_03285_));
 sky130_fd_sc_hd__xnor2_1 _15013_ (.A(_03218_),
    .B(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hd__xnor2_2 _15014_ (.A(_03141_),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__xnor2_4 _15015_ (.A(_03152_),
    .B(_03247_),
    .Y(_03288_));
 sky130_fd_sc_hd__a21oi_1 _15016_ (.A1(_03287_),
    .A2(_03288_),
    .B1(_05198_),
    .Y(_03289_));
 sky130_fd_sc_hd__o21ai_4 _15017_ (.A1(_03287_),
    .A2(_03288_),
    .B1(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__a22o_1 _15018_ (.A1(\sub1.data_o[83] ),
    .A2(_03209_),
    .B1(_03084_),
    .B2(\sub1.data_o[51] ),
    .X(_03291_));
 sky130_fd_sc_hd__a211o_1 _15019_ (.A1(\sub1.data_o[19] ),
    .A2(_03208_),
    .B1(_03081_),
    .C1(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__a21oi_1 _15020_ (.A1(\sub1.data_o[115] ),
    .A2(_03079_),
    .B1(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__a22o_1 _15021_ (.A1(\addroundkey_data_o[83] ),
    .A2(_03209_),
    .B1(_03084_),
    .B2(\addroundkey_data_o[51] ),
    .X(_03294_));
 sky130_fd_sc_hd__a211o_1 _15022_ (.A1(\addroundkey_data_o[19] ),
    .A2(_03208_),
    .B1(_03086_),
    .C1(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__a21oi_2 _15023_ (.A1(\addroundkey_data_o[115] ),
    .A2(_03079_),
    .B1(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__nor2_4 _15024_ (.A(_03293_),
    .B(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__a22o_1 _15025_ (.A1(\sub1.data_o[66] ),
    .A2(_03062_),
    .B1(_03091_),
    .B2(\sub1.data_o[34] ),
    .X(_03298_));
 sky130_fd_sc_hd__a211o_1 _15026_ (.A1(\sub1.data_o[2] ),
    .A2(_04375_),
    .B1(_04658_),
    .C1(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__a21oi_2 _15027_ (.A1(\sub1.data_o[98] ),
    .A2(_03077_),
    .B1(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__a22o_1 _15028_ (.A1(\addroundkey_data_o[66] ),
    .A2(_03062_),
    .B1(_03091_),
    .B2(\addroundkey_data_o[34] ),
    .X(_03301_));
 sky130_fd_sc_hd__a211o_1 _15029_ (.A1(\addroundkey_data_o[2] ),
    .A2(_04375_),
    .B1(_04900_),
    .C1(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__a21oi_4 _15030_ (.A1(\addroundkey_data_o[98] ),
    .A2(_03077_),
    .B1(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__nor2_8 _15031_ (.A(_03300_),
    .B(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__xnor2_2 _15032_ (.A(_03264_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__xnor2_2 _15033_ (.A(_03168_),
    .B(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__xnor2_2 _15034_ (.A(_03297_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__a22o_1 _15035_ (.A1(\sub1.data_o[91] ),
    .A2(_03064_),
    .B1(_03068_),
    .B2(\sub1.data_o[59] ),
    .X(_03308_));
 sky130_fd_sc_hd__a211o_1 _15036_ (.A1(\sub1.data_o[27] ),
    .A2(_04378_),
    .B1(_03059_),
    .C1(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__a21oi_4 _15037_ (.A1(\sub1.data_o[123] ),
    .A2(_03057_),
    .B1(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__a22o_1 _15038_ (.A1(\addroundkey_data_o[91] ),
    .A2(_03064_),
    .B1(_03084_),
    .B2(\addroundkey_data_o[59] ),
    .X(_03311_));
 sky130_fd_sc_hd__a211o_1 _15039_ (.A1(\addroundkey_data_o[27] ),
    .A2(_04378_),
    .B1(_05607_),
    .C1(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__a21oi_2 _15040_ (.A1(\addroundkey_data_o[123] ),
    .A2(_03057_),
    .B1(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__nor2_8 _15041_ (.A(_03310_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__a22o_1 _15042_ (.A1(\sub1.data_o[75] ),
    .A2(_03064_),
    .B1(_03084_),
    .B2(\sub1.data_o[43] ),
    .X(_03315_));
 sky130_fd_sc_hd__a211o_1 _15043_ (.A1(\sub1.data_o[11] ),
    .A2(_03208_),
    .B1(_03059_),
    .C1(_03315_),
    .X(_03316_));
 sky130_fd_sc_hd__a21oi_2 _15044_ (.A1(\sub1.data_o[107] ),
    .A2(_03079_),
    .B1(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__a22o_1 _15045_ (.A1(\addroundkey_data_o[75] ),
    .A2(_03064_),
    .B1(_03084_),
    .B2(\addroundkey_data_o[43] ),
    .X(_03318_));
 sky130_fd_sc_hd__a211o_1 _15046_ (.A1(\addroundkey_data_o[11] ),
    .A2(_03208_),
    .B1(_03086_),
    .C1(_03318_),
    .X(_03319_));
 sky130_fd_sc_hd__a21oi_2 _15047_ (.A1(\addroundkey_data_o[107] ),
    .A2(_03079_),
    .B1(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__nor2_8 _15048_ (.A(_03317_),
    .B(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor2_2 _15049_ (.A(_03314_),
    .B(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__xnor2_2 _15050_ (.A(_03307_),
    .B(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__xnor2_4 _15051_ (.A(_03290_),
    .B(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__mux2_1 _15052_ (.A0(\mix1.data_reg[67] ),
    .A1(_03324_),
    .S(_03171_),
    .X(_03325_));
 sky130_fd_sc_hd__clkbuf_1 _15053_ (.A(_03325_),
    .X(_01604_));
 sky130_fd_sc_hd__xnor2_2 _15054_ (.A(_03233_),
    .B(_03304_),
    .Y(_03326_));
 sky130_fd_sc_hd__xnor2_1 _15055_ (.A(_03282_),
    .B(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__o21ai_1 _15056_ (.A1(_03199_),
    .A2(_03327_),
    .B1(_04624_),
    .Y(_03328_));
 sky130_fd_sc_hd__a21o_1 _15057_ (.A1(_03199_),
    .A2(_03327_),
    .B1(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__a22o_1 _15058_ (.A1(\sub1.data_o[92] ),
    .A2(_03144_),
    .B1(_03145_),
    .B2(\sub1.data_o[60] ),
    .X(_03330_));
 sky130_fd_sc_hd__a211o_1 _15059_ (.A1(\sub1.data_o[28] ),
    .A2(_04379_),
    .B1(_03059_),
    .C1(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__a21oi_4 _15060_ (.A1(\sub1.data_o[124] ),
    .A2(_03143_),
    .B1(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__a22o_1 _15061_ (.A1(\addroundkey_data_o[92] ),
    .A2(_03144_),
    .B1(_03145_),
    .B2(\addroundkey_data_o[60] ),
    .X(_03333_));
 sky130_fd_sc_hd__a211o_1 _15062_ (.A1(\addroundkey_data_o[28] ),
    .A2(_04379_),
    .B1(_05607_),
    .C1(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__a21oi_2 _15063_ (.A1(\addroundkey_data_o[124] ),
    .A2(_03143_),
    .B1(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__nor2_8 _15064_ (.A(_03332_),
    .B(_03335_),
    .Y(_03336_));
 sky130_fd_sc_hd__a22o_1 _15065_ (.A1(\sub1.data_o[84] ),
    .A2(_03072_),
    .B1(_03068_),
    .B2(\sub1.data_o[52] ),
    .X(_03337_));
 sky130_fd_sc_hd__a211o_1 _15066_ (.A1(\sub1.data_o[20] ),
    .A2(_04378_),
    .B1(_03059_),
    .C1(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__a21oi_2 _15067_ (.A1(\sub1.data_o[116] ),
    .A2(_03057_),
    .B1(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__a22o_1 _15068_ (.A1(\addroundkey_data_o[84] ),
    .A2(_03072_),
    .B1(_03068_),
    .B2(\addroundkey_data_o[52] ),
    .X(_03340_));
 sky130_fd_sc_hd__a211o_1 _15069_ (.A1(\addroundkey_data_o[20] ),
    .A2(_04379_),
    .B1(_05607_),
    .C1(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__a21oi_4 _15070_ (.A1(\addroundkey_data_o[116] ),
    .A2(_03057_),
    .B1(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__nor2_8 _15071_ (.A(_03339_),
    .B(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__xnor2_4 _15072_ (.A(_03336_),
    .B(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__xnor2_2 _15073_ (.A(_03329_),
    .B(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__a22o_1 _15074_ (.A1(\sub1.data_o[67] ),
    .A2(_03064_),
    .B1(_03084_),
    .B2(\sub1.data_o[35] ),
    .X(_03346_));
 sky130_fd_sc_hd__a211o_1 _15075_ (.A1(\sub1.data_o[3] ),
    .A2(_04378_),
    .B1(_03059_),
    .C1(_03346_),
    .X(_03347_));
 sky130_fd_sc_hd__a21oi_1 _15076_ (.A1(\sub1.data_o[99] ),
    .A2(_03079_),
    .B1(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__a22o_1 _15077_ (.A1(\addroundkey_data_o[67] ),
    .A2(_03064_),
    .B1(_03084_),
    .B2(\addroundkey_data_o[35] ),
    .X(_03349_));
 sky130_fd_sc_hd__a211o_1 _15078_ (.A1(\addroundkey_data_o[3] ),
    .A2(_04378_),
    .B1(_05607_),
    .C1(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__a21oi_2 _15079_ (.A1(\addroundkey_data_o[99] ),
    .A2(_03079_),
    .B1(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__nor2_4 _15080_ (.A(_03348_),
    .B(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__xnor2_4 _15081_ (.A(_03314_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__xnor2_2 _15082_ (.A(_03168_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__a22o_1 _15083_ (.A1(\sub1.data_o[76] ),
    .A2(_03072_),
    .B1(_03068_),
    .B2(\sub1.data_o[44] ),
    .X(_03355_));
 sky130_fd_sc_hd__a211o_1 _15084_ (.A1(\sub1.data_o[12] ),
    .A2(_04378_),
    .B1(_03059_),
    .C1(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__a21oi_2 _15085_ (.A1(\sub1.data_o[108] ),
    .A2(_03057_),
    .B1(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__a22o_1 _15086_ (.A1(\addroundkey_data_o[76] ),
    .A2(_03072_),
    .B1(_03068_),
    .B2(\addroundkey_data_o[44] ),
    .X(_03358_));
 sky130_fd_sc_hd__a211o_1 _15087_ (.A1(\addroundkey_data_o[12] ),
    .A2(_04378_),
    .B1(_05607_),
    .C1(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__a21oi_2 _15088_ (.A1(\addroundkey_data_o[108] ),
    .A2(_03057_),
    .B1(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__nor2_8 _15089_ (.A(_03357_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__xnor2_2 _15090_ (.A(_03354_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__xnor2_4 _15091_ (.A(_03345_),
    .B(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__mux2_1 _15092_ (.A0(\mix1.data_reg[68] ),
    .A1(_03363_),
    .S(_03171_),
    .X(_03364_));
 sky130_fd_sc_hd__clkbuf_1 _15093_ (.A(_03364_),
    .X(_01605_));
 sky130_fd_sc_hd__a22o_1 _15094_ (.A1(\sub1.data_o[68] ),
    .A2(_03072_),
    .B1(_03068_),
    .B2(\sub1.data_o[36] ),
    .X(_03365_));
 sky130_fd_sc_hd__a211o_1 _15095_ (.A1(\sub1.data_o[4] ),
    .A2(_04379_),
    .B1(_03059_),
    .C1(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__a21oi_2 _15096_ (.A1(\sub1.data_o[100] ),
    .A2(_03057_),
    .B1(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__a22o_1 _15097_ (.A1(\addroundkey_data_o[68] ),
    .A2(_03072_),
    .B1(_03068_),
    .B2(\addroundkey_data_o[36] ),
    .X(_03368_));
 sky130_fd_sc_hd__a211o_1 _15098_ (.A1(\addroundkey_data_o[4] ),
    .A2(_04379_),
    .B1(_05607_),
    .C1(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__a21oi_4 _15099_ (.A1(\addroundkey_data_o[100] ),
    .A2(_03143_),
    .B1(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__nor2_8 _15100_ (.A(_03367_),
    .B(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__xnor2_4 _15101_ (.A(_03336_),
    .B(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__xor2_2 _15102_ (.A(_03257_),
    .B(_03273_),
    .X(_03373_));
 sky130_fd_sc_hd__xnor2_4 _15103_ (.A(_03246_),
    .B(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__xnor2_1 _15104_ (.A(_03307_),
    .B(_03352_),
    .Y(_03375_));
 sky130_fd_sc_hd__xnor2_2 _15105_ (.A(_03374_),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__o21ai_1 _15106_ (.A1(_03198_),
    .A2(_03376_),
    .B1(_06630_),
    .Y(_03377_));
 sky130_fd_sc_hd__a21oi_2 _15107_ (.A1(_03198_),
    .A2(_03376_),
    .B1(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__xnor2_4 _15108_ (.A(_03099_),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__xnor2_4 _15109_ (.A(_03115_),
    .B(_03138_),
    .Y(_03380_));
 sky130_fd_sc_hd__xor2_2 _15110_ (.A(_03379_),
    .B(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__xnor2_4 _15111_ (.A(_03372_),
    .B(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hd__mux2_1 _15112_ (.A0(net750),
    .A1(_03382_),
    .S(_03171_),
    .X(_03383_));
 sky130_fd_sc_hd__clkbuf_1 _15113_ (.A(_03383_),
    .X(_01606_));
 sky130_fd_sc_hd__xnor2_2 _15114_ (.A(_03246_),
    .B(_03297_),
    .Y(_03384_));
 sky130_fd_sc_hd__xnor2_4 _15115_ (.A(_03321_),
    .B(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__xnor2_4 _15116_ (.A(_03343_),
    .B(_03371_),
    .Y(_03386_));
 sky130_fd_sc_hd__xnor2_1 _15117_ (.A(_03354_),
    .B(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__a21oi_1 _15118_ (.A1(_03385_),
    .A2(_03387_),
    .B1(_05198_),
    .Y(_03388_));
 sky130_fd_sc_hd__o21a_2 _15119_ (.A1(_03385_),
    .A2(_03387_),
    .B1(_03388_),
    .X(_03389_));
 sky130_fd_sc_hd__xnor2_4 _15120_ (.A(_03179_),
    .B(_03195_),
    .Y(_03390_));
 sky130_fd_sc_hd__xnor2_4 _15121_ (.A(_03389_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__xor2_4 _15122_ (.A(_03140_),
    .B(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__mux2_1 _15123_ (.A0(net697),
    .A1(_03392_),
    .S(_03171_),
    .X(_03393_));
 sky130_fd_sc_hd__clkbuf_1 _15124_ (.A(_03393_),
    .X(_01607_));
 sky130_fd_sc_hd__xnor2_4 _15125_ (.A(_03167_),
    .B(_03187_),
    .Y(_03394_));
 sky130_fd_sc_hd__xnor2_4 _15126_ (.A(_03115_),
    .B(_03131_),
    .Y(_03395_));
 sky130_fd_sc_hd__xnor2_4 _15127_ (.A(_03343_),
    .B(_03361_),
    .Y(_03396_));
 sky130_fd_sc_hd__xnor2_1 _15128_ (.A(_03395_),
    .B(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__o21ai_1 _15129_ (.A1(_03372_),
    .A2(_03397_),
    .B1(_06630_),
    .Y(_03398_));
 sky130_fd_sc_hd__a21oi_1 _15130_ (.A1(_03372_),
    .A2(_03397_),
    .B1(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hd__xnor2_2 _15131_ (.A(_03245_),
    .B(_03399_),
    .Y(_03400_));
 sky130_fd_sc_hd__xor2_2 _15132_ (.A(_03180_),
    .B(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__xnor2_4 _15133_ (.A(_03394_),
    .B(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__mux2_1 _15134_ (.A0(net720),
    .A1(_03402_),
    .S(_03171_),
    .X(_03403_));
 sky130_fd_sc_hd__clkbuf_1 _15135_ (.A(_03403_),
    .X(_01608_));
 sky130_fd_sc_hd__xnor2_4 _15136_ (.A(_03099_),
    .B(_03131_),
    .Y(_03404_));
 sky130_fd_sc_hd__xor2_4 _15137_ (.A(_03380_),
    .B(_03404_),
    .X(_03405_));
 sky130_fd_sc_hd__xnor2_4 _15138_ (.A(_03390_),
    .B(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__nand2_4 _15139_ (.A(_05201_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__xnor2_1 _15140_ (.A(_03090_),
    .B(_03216_),
    .Y(_03408_));
 sky130_fd_sc_hd__xnor2_2 _15141_ (.A(_03407_),
    .B(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__xnor2_4 _15142_ (.A(_03160_),
    .B(_03245_),
    .Y(_03410_));
 sky130_fd_sc_hd__xnor2_4 _15143_ (.A(_03409_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__mux2_1 _15144_ (.A0(net769),
    .A1(_03411_),
    .S(_03171_),
    .X(_03412_));
 sky130_fd_sc_hd__clkbuf_1 _15145_ (.A(_03412_),
    .X(_01609_));
 sky130_fd_sc_hd__xnor2_4 _15146_ (.A(_03152_),
    .B(_03216_),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_2 _15147_ (.A(_03207_),
    .B(_03410_),
    .Y(_03414_));
 sky130_fd_sc_hd__xnor2_4 _15148_ (.A(_03413_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__xnor2_4 _15149_ (.A(_03107_),
    .B(_03195_),
    .Y(_03416_));
 sky130_fd_sc_hd__xor2_4 _15150_ (.A(_03167_),
    .B(_03416_),
    .X(_03417_));
 sky130_fd_sc_hd__xnor2_4 _15151_ (.A(_03124_),
    .B(_03179_),
    .Y(_03418_));
 sky130_fd_sc_hd__xnor2_2 _15152_ (.A(_03245_),
    .B(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__xnor2_4 _15153_ (.A(_03417_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__xor2_2 _15154_ (.A(_03406_),
    .B(_03420_),
    .X(_03421_));
 sky130_fd_sc_hd__nand2_2 _15155_ (.A(_05201_),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__xor2_4 _15156_ (.A(_03285_),
    .B(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__xor2_4 _15157_ (.A(_03415_),
    .B(_03423_),
    .X(_03424_));
 sky130_fd_sc_hd__buf_4 _15158_ (.A(_03144_),
    .X(_03425_));
 sky130_fd_sc_hd__mux2_1 _15159_ (.A0(net770),
    .A1(_03424_),
    .S(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__clkbuf_1 _15160_ (.A(_03426_),
    .X(_01610_));
 sky130_fd_sc_hd__xor2_1 _15161_ (.A(_03089_),
    .B(_03410_),
    .X(_03427_));
 sky130_fd_sc_hd__xnor2_1 _15162_ (.A(_03152_),
    .B(_03427_),
    .Y(_03428_));
 sky130_fd_sc_hd__xnor2_1 _15163_ (.A(_03394_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__o21ai_1 _15164_ (.A1(_03420_),
    .A2(_03429_),
    .B1(_05202_),
    .Y(_03430_));
 sky130_fd_sc_hd__a21o_4 _15165_ (.A1(_03420_),
    .A2(_03429_),
    .B1(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__xor2_2 _15166_ (.A(_03225_),
    .B(_03280_),
    .X(_03432_));
 sky130_fd_sc_hd__xor2_1 _15167_ (.A(_03273_),
    .B(_03305_),
    .X(_03433_));
 sky130_fd_sc_hd__xnor2_2 _15168_ (.A(_03432_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__xnor2_4 _15169_ (.A(_03431_),
    .B(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__mux2_1 _15170_ (.A0(net727),
    .A1(_03435_),
    .S(_03425_),
    .X(_03436_));
 sky130_fd_sc_hd__clkbuf_1 _15171_ (.A(_03436_),
    .X(_01611_));
 sky130_fd_sc_hd__xor2_2 _15172_ (.A(_03090_),
    .B(_03225_),
    .X(_03437_));
 sky130_fd_sc_hd__xnor2_4 _15173_ (.A(_03394_),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__xnor2_2 _15174_ (.A(_03406_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__a21oi_1 _15175_ (.A1(_03415_),
    .A2(_03439_),
    .B1(_05198_),
    .Y(_03440_));
 sky130_fd_sc_hd__o21ai_4 _15176_ (.A1(_03415_),
    .A2(_03439_),
    .B1(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__xnor2_2 _15177_ (.A(_03257_),
    .B(_03304_),
    .Y(_03442_));
 sky130_fd_sc_hd__xor2_1 _15178_ (.A(_03410_),
    .B(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__xor2_1 _15179_ (.A(_03297_),
    .B(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__xnor2_2 _15180_ (.A(_03353_),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__xnor2_4 _15181_ (.A(_03441_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__mux2_1 _15182_ (.A0(net760),
    .A1(_03446_),
    .S(_03425_),
    .X(_03447_));
 sky130_fd_sc_hd__clkbuf_1 _15183_ (.A(_03447_),
    .X(_01612_));
 sky130_fd_sc_hd__xor2_1 _15184_ (.A(_03233_),
    .B(_03265_),
    .X(_03448_));
 sky130_fd_sc_hd__xnor2_1 _15185_ (.A(_03281_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__a21oi_1 _15186_ (.A1(_03421_),
    .A2(_03449_),
    .B1(_05198_),
    .Y(_03450_));
 sky130_fd_sc_hd__o21a_1 _15187_ (.A1(_03421_),
    .A2(_03449_),
    .B1(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__xnor2_4 _15188_ (.A(_03386_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__xnor2_4 _15189_ (.A(_03321_),
    .B(_03352_),
    .Y(_03453_));
 sky130_fd_sc_hd__xnor2_2 _15190_ (.A(_03410_),
    .B(_03453_),
    .Y(_03454_));
 sky130_fd_sc_hd__xnor2_4 _15191_ (.A(_03336_),
    .B(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__xor2_4 _15192_ (.A(_03452_),
    .B(_03455_),
    .X(_03456_));
 sky130_fd_sc_hd__mux2_1 _15193_ (.A0(net777),
    .A1(_03456_),
    .S(_03425_),
    .X(_03457_));
 sky130_fd_sc_hd__clkbuf_1 _15194_ (.A(_03457_),
    .X(_01613_));
 sky130_fd_sc_hd__xor2_1 _15195_ (.A(_03264_),
    .B(_03273_),
    .X(_03458_));
 sky130_fd_sc_hd__xnor2_2 _15196_ (.A(_03394_),
    .B(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__xor2_1 _15197_ (.A(_03322_),
    .B(_03443_),
    .X(_03460_));
 sky130_fd_sc_hd__xnor2_1 _15198_ (.A(_03459_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__a21oi_1 _15199_ (.A1(_03420_),
    .A2(_03461_),
    .B1(_04617_),
    .Y(_03462_));
 sky130_fd_sc_hd__o21a_1 _15200_ (.A1(_03420_),
    .A2(_03461_),
    .B1(_03462_),
    .X(_03463_));
 sky130_fd_sc_hd__xnor2_4 _15201_ (.A(_03395_),
    .B(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__xnor2_2 _15202_ (.A(_03361_),
    .B(_03371_),
    .Y(_03465_));
 sky130_fd_sc_hd__xnor2_4 _15203_ (.A(_03138_),
    .B(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__xor2_4 _15204_ (.A(_03464_),
    .B(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__mux2_1 _15205_ (.A0(net780),
    .A1(_03467_),
    .S(_03425_),
    .X(_03468_));
 sky130_fd_sc_hd__clkbuf_1 _15206_ (.A(_03468_),
    .X(_01614_));
 sky130_fd_sc_hd__xor2_4 _15207_ (.A(_03107_),
    .B(_03404_),
    .X(_03469_));
 sky130_fd_sc_hd__xnor2_2 _15208_ (.A(_03297_),
    .B(_03314_),
    .Y(_03470_));
 sky130_fd_sc_hd__xor2_2 _15209_ (.A(_03361_),
    .B(_03394_),
    .X(_03471_));
 sky130_fd_sc_hd__xnor2_4 _15210_ (.A(_03470_),
    .B(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__nand2_1 _15211_ (.A(_03455_),
    .B(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__or2_1 _15212_ (.A(_03455_),
    .B(_03472_),
    .X(_03474_));
 sky130_fd_sc_hd__a21o_2 _15213_ (.A1(_03473_),
    .A2(_03474_),
    .B1(_05198_),
    .X(_03475_));
 sky130_fd_sc_hd__xor2_2 _15214_ (.A(_03418_),
    .B(_03475_),
    .X(_03476_));
 sky130_fd_sc_hd__xnor2_4 _15215_ (.A(_03469_),
    .B(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__mux2_1 _15216_ (.A0(net737),
    .A1(_03477_),
    .S(_03425_),
    .X(_03478_));
 sky130_fd_sc_hd__clkbuf_1 _15217_ (.A(_03478_),
    .X(_01615_));
 sky130_fd_sc_hd__xor2_4 _15218_ (.A(_03099_),
    .B(_03344_),
    .X(_03479_));
 sky130_fd_sc_hd__or2_1 _15219_ (.A(_03466_),
    .B(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__nand2_1 _15220_ (.A(_03466_),
    .B(_03479_),
    .Y(_03481_));
 sky130_fd_sc_hd__a21o_2 _15221_ (.A1(_03480_),
    .A2(_03481_),
    .B1(_05198_),
    .X(_03482_));
 sky130_fd_sc_hd__xor2_1 _15222_ (.A(_03188_),
    .B(_03417_),
    .X(_03483_));
 sky130_fd_sc_hd__xnor2_2 _15223_ (.A(_03482_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__mux2_1 _15224_ (.A0(net731),
    .A1(_03484_),
    .S(_03425_),
    .X(_03485_));
 sky130_fd_sc_hd__clkbuf_1 _15225_ (.A(_03485_),
    .X(_01616_));
 sky130_fd_sc_hd__xnor2_1 _15226_ (.A(_03153_),
    .B(_03246_),
    .Y(_03486_));
 sky130_fd_sc_hd__xnor2_2 _15227_ (.A(_03217_),
    .B(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__mux2_1 _15228_ (.A0(net778),
    .A1(_03487_),
    .S(_03425_),
    .X(_03488_));
 sky130_fd_sc_hd__clkbuf_1 _15229_ (.A(_03488_),
    .X(_01617_));
 sky130_fd_sc_hd__xor2_1 _15230_ (.A(_03281_),
    .B(_03288_),
    .X(_03489_));
 sky130_fd_sc_hd__xnor2_1 _15231_ (.A(_03200_),
    .B(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__xnor2_2 _15232_ (.A(_03225_),
    .B(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__mux2_1 _15233_ (.A0(net755),
    .A1(_03491_),
    .S(_03425_),
    .X(_03492_));
 sky130_fd_sc_hd__clkbuf_1 _15234_ (.A(_03492_),
    .X(_01618_));
 sky130_fd_sc_hd__xor2_2 _15235_ (.A(_03266_),
    .B(_03326_),
    .X(_03493_));
 sky130_fd_sc_hd__mux2_1 _15236_ (.A0(net748),
    .A1(_03493_),
    .S(_03425_),
    .X(_03494_));
 sky130_fd_sc_hd__clkbuf_1 _15237_ (.A(_03494_),
    .X(_01619_));
 sky130_fd_sc_hd__xor2_2 _15238_ (.A(_03314_),
    .B(_03453_),
    .X(_03495_));
 sky130_fd_sc_hd__xnor2_2 _15239_ (.A(_03290_),
    .B(_03374_),
    .Y(_03496_));
 sky130_fd_sc_hd__xnor2_4 _15240_ (.A(_03495_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__clkbuf_4 _15241_ (.A(_03144_),
    .X(_03498_));
 sky130_fd_sc_hd__mux2_1 _15242_ (.A0(net786),
    .A1(_03497_),
    .S(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__clkbuf_1 _15243_ (.A(_03499_),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_1 _15244_ (.A(_03329_),
    .B(_03361_),
    .Y(_03500_));
 sky130_fd_sc_hd__xnor2_2 _15245_ (.A(_03372_),
    .B(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__xnor2_4 _15246_ (.A(_03385_),
    .B(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__mux2_1 _15247_ (.A0(net783),
    .A1(_03502_),
    .S(_03498_),
    .X(_03503_));
 sky130_fd_sc_hd__clkbuf_1 _15248_ (.A(_03503_),
    .X(_01621_));
 sky130_fd_sc_hd__xor2_4 _15249_ (.A(_03139_),
    .B(_03379_),
    .X(_03504_));
 sky130_fd_sc_hd__xnor2_4 _15250_ (.A(_03396_),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__mux2_1 _15251_ (.A0(net775),
    .A1(_03505_),
    .S(_03498_),
    .X(_03506_));
 sky130_fd_sc_hd__clkbuf_1 _15252_ (.A(_03506_),
    .X(_01622_));
 sky130_fd_sc_hd__xnor2_4 _15253_ (.A(_03117_),
    .B(_03391_),
    .Y(_03507_));
 sky130_fd_sc_hd__mux2_1 _15254_ (.A0(net792),
    .A1(_03507_),
    .S(_03498_),
    .X(_03508_));
 sky130_fd_sc_hd__clkbuf_1 _15255_ (.A(_03508_),
    .X(_01623_));
 sky130_fd_sc_hd__xor2_2 _15256_ (.A(_03168_),
    .B(_03400_),
    .X(_03509_));
 sky130_fd_sc_hd__xnor2_4 _15257_ (.A(_03196_),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__mux2_1 _15258_ (.A0(net747),
    .A1(_03510_),
    .S(_03498_),
    .X(_03511_));
 sky130_fd_sc_hd__clkbuf_1 _15259_ (.A(_03511_),
    .X(_01624_));
 sky130_fd_sc_hd__xnor2_1 _15260_ (.A(_03394_),
    .B(_03413_),
    .Y(_03512_));
 sky130_fd_sc_hd__xnor2_2 _15261_ (.A(_03076_),
    .B(_03512_),
    .Y(_03513_));
 sky130_fd_sc_hd__xnor2_4 _15262_ (.A(_03407_),
    .B(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__mux2_1 _15263_ (.A0(net761),
    .A1(_03514_),
    .S(_03498_),
    .X(_03515_));
 sky130_fd_sc_hd__clkbuf_1 _15264_ (.A(_03515_),
    .X(_01625_));
 sky130_fd_sc_hd__xnor2_4 _15265_ (.A(_03423_),
    .B(_03438_),
    .Y(_03516_));
 sky130_fd_sc_hd__mux2_1 _15266_ (.A0(net785),
    .A1(_03516_),
    .S(_03498_),
    .X(_03517_));
 sky130_fd_sc_hd__clkbuf_1 _15267_ (.A(_03517_),
    .X(_01626_));
 sky130_fd_sc_hd__xnor2_1 _15268_ (.A(_03207_),
    .B(_03273_),
    .Y(_03518_));
 sky130_fd_sc_hd__xnor2_1 _15269_ (.A(_03232_),
    .B(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__xnor2_2 _15270_ (.A(_03442_),
    .B(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hd__xnor2_4 _15271_ (.A(_03431_),
    .B(_03520_),
    .Y(_03521_));
 sky130_fd_sc_hd__mux2_1 _15272_ (.A0(net752),
    .A1(_03521_),
    .S(_03498_),
    .X(_03522_));
 sky130_fd_sc_hd__clkbuf_1 _15273_ (.A(_03522_),
    .X(_01627_));
 sky130_fd_sc_hd__xor2_1 _15274_ (.A(_03297_),
    .B(_03453_),
    .X(_03523_));
 sky130_fd_sc_hd__xnor2_2 _15275_ (.A(_03459_),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__xnor2_4 _15276_ (.A(_03441_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__mux2_1 _15277_ (.A0(net736),
    .A1(_03525_),
    .S(_03498_),
    .X(_03526_));
 sky130_fd_sc_hd__clkbuf_1 _15278_ (.A(_03526_),
    .X(_01628_));
 sky130_fd_sc_hd__xnor2_4 _15279_ (.A(_03452_),
    .B(_03472_),
    .Y(_03527_));
 sky130_fd_sc_hd__mux2_1 _15280_ (.A0(net782),
    .A1(_03527_),
    .S(_03498_),
    .X(_03528_));
 sky130_fd_sc_hd__clkbuf_1 _15281_ (.A(_03528_),
    .X(_01629_));
 sky130_fd_sc_hd__xnor2_4 _15282_ (.A(_03464_),
    .B(_03479_),
    .Y(_03529_));
 sky130_fd_sc_hd__mux2_1 _15283_ (.A0(net773),
    .A1(_03529_),
    .S(_03144_),
    .X(_03530_));
 sky130_fd_sc_hd__clkbuf_1 _15284_ (.A(_03530_),
    .X(_01630_));
 sky130_fd_sc_hd__xnor2_1 _15285_ (.A(_03124_),
    .B(_03416_),
    .Y(_03531_));
 sky130_fd_sc_hd__xnor2_1 _15286_ (.A(_03380_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__xnor2_2 _15287_ (.A(_03475_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__mux2_1 _15288_ (.A0(net716),
    .A1(_03533_),
    .S(_03144_),
    .X(_03534_));
 sky130_fd_sc_hd__clkbuf_1 _15289_ (.A(_03534_),
    .X(_01631_));
 sky130_fd_sc_hd__xnor2_1 _15290_ (.A(_03187_),
    .B(_03418_),
    .Y(_03535_));
 sky130_fd_sc_hd__xnor2_1 _15291_ (.A(_03410_),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__xnor2_2 _15292_ (.A(_03482_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__mux2_1 _15293_ (.A0(net725),
    .A1(_03537_),
    .S(_03144_),
    .X(_03538_));
 sky130_fd_sc_hd__clkbuf_1 _15294_ (.A(_03538_),
    .X(_01632_));
 sky130_fd_sc_hd__clkbuf_4 _15295_ (.A(_03145_),
    .X(_03539_));
 sky130_fd_sc_hd__mux2_1 _15296_ (.A0(net694),
    .A1(_03170_),
    .S(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__clkbuf_1 _15297_ (.A(_03540_),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _15298_ (.A0(net772),
    .A1(_03236_),
    .S(_03539_),
    .X(_03541_));
 sky130_fd_sc_hd__clkbuf_1 _15299_ (.A(_03541_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _15300_ (.A0(net693),
    .A1(_03283_),
    .S(_03539_),
    .X(_03542_));
 sky130_fd_sc_hd__clkbuf_1 _15301_ (.A(_03542_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _15302_ (.A0(net735),
    .A1(_03324_),
    .S(_03539_),
    .X(_03543_));
 sky130_fd_sc_hd__clkbuf_1 _15303_ (.A(_03543_),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _15304_ (.A0(net700),
    .A1(_03363_),
    .S(_03539_),
    .X(_03544_));
 sky130_fd_sc_hd__clkbuf_1 _15305_ (.A(_03544_),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _15306_ (.A0(net789),
    .A1(_03382_),
    .S(_03539_),
    .X(_03545_));
 sky130_fd_sc_hd__clkbuf_1 _15307_ (.A(_03545_),
    .X(_01638_));
 sky130_fd_sc_hd__mux2_1 _15308_ (.A0(net762),
    .A1(_03392_),
    .S(_03539_),
    .X(_03546_));
 sky130_fd_sc_hd__clkbuf_1 _15309_ (.A(_03546_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _15310_ (.A0(net791),
    .A1(_03402_),
    .S(_03539_),
    .X(_03547_));
 sky130_fd_sc_hd__clkbuf_1 _15311_ (.A(_03547_),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _15312_ (.A0(net726),
    .A1(_03411_),
    .S(_03539_),
    .X(_03548_));
 sky130_fd_sc_hd__clkbuf_1 _15313_ (.A(_03548_),
    .X(_01641_));
 sky130_fd_sc_hd__buf_4 _15314_ (.A(_03145_),
    .X(_03549_));
 sky130_fd_sc_hd__mux2_1 _15315_ (.A0(net754),
    .A1(_03424_),
    .S(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__clkbuf_1 _15316_ (.A(_03550_),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _15317_ (.A0(net732),
    .A1(_03435_),
    .S(_03549_),
    .X(_03551_));
 sky130_fd_sc_hd__clkbuf_1 _15318_ (.A(_03551_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _15319_ (.A0(net723),
    .A1(_03446_),
    .S(_03549_),
    .X(_03552_));
 sky130_fd_sc_hd__clkbuf_1 _15320_ (.A(_03552_),
    .X(_01644_));
 sky130_fd_sc_hd__mux2_1 _15321_ (.A0(net767),
    .A1(_03456_),
    .S(_03549_),
    .X(_03553_));
 sky130_fd_sc_hd__clkbuf_1 _15322_ (.A(_03553_),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _15323_ (.A0(net718),
    .A1(_03467_),
    .S(_03549_),
    .X(_03554_));
 sky130_fd_sc_hd__clkbuf_1 _15324_ (.A(_03554_),
    .X(_01646_));
 sky130_fd_sc_hd__mux2_1 _15325_ (.A0(net730),
    .A1(_03477_),
    .S(_03549_),
    .X(_03555_));
 sky130_fd_sc_hd__clkbuf_1 _15326_ (.A(_03555_),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _15327_ (.A0(net768),
    .A1(_03484_),
    .S(_03549_),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_1 _15328_ (.A(_03556_),
    .X(_01648_));
 sky130_fd_sc_hd__mux2_1 _15329_ (.A0(net741),
    .A1(_03487_),
    .S(_03549_),
    .X(_03557_));
 sky130_fd_sc_hd__clkbuf_1 _15330_ (.A(_03557_),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _15331_ (.A0(\mix1.data_reg[49] ),
    .A1(_03491_),
    .S(_03549_),
    .X(_03558_));
 sky130_fd_sc_hd__clkbuf_1 _15332_ (.A(_03558_),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _15333_ (.A0(\mix1.data_reg[50] ),
    .A1(_03493_),
    .S(_03549_),
    .X(_03559_));
 sky130_fd_sc_hd__clkbuf_1 _15334_ (.A(_03559_),
    .X(_01651_));
 sky130_fd_sc_hd__clkbuf_4 _15335_ (.A(_03145_),
    .X(_03560_));
 sky130_fd_sc_hd__mux2_1 _15336_ (.A0(net763),
    .A1(_03497_),
    .S(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__clkbuf_1 _15337_ (.A(_03561_),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _15338_ (.A0(net764),
    .A1(_03502_),
    .S(_03560_),
    .X(_03562_));
 sky130_fd_sc_hd__clkbuf_1 _15339_ (.A(_03562_),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _15340_ (.A0(net740),
    .A1(_03505_),
    .S(_03560_),
    .X(_03563_));
 sky130_fd_sc_hd__clkbuf_1 _15341_ (.A(_03563_),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _15342_ (.A0(net710),
    .A1(_03507_),
    .S(_03560_),
    .X(_03564_));
 sky130_fd_sc_hd__clkbuf_1 _15343_ (.A(_03564_),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _15344_ (.A0(net734),
    .A1(_03510_),
    .S(_03560_),
    .X(_03565_));
 sky130_fd_sc_hd__clkbuf_1 _15345_ (.A(_03565_),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _15346_ (.A0(net756),
    .A1(_03514_),
    .S(_03560_),
    .X(_03566_));
 sky130_fd_sc_hd__clkbuf_1 _15347_ (.A(_03566_),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _15348_ (.A0(net715),
    .A1(_03516_),
    .S(_03560_),
    .X(_03567_));
 sky130_fd_sc_hd__clkbuf_1 _15349_ (.A(_03567_),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _15350_ (.A0(net798),
    .A1(_03521_),
    .S(_03560_),
    .X(_03568_));
 sky130_fd_sc_hd__clkbuf_1 _15351_ (.A(_03568_),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _15352_ (.A0(net743),
    .A1(_03525_),
    .S(_03560_),
    .X(_03569_));
 sky130_fd_sc_hd__clkbuf_1 _15353_ (.A(_03569_),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _15354_ (.A0(net742),
    .A1(_03527_),
    .S(_03560_),
    .X(_03570_));
 sky130_fd_sc_hd__clkbuf_1 _15355_ (.A(_03570_),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _15356_ (.A0(net724),
    .A1(_03529_),
    .S(_03145_),
    .X(_03571_));
 sky130_fd_sc_hd__clkbuf_1 _15357_ (.A(_03571_),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _15358_ (.A0(\mix1.data_reg[62] ),
    .A1(_03533_),
    .S(_03145_),
    .X(_03572_));
 sky130_fd_sc_hd__clkbuf_1 _15359_ (.A(_03572_),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _15360_ (.A0(\mix1.data_reg[63] ),
    .A1(_03537_),
    .S(_03145_),
    .X(_03573_));
 sky130_fd_sc_hd__clkbuf_1 _15361_ (.A(_03573_),
    .X(_01664_));
 sky130_fd_sc_hd__buf_4 _15362_ (.A(_05202_),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_1 _15363_ (.A0(\sub1.data_o[32] ),
    .A1(\sub1.data_o[96] ),
    .S(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__buf_4 _15364_ (.A(_04368_),
    .X(_03576_));
 sky130_fd_sc_hd__mux2_1 _15365_ (.A0(\sub1.data_o[0] ),
    .A1(_03575_),
    .S(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__clkbuf_1 _15366_ (.A(_03577_),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _15367_ (.A0(\sub1.data_o[33] ),
    .A1(\sub1.data_o[97] ),
    .S(_03574_),
    .X(_03578_));
 sky130_fd_sc_hd__mux2_1 _15368_ (.A0(\sub1.data_o[1] ),
    .A1(_03578_),
    .S(_03576_),
    .X(_03579_));
 sky130_fd_sc_hd__clkbuf_1 _15369_ (.A(_03579_),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _15370_ (.A0(\sub1.data_o[34] ),
    .A1(\sub1.data_o[98] ),
    .S(_03574_),
    .X(_03580_));
 sky130_fd_sc_hd__clkbuf_8 _15371_ (.A(_04368_),
    .X(_03581_));
 sky130_fd_sc_hd__mux2_1 _15372_ (.A0(\sub1.data_o[2] ),
    .A1(_03580_),
    .S(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__clkbuf_1 _15373_ (.A(_03582_),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_1 _15374_ (.A0(\sub1.data_o[35] ),
    .A1(\sub1.data_o[99] ),
    .S(_03574_),
    .X(_03583_));
 sky130_fd_sc_hd__mux2_1 _15375_ (.A0(\sub1.data_o[3] ),
    .A1(_03583_),
    .S(_03581_),
    .X(_03584_));
 sky130_fd_sc_hd__clkbuf_1 _15376_ (.A(_03584_),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _15377_ (.A0(\sub1.data_o[36] ),
    .A1(\sub1.data_o[100] ),
    .S(_05202_),
    .X(_03585_));
 sky130_fd_sc_hd__mux2_1 _15378_ (.A0(\sub1.data_o[4] ),
    .A1(_03585_),
    .S(_03581_),
    .X(_03586_));
 sky130_fd_sc_hd__clkbuf_1 _15379_ (.A(_03586_),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _15380_ (.A0(\sub1.data_o[37] ),
    .A1(\sub1.data_o[101] ),
    .S(_05202_),
    .X(_03587_));
 sky130_fd_sc_hd__mux2_1 _15381_ (.A0(\sub1.data_o[5] ),
    .A1(_03587_),
    .S(_03581_),
    .X(_03588_));
 sky130_fd_sc_hd__clkbuf_1 _15382_ (.A(_03588_),
    .X(_01670_));
 sky130_fd_sc_hd__mux2_1 _15383_ (.A0(\sub1.data_o[38] ),
    .A1(\sub1.data_o[102] ),
    .S(_05202_),
    .X(_03589_));
 sky130_fd_sc_hd__mux2_1 _15384_ (.A0(\sub1.data_o[6] ),
    .A1(_03589_),
    .S(_03581_),
    .X(_03590_));
 sky130_fd_sc_hd__clkbuf_1 _15385_ (.A(_03590_),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _15386_ (.A0(\sub1.data_o[39] ),
    .A1(\sub1.data_o[103] ),
    .S(_05202_),
    .X(_03591_));
 sky130_fd_sc_hd__mux2_1 _15387_ (.A0(\sub1.data_o[7] ),
    .A1(_03591_),
    .S(_03581_),
    .X(_03592_));
 sky130_fd_sc_hd__clkbuf_1 _15388_ (.A(_03592_),
    .X(_01672_));
 sky130_fd_sc_hd__clkbuf_4 _15389_ (.A(_04689_),
    .X(_03593_));
 sky130_fd_sc_hd__buf_4 _15390_ (.A(_04369_),
    .X(_03594_));
 sky130_fd_sc_hd__nor2_2 _15391_ (.A(_03581_),
    .B(_04689_),
    .Y(_03595_));
 sky130_fd_sc_hd__a22o_1 _15392_ (.A1(\sub1.data_o[72] ),
    .A2(_03594_),
    .B1(_03595_),
    .B2(\sub1.data_o[8] ),
    .X(_03596_));
 sky130_fd_sc_hd__a31o_1 _15393_ (.A1(_03019_),
    .A2(_03593_),
    .A3(_05548_),
    .B1(_03596_),
    .X(_01673_));
 sky130_fd_sc_hd__a22o_1 _15394_ (.A1(\sub1.data_o[73] ),
    .A2(_03594_),
    .B1(_03595_),
    .B2(\sub1.data_o[9] ),
    .X(_03597_));
 sky130_fd_sc_hd__a31o_1 _15395_ (.A1(_03019_),
    .A2(_03593_),
    .A3(_05554_),
    .B1(_03597_),
    .X(_01674_));
 sky130_fd_sc_hd__a22o_1 _15396_ (.A1(\sub1.data_o[74] ),
    .A2(_03594_),
    .B1(_03595_),
    .B2(\sub1.data_o[10] ),
    .X(_03598_));
 sky130_fd_sc_hd__a31o_1 _15397_ (.A1(_03019_),
    .A2(_03593_),
    .A3(_05560_),
    .B1(_03598_),
    .X(_01675_));
 sky130_fd_sc_hd__a22o_1 _15398_ (.A1(\sub1.data_o[75] ),
    .A2(_03594_),
    .B1(_03595_),
    .B2(\sub1.data_o[11] ),
    .X(_03599_));
 sky130_fd_sc_hd__a31o_1 _15399_ (.A1(_03019_),
    .A2(_03593_),
    .A3(_05196_),
    .B1(_03599_),
    .X(_01676_));
 sky130_fd_sc_hd__clkbuf_4 _15400_ (.A(_04369_),
    .X(_03600_));
 sky130_fd_sc_hd__a22o_1 _15401_ (.A1(\sub1.data_o[76] ),
    .A2(_03600_),
    .B1(_03595_),
    .B2(\sub1.data_o[12] ),
    .X(_03601_));
 sky130_fd_sc_hd__a31o_1 _15402_ (.A1(_03019_),
    .A2(_03593_),
    .A3(_05219_),
    .B1(_03601_),
    .X(_01677_));
 sky130_fd_sc_hd__a22o_1 _15403_ (.A1(\sub1.data_o[77] ),
    .A2(_03600_),
    .B1(_03595_),
    .B2(\sub1.data_o[13] ),
    .X(_03602_));
 sky130_fd_sc_hd__a31o_1 _15404_ (.A1(_03019_),
    .A2(_03593_),
    .A3(_05228_),
    .B1(_03602_),
    .X(_01678_));
 sky130_fd_sc_hd__clkbuf_4 _15405_ (.A(_05103_),
    .X(_03603_));
 sky130_fd_sc_hd__a22o_1 _15406_ (.A1(\sub1.data_o[78] ),
    .A2(_03600_),
    .B1(_03595_),
    .B2(\sub1.data_o[14] ),
    .X(_03604_));
 sky130_fd_sc_hd__a31o_1 _15407_ (.A1(_03603_),
    .A2(_03593_),
    .A3(_05236_),
    .B1(_03604_),
    .X(_01679_));
 sky130_fd_sc_hd__a22o_1 _15408_ (.A1(\sub1.data_o[79] ),
    .A2(_03600_),
    .B1(_03595_),
    .B2(\sub1.data_o[15] ),
    .X(_03605_));
 sky130_fd_sc_hd__a31o_1 _15409_ (.A1(_03603_),
    .A2(_03593_),
    .A3(_05245_),
    .B1(_03605_),
    .X(_01680_));
 sky130_fd_sc_hd__nor2_2 _15410_ (.A(_04369_),
    .B(_04949_),
    .Y(_03606_));
 sky130_fd_sc_hd__mux2_1 _15411_ (.A0(\sub1.data_o[112] ),
    .A1(\sub1.data_o[48] ),
    .S(_05598_),
    .X(_03607_));
 sky130_fd_sc_hd__a22o_1 _15412_ (.A1(\sub1.data_o[16] ),
    .A2(_03606_),
    .B1(_03607_),
    .B2(\sub1.next_ready_o ),
    .X(_03608_));
 sky130_fd_sc_hd__a31o_1 _15413_ (.A1(_03603_),
    .A2(_04949_),
    .A3(_05548_),
    .B1(_03608_),
    .X(_01681_));
 sky130_fd_sc_hd__clkbuf_4 _15414_ (.A(_05202_),
    .X(_03609_));
 sky130_fd_sc_hd__mux2_1 _15415_ (.A0(\sub1.data_o[113] ),
    .A1(\sub1.data_o[49] ),
    .S(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__clkbuf_4 _15416_ (.A(_03581_),
    .X(_03611_));
 sky130_fd_sc_hd__a22o_1 _15417_ (.A1(\sub1.data_o[17] ),
    .A2(_03606_),
    .B1(_03610_),
    .B2(_03611_),
    .X(_03612_));
 sky130_fd_sc_hd__a31o_1 _15418_ (.A1(_03603_),
    .A2(_04949_),
    .A3(_05554_),
    .B1(_03612_),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _15419_ (.A0(\sub1.data_o[114] ),
    .A1(\sub1.data_o[50] ),
    .S(_03609_),
    .X(_03613_));
 sky130_fd_sc_hd__a22o_1 _15420_ (.A1(\sub1.data_o[18] ),
    .A2(_03606_),
    .B1(_03613_),
    .B2(_03611_),
    .X(_03614_));
 sky130_fd_sc_hd__a31o_1 _15421_ (.A1(_03603_),
    .A2(_04949_),
    .A3(_05560_),
    .B1(_03614_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _15422_ (.A0(\sub1.data_o[115] ),
    .A1(\sub1.data_o[51] ),
    .S(_03609_),
    .X(_03615_));
 sky130_fd_sc_hd__a22o_1 _15423_ (.A1(\sub1.data_o[19] ),
    .A2(_03606_),
    .B1(_03615_),
    .B2(_03611_),
    .X(_03616_));
 sky130_fd_sc_hd__a31o_1 _15424_ (.A1(_03603_),
    .A2(_04949_),
    .A3(_05196_),
    .B1(_03616_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _15425_ (.A0(\sub1.data_o[116] ),
    .A1(\sub1.data_o[52] ),
    .S(_03609_),
    .X(_03617_));
 sky130_fd_sc_hd__a22o_1 _15426_ (.A1(\sub1.data_o[20] ),
    .A2(_03606_),
    .B1(_03617_),
    .B2(_03611_),
    .X(_03618_));
 sky130_fd_sc_hd__a31o_1 _15427_ (.A1(_03603_),
    .A2(_04949_),
    .A3(_05219_),
    .B1(_03618_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _15428_ (.A0(\sub1.data_o[117] ),
    .A1(\sub1.data_o[53] ),
    .S(_03609_),
    .X(_03619_));
 sky130_fd_sc_hd__a22o_1 _15429_ (.A1(\sub1.data_o[21] ),
    .A2(_03606_),
    .B1(_03619_),
    .B2(_03611_),
    .X(_03620_));
 sky130_fd_sc_hd__a31o_1 _15430_ (.A1(_03603_),
    .A2(_04949_),
    .A3(_05228_),
    .B1(_03620_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _15431_ (.A0(\sub1.data_o[118] ),
    .A1(\sub1.data_o[54] ),
    .S(_03609_),
    .X(_03621_));
 sky130_fd_sc_hd__a22o_1 _15432_ (.A1(\sub1.data_o[22] ),
    .A2(_03606_),
    .B1(_03621_),
    .B2(_03611_),
    .X(_03622_));
 sky130_fd_sc_hd__a31o_1 _15433_ (.A1(_03603_),
    .A2(_04949_),
    .A3(_05236_),
    .B1(_03622_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _15434_ (.A0(\sub1.data_o[119] ),
    .A1(\sub1.data_o[55] ),
    .S(_03609_),
    .X(_03623_));
 sky130_fd_sc_hd__a22o_1 _15435_ (.A1(\sub1.data_o[23] ),
    .A2(_03606_),
    .B1(_03623_),
    .B2(_03611_),
    .X(_03624_));
 sky130_fd_sc_hd__a31o_1 _15436_ (.A1(_03603_),
    .A2(_04949_),
    .A3(_05245_),
    .B1(_03624_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _15437_ (.A0(\sub1.data_o[24] ),
    .A1(_05547_),
    .S(_04879_),
    .X(_03625_));
 sky130_fd_sc_hd__clkbuf_1 _15438_ (.A(_03625_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _15439_ (.A0(\sub1.data_o[25] ),
    .A1(_05553_),
    .S(_04879_),
    .X(_03626_));
 sky130_fd_sc_hd__clkbuf_1 _15440_ (.A(_03626_),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _15441_ (.A0(\sub1.data_o[26] ),
    .A1(_05559_),
    .S(_04879_),
    .X(_03627_));
 sky130_fd_sc_hd__clkbuf_1 _15442_ (.A(_03627_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _15443_ (.A0(\sub1.data_o[27] ),
    .A1(_05195_),
    .S(_04879_),
    .X(_03628_));
 sky130_fd_sc_hd__clkbuf_1 _15444_ (.A(_03628_),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _15445_ (.A0(\sub1.data_o[28] ),
    .A1(_05218_),
    .S(_04879_),
    .X(_03629_));
 sky130_fd_sc_hd__clkbuf_1 _15446_ (.A(_03629_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _15447_ (.A0(\sub1.data_o[29] ),
    .A1(_05227_),
    .S(_04879_),
    .X(_03630_));
 sky130_fd_sc_hd__clkbuf_1 _15448_ (.A(_03630_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _15449_ (.A0(\sub1.data_o[30] ),
    .A1(_05235_),
    .S(_04879_),
    .X(_03631_));
 sky130_fd_sc_hd__clkbuf_1 _15450_ (.A(_03631_),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_1 _15451_ (.A0(\sub1.data_o[31] ),
    .A1(_05244_),
    .S(_04879_),
    .X(_03632_));
 sky130_fd_sc_hd__clkbuf_1 _15452_ (.A(_03632_),
    .X(_01696_));
 sky130_fd_sc_hd__nand2_4 _15453_ (.A(_05198_),
    .B(_04368_),
    .Y(_03633_));
 sky130_fd_sc_hd__mux2_1 _15454_ (.A0(\sub1.data_o[64] ),
    .A1(_05547_),
    .S(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__or2_1 _15455_ (.A(_04368_),
    .B(_04675_),
    .X(_03635_));
 sky130_fd_sc_hd__clkbuf_4 _15456_ (.A(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__mux2_1 _15457_ (.A0(\sub1.data_o[32] ),
    .A1(_03634_),
    .S(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__clkbuf_1 _15458_ (.A(_03637_),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _15459_ (.A0(\sub1.data_o[65] ),
    .A1(_05553_),
    .S(_03633_),
    .X(_03638_));
 sky130_fd_sc_hd__mux2_1 _15460_ (.A0(\sub1.data_o[33] ),
    .A1(_03638_),
    .S(_03636_),
    .X(_03639_));
 sky130_fd_sc_hd__clkbuf_1 _15461_ (.A(_03639_),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _15462_ (.A0(\sub1.data_o[66] ),
    .A1(_05559_),
    .S(_03633_),
    .X(_03640_));
 sky130_fd_sc_hd__mux2_1 _15463_ (.A0(\sub1.data_o[34] ),
    .A1(_03640_),
    .S(_03636_),
    .X(_03641_));
 sky130_fd_sc_hd__clkbuf_1 _15464_ (.A(_03641_),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _15465_ (.A0(\sub1.data_o[67] ),
    .A1(_05195_),
    .S(_03633_),
    .X(_03642_));
 sky130_fd_sc_hd__mux2_1 _15466_ (.A0(\sub1.data_o[35] ),
    .A1(_03642_),
    .S(_03636_),
    .X(_03643_));
 sky130_fd_sc_hd__clkbuf_1 _15467_ (.A(_03643_),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _15468_ (.A0(\sub1.data_o[68] ),
    .A1(_05218_),
    .S(_03633_),
    .X(_03644_));
 sky130_fd_sc_hd__mux2_1 _15469_ (.A0(\sub1.data_o[36] ),
    .A1(_03644_),
    .S(_03636_),
    .X(_03645_));
 sky130_fd_sc_hd__clkbuf_1 _15470_ (.A(_03645_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _15471_ (.A0(\sub1.data_o[69] ),
    .A1(_05227_),
    .S(_03633_),
    .X(_03646_));
 sky130_fd_sc_hd__mux2_1 _15472_ (.A0(\sub1.data_o[37] ),
    .A1(_03646_),
    .S(_03636_),
    .X(_03647_));
 sky130_fd_sc_hd__clkbuf_1 _15473_ (.A(_03647_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _15474_ (.A0(\sub1.data_o[70] ),
    .A1(_05235_),
    .S(_03633_),
    .X(_03648_));
 sky130_fd_sc_hd__mux2_1 _15475_ (.A0(\sub1.data_o[38] ),
    .A1(_03648_),
    .S(_03636_),
    .X(_03649_));
 sky130_fd_sc_hd__clkbuf_1 _15476_ (.A(_03649_),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _15477_ (.A0(\sub1.data_o[71] ),
    .A1(_05244_),
    .S(_03633_),
    .X(_03650_));
 sky130_fd_sc_hd__mux2_1 _15478_ (.A0(\sub1.data_o[39] ),
    .A1(_03650_),
    .S(_03636_),
    .X(_03651_));
 sky130_fd_sc_hd__clkbuf_1 _15479_ (.A(_03651_),
    .X(_01704_));
 sky130_fd_sc_hd__buf_4 _15480_ (.A(_05103_),
    .X(_03652_));
 sky130_fd_sc_hd__nor2_2 _15481_ (.A(_03581_),
    .B(_04784_),
    .Y(_03653_));
 sky130_fd_sc_hd__a22o_1 _15482_ (.A1(\sub1.data_o[104] ),
    .A2(_03600_),
    .B1(_03653_),
    .B2(\sub1.data_o[40] ),
    .X(_03654_));
 sky130_fd_sc_hd__a31o_1 _15483_ (.A1(_03652_),
    .A2(_04784_),
    .A3(_05548_),
    .B1(_03654_),
    .X(_01705_));
 sky130_fd_sc_hd__a22o_1 _15484_ (.A1(\sub1.data_o[105] ),
    .A2(_03600_),
    .B1(_03653_),
    .B2(\sub1.data_o[41] ),
    .X(_03655_));
 sky130_fd_sc_hd__a31o_1 _15485_ (.A1(_03652_),
    .A2(_04784_),
    .A3(_05554_),
    .B1(_03655_),
    .X(_01706_));
 sky130_fd_sc_hd__a22o_1 _15486_ (.A1(\sub1.data_o[106] ),
    .A2(_03600_),
    .B1(_03653_),
    .B2(\sub1.data_o[42] ),
    .X(_03656_));
 sky130_fd_sc_hd__a31o_1 _15487_ (.A1(_03652_),
    .A2(_04784_),
    .A3(_05560_),
    .B1(_03656_),
    .X(_01707_));
 sky130_fd_sc_hd__a22o_1 _15488_ (.A1(\sub1.data_o[107] ),
    .A2(_03600_),
    .B1(_03653_),
    .B2(\sub1.data_o[43] ),
    .X(_03657_));
 sky130_fd_sc_hd__a31o_1 _15489_ (.A1(_03652_),
    .A2(_04784_),
    .A3(_05196_),
    .B1(_03657_),
    .X(_01708_));
 sky130_fd_sc_hd__a22o_1 _15490_ (.A1(\sub1.data_o[108] ),
    .A2(_03600_),
    .B1(_03653_),
    .B2(\sub1.data_o[44] ),
    .X(_03658_));
 sky130_fd_sc_hd__a31o_1 _15491_ (.A1(_03652_),
    .A2(_04784_),
    .A3(_05219_),
    .B1(_03658_),
    .X(_01709_));
 sky130_fd_sc_hd__a22o_1 _15492_ (.A1(\sub1.data_o[109] ),
    .A2(_03600_),
    .B1(_03653_),
    .B2(\sub1.data_o[45] ),
    .X(_03659_));
 sky130_fd_sc_hd__a31o_1 _15493_ (.A1(_03652_),
    .A2(_04784_),
    .A3(_05228_),
    .B1(_03659_),
    .X(_01710_));
 sky130_fd_sc_hd__clkbuf_4 _15494_ (.A(_04369_),
    .X(_03660_));
 sky130_fd_sc_hd__a22o_1 _15495_ (.A1(\sub1.data_o[110] ),
    .A2(_03660_),
    .B1(_03653_),
    .B2(\sub1.data_o[46] ),
    .X(_03661_));
 sky130_fd_sc_hd__a31o_1 _15496_ (.A1(_03652_),
    .A2(_04784_),
    .A3(_05236_),
    .B1(_03661_),
    .X(_01711_));
 sky130_fd_sc_hd__a22o_1 _15497_ (.A1(\sub1.data_o[111] ),
    .A2(_03660_),
    .B1(_03653_),
    .B2(\sub1.data_o[47] ),
    .X(_03662_));
 sky130_fd_sc_hd__a31o_1 _15498_ (.A1(_03652_),
    .A2(_04784_),
    .A3(_05245_),
    .B1(_03662_),
    .X(_01712_));
 sky130_fd_sc_hd__nor2_4 _15499_ (.A(_04369_),
    .B(_04777_),
    .Y(_03663_));
 sky130_fd_sc_hd__mux2_1 _15500_ (.A0(\sub1.data_o[16] ),
    .A1(\sub1.data_o[80] ),
    .S(_03609_),
    .X(_03664_));
 sky130_fd_sc_hd__a22o_1 _15501_ (.A1(\sub1.data_o[48] ),
    .A2(_03663_),
    .B1(_03664_),
    .B2(_03611_),
    .X(_03665_));
 sky130_fd_sc_hd__a31o_1 _15502_ (.A1(_03652_),
    .A2(_04777_),
    .A3(_05548_),
    .B1(_03665_),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _15503_ (.A0(\sub1.data_o[17] ),
    .A1(\sub1.data_o[81] ),
    .S(_03609_),
    .X(_03666_));
 sky130_fd_sc_hd__a22o_1 _15504_ (.A1(\sub1.data_o[49] ),
    .A2(_03663_),
    .B1(_03666_),
    .B2(_03611_),
    .X(_03667_));
 sky130_fd_sc_hd__a31o_1 _15505_ (.A1(_03652_),
    .A2(_04777_),
    .A3(_05554_),
    .B1(_03667_),
    .X(_01714_));
 sky130_fd_sc_hd__clkbuf_4 _15506_ (.A(_05103_),
    .X(_03668_));
 sky130_fd_sc_hd__mux2_1 _15507_ (.A0(\sub1.data_o[18] ),
    .A1(\sub1.data_o[82] ),
    .S(_03609_),
    .X(_03669_));
 sky130_fd_sc_hd__a22o_1 _15508_ (.A1(\sub1.data_o[50] ),
    .A2(_03663_),
    .B1(_03669_),
    .B2(_03611_),
    .X(_03670_));
 sky130_fd_sc_hd__a31o_1 _15509_ (.A1(_03668_),
    .A2(_04777_),
    .A3(_05560_),
    .B1(_03670_),
    .X(_01715_));
 sky130_fd_sc_hd__clkbuf_4 _15510_ (.A(_05202_),
    .X(_03671_));
 sky130_fd_sc_hd__mux2_1 _15511_ (.A0(\sub1.data_o[19] ),
    .A1(\sub1.data_o[83] ),
    .S(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__clkbuf_4 _15512_ (.A(_03581_),
    .X(_03673_));
 sky130_fd_sc_hd__a22o_1 _15513_ (.A1(\sub1.data_o[51] ),
    .A2(_03663_),
    .B1(_03672_),
    .B2(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__a31o_1 _15514_ (.A1(_03668_),
    .A2(_04777_),
    .A3(_05196_),
    .B1(_03674_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _15515_ (.A0(\sub1.data_o[20] ),
    .A1(\sub1.data_o[84] ),
    .S(_03671_),
    .X(_03675_));
 sky130_fd_sc_hd__a22o_1 _15516_ (.A1(\sub1.data_o[52] ),
    .A2(_03663_),
    .B1(_03675_),
    .B2(_03673_),
    .X(_03676_));
 sky130_fd_sc_hd__a31o_1 _15517_ (.A1(_03668_),
    .A2(_04777_),
    .A3(_05219_),
    .B1(_03676_),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _15518_ (.A0(\sub1.data_o[21] ),
    .A1(\sub1.data_o[85] ),
    .S(_03671_),
    .X(_03677_));
 sky130_fd_sc_hd__a22o_1 _15519_ (.A1(\sub1.data_o[53] ),
    .A2(_03663_),
    .B1(_03677_),
    .B2(_03673_),
    .X(_03678_));
 sky130_fd_sc_hd__a31o_1 _15520_ (.A1(_03668_),
    .A2(_04777_),
    .A3(_05228_),
    .B1(_03678_),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _15521_ (.A0(\sub1.data_o[22] ),
    .A1(\sub1.data_o[86] ),
    .S(_03671_),
    .X(_03679_));
 sky130_fd_sc_hd__a22o_1 _15522_ (.A1(\sub1.data_o[54] ),
    .A2(_03663_),
    .B1(_03679_),
    .B2(_03673_),
    .X(_03680_));
 sky130_fd_sc_hd__a31o_1 _15523_ (.A1(_03668_),
    .A2(_04777_),
    .A3(_05236_),
    .B1(_03680_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _15524_ (.A0(\sub1.data_o[23] ),
    .A1(\sub1.data_o[87] ),
    .S(_03671_),
    .X(_03681_));
 sky130_fd_sc_hd__a22o_1 _15525_ (.A1(\sub1.data_o[55] ),
    .A2(_03663_),
    .B1(_03681_),
    .B2(_03673_),
    .X(_03682_));
 sky130_fd_sc_hd__a31o_1 _15526_ (.A1(_03668_),
    .A2(_04777_),
    .A3(_05245_),
    .B1(_03682_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _15527_ (.A0(\sub1.data_o[56] ),
    .A1(_05547_),
    .S(_04884_),
    .X(_03683_));
 sky130_fd_sc_hd__clkbuf_1 _15528_ (.A(_03683_),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _15529_ (.A0(\sub1.data_o[57] ),
    .A1(_05553_),
    .S(_04884_),
    .X(_03684_));
 sky130_fd_sc_hd__clkbuf_1 _15530_ (.A(_03684_),
    .X(_01722_));
 sky130_fd_sc_hd__mux2_1 _15531_ (.A0(\sub1.data_o[58] ),
    .A1(_05559_),
    .S(_04884_),
    .X(_03685_));
 sky130_fd_sc_hd__clkbuf_1 _15532_ (.A(_03685_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _15533_ (.A0(\sub1.data_o[59] ),
    .A1(_05195_),
    .S(_04884_),
    .X(_03686_));
 sky130_fd_sc_hd__clkbuf_1 _15534_ (.A(_03686_),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _15535_ (.A0(\sub1.data_o[60] ),
    .A1(_05218_),
    .S(_04884_),
    .X(_03687_));
 sky130_fd_sc_hd__clkbuf_1 _15536_ (.A(_03687_),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _15537_ (.A0(\sub1.data_o[61] ),
    .A1(_05227_),
    .S(_04884_),
    .X(_03688_));
 sky130_fd_sc_hd__clkbuf_1 _15538_ (.A(_03688_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _15539_ (.A0(\sub1.data_o[62] ),
    .A1(_05235_),
    .S(_04884_),
    .X(_03689_));
 sky130_fd_sc_hd__clkbuf_1 _15540_ (.A(_03689_),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _15541_ (.A0(\sub1.data_o[63] ),
    .A1(_05244_),
    .S(_04884_),
    .X(_03690_));
 sky130_fd_sc_hd__clkbuf_1 _15542_ (.A(_03690_),
    .X(_01728_));
 sky130_fd_sc_hd__nor2_2 _15543_ (.A(_04368_),
    .B(_04935_),
    .Y(_03691_));
 sky130_fd_sc_hd__mux2_1 _15544_ (.A0(\sub1.data_o[96] ),
    .A1(\sub1.data_o[32] ),
    .S(_03671_),
    .X(_03692_));
 sky130_fd_sc_hd__a22o_1 _15545_ (.A1(\sub1.data_o[64] ),
    .A2(_03691_),
    .B1(_03692_),
    .B2(_03673_),
    .X(_03693_));
 sky130_fd_sc_hd__a31o_1 _15546_ (.A1(_03668_),
    .A2(_04935_),
    .A3(_05548_),
    .B1(_03693_),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_1 _15547_ (.A0(\sub1.data_o[97] ),
    .A1(\sub1.data_o[33] ),
    .S(_03671_),
    .X(_03694_));
 sky130_fd_sc_hd__a22o_1 _15548_ (.A1(\sub1.data_o[65] ),
    .A2(_03691_),
    .B1(_03694_),
    .B2(_03673_),
    .X(_03695_));
 sky130_fd_sc_hd__a31o_1 _15549_ (.A1(_03668_),
    .A2(_04935_),
    .A3(_05554_),
    .B1(_03695_),
    .X(_01730_));
 sky130_fd_sc_hd__mux2_1 _15550_ (.A0(\sub1.data_o[98] ),
    .A1(\sub1.data_o[34] ),
    .S(_03671_),
    .X(_03696_));
 sky130_fd_sc_hd__a22o_1 _15551_ (.A1(\sub1.data_o[66] ),
    .A2(_03691_),
    .B1(_03696_),
    .B2(_03673_),
    .X(_03697_));
 sky130_fd_sc_hd__a31o_1 _15552_ (.A1(_03668_),
    .A2(_04935_),
    .A3(_05560_),
    .B1(_03697_),
    .X(_01731_));
 sky130_fd_sc_hd__mux2_1 _15553_ (.A0(\sub1.data_o[99] ),
    .A1(\sub1.data_o[35] ),
    .S(_03671_),
    .X(_03698_));
 sky130_fd_sc_hd__a22o_1 _15554_ (.A1(\sub1.data_o[67] ),
    .A2(_03691_),
    .B1(_03698_),
    .B2(_03673_),
    .X(_03699_));
 sky130_fd_sc_hd__a31o_1 _15555_ (.A1(_03668_),
    .A2(_04935_),
    .A3(_05196_),
    .B1(_03699_),
    .X(_01732_));
 sky130_fd_sc_hd__buf_4 _15556_ (.A(_05103_),
    .X(_03700_));
 sky130_fd_sc_hd__mux2_1 _15557_ (.A0(\sub1.data_o[100] ),
    .A1(\sub1.data_o[36] ),
    .S(_03671_),
    .X(_03701_));
 sky130_fd_sc_hd__a22o_1 _15558_ (.A1(\sub1.data_o[68] ),
    .A2(_03691_),
    .B1(_03701_),
    .B2(_03673_),
    .X(_03702_));
 sky130_fd_sc_hd__a31o_1 _15559_ (.A1(_03700_),
    .A2(_04935_),
    .A3(_05219_),
    .B1(_03702_),
    .X(_01733_));
 sky130_fd_sc_hd__mux2_1 _15560_ (.A0(\sub1.data_o[101] ),
    .A1(\sub1.data_o[37] ),
    .S(_03574_),
    .X(_03703_));
 sky130_fd_sc_hd__a22o_1 _15561_ (.A1(\sub1.data_o[69] ),
    .A2(_03691_),
    .B1(_03703_),
    .B2(_03594_),
    .X(_03704_));
 sky130_fd_sc_hd__a31o_1 _15562_ (.A1(_03700_),
    .A2(_04935_),
    .A3(_05228_),
    .B1(_03704_),
    .X(_01734_));
 sky130_fd_sc_hd__mux2_1 _15563_ (.A0(\sub1.data_o[102] ),
    .A1(\sub1.data_o[38] ),
    .S(_03574_),
    .X(_03705_));
 sky130_fd_sc_hd__a22o_1 _15564_ (.A1(\sub1.data_o[70] ),
    .A2(_03691_),
    .B1(_03705_),
    .B2(_03594_),
    .X(_03706_));
 sky130_fd_sc_hd__a31o_1 _15565_ (.A1(_03700_),
    .A2(_04935_),
    .A3(_05236_),
    .B1(_03706_),
    .X(_01735_));
 sky130_fd_sc_hd__mux2_1 _15566_ (.A0(\sub1.data_o[103] ),
    .A1(\sub1.data_o[39] ),
    .S(_03574_),
    .X(_03707_));
 sky130_fd_sc_hd__a22o_1 _15567_ (.A1(\sub1.data_o[71] ),
    .A2(_03691_),
    .B1(_03707_),
    .B2(_03594_),
    .X(_03708_));
 sky130_fd_sc_hd__a31o_1 _15568_ (.A1(_03700_),
    .A2(_04935_),
    .A3(_05245_),
    .B1(_03708_),
    .X(_01736_));
 sky130_fd_sc_hd__clkbuf_4 _15569_ (.A(_04713_),
    .X(_03709_));
 sky130_fd_sc_hd__nor2_2 _15570_ (.A(_04369_),
    .B(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__a22o_1 _15571_ (.A1(\sub1.data_o[8] ),
    .A2(_03660_),
    .B1(_03710_),
    .B2(\sub1.data_o[72] ),
    .X(_03711_));
 sky130_fd_sc_hd__a31o_1 _15572_ (.A1(_03700_),
    .A2(_03709_),
    .A3(_05548_),
    .B1(_03711_),
    .X(_01737_));
 sky130_fd_sc_hd__a22o_1 _15573_ (.A1(\sub1.data_o[9] ),
    .A2(_03660_),
    .B1(_03710_),
    .B2(\sub1.data_o[73] ),
    .X(_03712_));
 sky130_fd_sc_hd__a31o_1 _15574_ (.A1(_03700_),
    .A2(_03709_),
    .A3(_05554_),
    .B1(_03712_),
    .X(_01738_));
 sky130_fd_sc_hd__a22o_1 _15575_ (.A1(\sub1.data_o[10] ),
    .A2(_03660_),
    .B1(_03710_),
    .B2(\sub1.data_o[74] ),
    .X(_03713_));
 sky130_fd_sc_hd__a31o_1 _15576_ (.A1(_03700_),
    .A2(_03709_),
    .A3(_05560_),
    .B1(_03713_),
    .X(_01739_));
 sky130_fd_sc_hd__a22o_1 _15577_ (.A1(\sub1.data_o[11] ),
    .A2(_03660_),
    .B1(_03710_),
    .B2(\sub1.data_o[75] ),
    .X(_03714_));
 sky130_fd_sc_hd__a31o_1 _15578_ (.A1(_03700_),
    .A2(_03709_),
    .A3(_05196_),
    .B1(_03714_),
    .X(_01740_));
 sky130_fd_sc_hd__a22o_1 _15579_ (.A1(\sub1.data_o[12] ),
    .A2(_03660_),
    .B1(_03710_),
    .B2(\sub1.data_o[76] ),
    .X(_03715_));
 sky130_fd_sc_hd__a31o_1 _15580_ (.A1(_03700_),
    .A2(_03709_),
    .A3(_05219_),
    .B1(_03715_),
    .X(_01741_));
 sky130_fd_sc_hd__a22o_1 _15581_ (.A1(\sub1.data_o[13] ),
    .A2(_03660_),
    .B1(_03710_),
    .B2(\sub1.data_o[77] ),
    .X(_03716_));
 sky130_fd_sc_hd__a31o_1 _15582_ (.A1(_03700_),
    .A2(_03709_),
    .A3(_05228_),
    .B1(_03716_),
    .X(_01742_));
 sky130_fd_sc_hd__clkbuf_4 _15583_ (.A(_05103_),
    .X(_03717_));
 sky130_fd_sc_hd__a22o_1 _15584_ (.A1(\sub1.data_o[14] ),
    .A2(_03660_),
    .B1(_03710_),
    .B2(\sub1.data_o[78] ),
    .X(_03718_));
 sky130_fd_sc_hd__a31o_1 _15585_ (.A1(_03717_),
    .A2(_03709_),
    .A3(_05236_),
    .B1(_03718_),
    .X(_01743_));
 sky130_fd_sc_hd__a22o_1 _15586_ (.A1(\sub1.data_o[15] ),
    .A2(_03660_),
    .B1(_03710_),
    .B2(\sub1.data_o[79] ),
    .X(_03719_));
 sky130_fd_sc_hd__a31o_1 _15587_ (.A1(_03717_),
    .A2(_03709_),
    .A3(_05245_),
    .B1(_03719_),
    .X(_01744_));
 sky130_fd_sc_hd__mux2_1 _15588_ (.A0(\mix1.data_o[0] ),
    .A1(_03170_),
    .S(\mix1.next_ready_o ),
    .X(_03720_));
 sky130_fd_sc_hd__clkbuf_1 _15589_ (.A(_03720_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _15590_ (.A0(\mix1.data_o[1] ),
    .A1(_03236_),
    .S(\mix1.next_ready_o ),
    .X(_03721_));
 sky130_fd_sc_hd__clkbuf_1 _15591_ (.A(_03721_),
    .X(_01746_));
 sky130_fd_sc_hd__mux2_1 _15592_ (.A0(\mix1.data_o[2] ),
    .A1(_03283_),
    .S(\mix1.next_ready_o ),
    .X(_03722_));
 sky130_fd_sc_hd__clkbuf_1 _15593_ (.A(_03722_),
    .X(_01747_));
 sky130_fd_sc_hd__mux2_1 _15594_ (.A0(\mix1.data_o[3] ),
    .A1(_03324_),
    .S(\mix1.next_ready_o ),
    .X(_03723_));
 sky130_fd_sc_hd__clkbuf_1 _15595_ (.A(_03723_),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_1 _15596_ (.A0(\mix1.data_o[4] ),
    .A1(_03363_),
    .S(\mix1.next_ready_o ),
    .X(_03724_));
 sky130_fd_sc_hd__clkbuf_1 _15597_ (.A(_03724_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _15598_ (.A0(\mix1.data_o[5] ),
    .A1(_03382_),
    .S(\mix1.next_ready_o ),
    .X(_03725_));
 sky130_fd_sc_hd__clkbuf_1 _15599_ (.A(_03725_),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _15600_ (.A0(\mix1.data_o[6] ),
    .A1(_03392_),
    .S(\mix1.next_ready_o ),
    .X(_03726_));
 sky130_fd_sc_hd__clkbuf_1 _15601_ (.A(_03726_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _15602_ (.A0(\mix1.data_o[7] ),
    .A1(_03402_),
    .S(\mix1.next_ready_o ),
    .X(_03727_));
 sky130_fd_sc_hd__clkbuf_1 _15603_ (.A(_03727_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _15604_ (.A0(\mix1.data_o[8] ),
    .A1(_03411_),
    .S(\mix1.next_ready_o ),
    .X(_03728_));
 sky130_fd_sc_hd__clkbuf_1 _15605_ (.A(_03728_),
    .X(_01753_));
 sky130_fd_sc_hd__buf_6 _15606_ (.A(_04379_),
    .X(_03729_));
 sky130_fd_sc_hd__clkbuf_4 _15607_ (.A(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__mux2_1 _15608_ (.A0(\mix1.data_o[9] ),
    .A1(_03424_),
    .S(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__clkbuf_1 _15609_ (.A(_03731_),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _15610_ (.A0(\mix1.data_o[10] ),
    .A1(_03435_),
    .S(_03730_),
    .X(_03732_));
 sky130_fd_sc_hd__clkbuf_1 _15611_ (.A(_03732_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _15612_ (.A0(\mix1.data_o[11] ),
    .A1(_03446_),
    .S(_03730_),
    .X(_03733_));
 sky130_fd_sc_hd__clkbuf_1 _15613_ (.A(_03733_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _15614_ (.A0(\mix1.data_o[12] ),
    .A1(_03456_),
    .S(_03730_),
    .X(_03734_));
 sky130_fd_sc_hd__clkbuf_1 _15615_ (.A(_03734_),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_1 _15616_ (.A0(\mix1.data_o[13] ),
    .A1(_03467_),
    .S(_03730_),
    .X(_03735_));
 sky130_fd_sc_hd__clkbuf_1 _15617_ (.A(_03735_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _15618_ (.A0(\mix1.data_o[14] ),
    .A1(_03477_),
    .S(_03730_),
    .X(_03736_));
 sky130_fd_sc_hd__clkbuf_1 _15619_ (.A(_03736_),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_1 _15620_ (.A0(\mix1.data_o[15] ),
    .A1(_03484_),
    .S(_03730_),
    .X(_03737_));
 sky130_fd_sc_hd__clkbuf_1 _15621_ (.A(_03737_),
    .X(_01760_));
 sky130_fd_sc_hd__mux2_1 _15622_ (.A0(\mix1.data_o[16] ),
    .A1(_03487_),
    .S(_03730_),
    .X(_03738_));
 sky130_fd_sc_hd__clkbuf_1 _15623_ (.A(_03738_),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_1 _15624_ (.A0(\mix1.data_o[17] ),
    .A1(_03491_),
    .S(_03730_),
    .X(_03739_));
 sky130_fd_sc_hd__clkbuf_1 _15625_ (.A(_03739_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _15626_ (.A0(\mix1.data_o[18] ),
    .A1(_03493_),
    .S(_03730_),
    .X(_03740_));
 sky130_fd_sc_hd__clkbuf_1 _15627_ (.A(_03740_),
    .X(_01763_));
 sky130_fd_sc_hd__buf_4 _15628_ (.A(_04379_),
    .X(_03741_));
 sky130_fd_sc_hd__clkbuf_4 _15629_ (.A(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__mux2_1 _15630_ (.A0(\mix1.data_o[19] ),
    .A1(_03497_),
    .S(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__clkbuf_1 _15631_ (.A(_03743_),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _15632_ (.A0(\mix1.data_o[20] ),
    .A1(_03502_),
    .S(_03742_),
    .X(_03744_));
 sky130_fd_sc_hd__clkbuf_1 _15633_ (.A(_03744_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _15634_ (.A0(\mix1.data_o[21] ),
    .A1(_03505_),
    .S(_03742_),
    .X(_03745_));
 sky130_fd_sc_hd__clkbuf_1 _15635_ (.A(_03745_),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _15636_ (.A0(\mix1.data_o[22] ),
    .A1(_03507_),
    .S(_03742_),
    .X(_03746_));
 sky130_fd_sc_hd__clkbuf_1 _15637_ (.A(_03746_),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _15638_ (.A0(\mix1.data_o[23] ),
    .A1(_03510_),
    .S(_03742_),
    .X(_03747_));
 sky130_fd_sc_hd__clkbuf_1 _15639_ (.A(_03747_),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _15640_ (.A0(\mix1.data_o[24] ),
    .A1(_03514_),
    .S(_03742_),
    .X(_03748_));
 sky130_fd_sc_hd__clkbuf_1 _15641_ (.A(_03748_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _15642_ (.A0(\mix1.data_o[25] ),
    .A1(_03516_),
    .S(_03742_),
    .X(_03749_));
 sky130_fd_sc_hd__clkbuf_1 _15643_ (.A(_03749_),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_1 _15644_ (.A0(\mix1.data_o[26] ),
    .A1(_03521_),
    .S(_03742_),
    .X(_03750_));
 sky130_fd_sc_hd__clkbuf_1 _15645_ (.A(_03750_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _15646_ (.A0(\mix1.data_o[27] ),
    .A1(_03525_),
    .S(_03742_),
    .X(_03751_));
 sky130_fd_sc_hd__clkbuf_1 _15647_ (.A(_03751_),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_1 _15648_ (.A0(\mix1.data_o[28] ),
    .A1(_03527_),
    .S(_03742_),
    .X(_03752_));
 sky130_fd_sc_hd__clkbuf_1 _15649_ (.A(_03752_),
    .X(_01773_));
 sky130_fd_sc_hd__buf_4 _15650_ (.A(_03741_),
    .X(_03753_));
 sky130_fd_sc_hd__mux2_1 _15651_ (.A0(\mix1.data_o[29] ),
    .A1(_03529_),
    .S(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__clkbuf_1 _15652_ (.A(_03754_),
    .X(_01774_));
 sky130_fd_sc_hd__mux2_1 _15653_ (.A0(\mix1.data_o[30] ),
    .A1(_03533_),
    .S(_03753_),
    .X(_03755_));
 sky130_fd_sc_hd__clkbuf_1 _15654_ (.A(_03755_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _15655_ (.A0(\mix1.data_o[31] ),
    .A1(_03537_),
    .S(_03753_),
    .X(_03756_));
 sky130_fd_sc_hd__clkbuf_1 _15656_ (.A(_03756_),
    .X(_01776_));
 sky130_fd_sc_hd__mux2_1 _15657_ (.A0(\mix1.data_o[32] ),
    .A1(net694),
    .S(_03753_),
    .X(_03757_));
 sky130_fd_sc_hd__clkbuf_1 _15658_ (.A(_03757_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _15659_ (.A0(\mix1.data_o[33] ),
    .A1(net772),
    .S(_03753_),
    .X(_03758_));
 sky130_fd_sc_hd__clkbuf_1 _15660_ (.A(_03758_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _15661_ (.A0(\mix1.data_o[34] ),
    .A1(net693),
    .S(_03753_),
    .X(_03759_));
 sky130_fd_sc_hd__clkbuf_1 _15662_ (.A(_03759_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _15663_ (.A0(\mix1.data_o[35] ),
    .A1(net735),
    .S(_03753_),
    .X(_03760_));
 sky130_fd_sc_hd__clkbuf_1 _15664_ (.A(_03760_),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _15665_ (.A0(\mix1.data_o[36] ),
    .A1(net700),
    .S(_03753_),
    .X(_03761_));
 sky130_fd_sc_hd__clkbuf_1 _15666_ (.A(_03761_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _15667_ (.A0(\mix1.data_o[37] ),
    .A1(net789),
    .S(_03753_),
    .X(_03762_));
 sky130_fd_sc_hd__clkbuf_1 _15668_ (.A(_03762_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _15669_ (.A0(\mix1.data_o[38] ),
    .A1(net762),
    .S(_03753_),
    .X(_03763_));
 sky130_fd_sc_hd__clkbuf_1 _15670_ (.A(_03763_),
    .X(_01783_));
 sky130_fd_sc_hd__buf_4 _15671_ (.A(_03741_),
    .X(_03764_));
 sky130_fd_sc_hd__mux2_1 _15672_ (.A0(\mix1.data_o[39] ),
    .A1(net791),
    .S(_03764_),
    .X(_03765_));
 sky130_fd_sc_hd__clkbuf_1 _15673_ (.A(_03765_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _15674_ (.A0(\mix1.data_o[40] ),
    .A1(net726),
    .S(_03764_),
    .X(_03766_));
 sky130_fd_sc_hd__clkbuf_1 _15675_ (.A(_03766_),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _15676_ (.A0(\mix1.data_o[41] ),
    .A1(net754),
    .S(_03764_),
    .X(_03767_));
 sky130_fd_sc_hd__clkbuf_1 _15677_ (.A(_03767_),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _15678_ (.A0(\mix1.data_o[42] ),
    .A1(net732),
    .S(_03764_),
    .X(_03768_));
 sky130_fd_sc_hd__clkbuf_1 _15679_ (.A(_03768_),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _15680_ (.A0(\mix1.data_o[43] ),
    .A1(net723),
    .S(_03764_),
    .X(_03769_));
 sky130_fd_sc_hd__clkbuf_1 _15681_ (.A(_03769_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _15682_ (.A0(\mix1.data_o[44] ),
    .A1(net767),
    .S(_03764_),
    .X(_03770_));
 sky130_fd_sc_hd__clkbuf_1 _15683_ (.A(_03770_),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _15684_ (.A0(\mix1.data_o[45] ),
    .A1(net718),
    .S(_03764_),
    .X(_03771_));
 sky130_fd_sc_hd__clkbuf_1 _15685_ (.A(_03771_),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _15686_ (.A0(\mix1.data_o[46] ),
    .A1(net730),
    .S(_03764_),
    .X(_03772_));
 sky130_fd_sc_hd__clkbuf_1 _15687_ (.A(_03772_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _15688_ (.A0(\mix1.data_o[47] ),
    .A1(net768),
    .S(_03764_),
    .X(_03773_));
 sky130_fd_sc_hd__clkbuf_1 _15689_ (.A(_03773_),
    .X(_01792_));
 sky130_fd_sc_hd__mux2_1 _15690_ (.A0(\mix1.data_o[48] ),
    .A1(net741),
    .S(_03764_),
    .X(_03774_));
 sky130_fd_sc_hd__clkbuf_1 _15691_ (.A(_03774_),
    .X(_01793_));
 sky130_fd_sc_hd__buf_4 _15692_ (.A(_03741_),
    .X(_03775_));
 sky130_fd_sc_hd__mux2_1 _15693_ (.A0(\mix1.data_o[49] ),
    .A1(net788),
    .S(_03775_),
    .X(_03776_));
 sky130_fd_sc_hd__clkbuf_1 _15694_ (.A(_03776_),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _15695_ (.A0(\mix1.data_o[50] ),
    .A1(net753),
    .S(_03775_),
    .X(_03777_));
 sky130_fd_sc_hd__clkbuf_1 _15696_ (.A(_03777_),
    .X(_01795_));
 sky130_fd_sc_hd__mux2_1 _15697_ (.A0(\mix1.data_o[51] ),
    .A1(net763),
    .S(_03775_),
    .X(_03778_));
 sky130_fd_sc_hd__clkbuf_1 _15698_ (.A(_03778_),
    .X(_01796_));
 sky130_fd_sc_hd__mux2_1 _15699_ (.A0(\mix1.data_o[52] ),
    .A1(net764),
    .S(_03775_),
    .X(_03779_));
 sky130_fd_sc_hd__clkbuf_1 _15700_ (.A(_03779_),
    .X(_01797_));
 sky130_fd_sc_hd__mux2_1 _15701_ (.A0(\mix1.data_o[53] ),
    .A1(net740),
    .S(_03775_),
    .X(_03780_));
 sky130_fd_sc_hd__clkbuf_1 _15702_ (.A(_03780_),
    .X(_01798_));
 sky130_fd_sc_hd__mux2_1 _15703_ (.A0(\mix1.data_o[54] ),
    .A1(net710),
    .S(_03775_),
    .X(_03781_));
 sky130_fd_sc_hd__clkbuf_1 _15704_ (.A(_03781_),
    .X(_01799_));
 sky130_fd_sc_hd__mux2_1 _15705_ (.A0(\mix1.data_o[55] ),
    .A1(net734),
    .S(_03775_),
    .X(_03782_));
 sky130_fd_sc_hd__clkbuf_1 _15706_ (.A(_03782_),
    .X(_01800_));
 sky130_fd_sc_hd__mux2_1 _15707_ (.A0(\mix1.data_o[56] ),
    .A1(net756),
    .S(_03775_),
    .X(_03783_));
 sky130_fd_sc_hd__clkbuf_1 _15708_ (.A(_03783_),
    .X(_01801_));
 sky130_fd_sc_hd__mux2_1 _15709_ (.A0(\mix1.data_o[57] ),
    .A1(net715),
    .S(_03775_),
    .X(_03784_));
 sky130_fd_sc_hd__clkbuf_1 _15710_ (.A(_03784_),
    .X(_01802_));
 sky130_fd_sc_hd__mux2_1 _15711_ (.A0(\mix1.data_o[58] ),
    .A1(net798),
    .S(_03775_),
    .X(_03785_));
 sky130_fd_sc_hd__clkbuf_1 _15712_ (.A(_03785_),
    .X(_01803_));
 sky130_fd_sc_hd__clkbuf_8 _15713_ (.A(_03741_),
    .X(_03786_));
 sky130_fd_sc_hd__mux2_1 _15714_ (.A0(\mix1.data_o[59] ),
    .A1(net743),
    .S(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__clkbuf_1 _15715_ (.A(_03787_),
    .X(_01804_));
 sky130_fd_sc_hd__mux2_1 _15716_ (.A0(\mix1.data_o[60] ),
    .A1(net742),
    .S(_03786_),
    .X(_03788_));
 sky130_fd_sc_hd__clkbuf_1 _15717_ (.A(_03788_),
    .X(_01805_));
 sky130_fd_sc_hd__mux2_1 _15718_ (.A0(\mix1.data_o[61] ),
    .A1(net724),
    .S(_03786_),
    .X(_03789_));
 sky130_fd_sc_hd__clkbuf_1 _15719_ (.A(_03789_),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _15720_ (.A0(\mix1.data_o[62] ),
    .A1(\mix1.data_reg[62] ),
    .S(_03786_),
    .X(_03790_));
 sky130_fd_sc_hd__clkbuf_1 _15721_ (.A(_03790_),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _15722_ (.A0(\mix1.data_o[63] ),
    .A1(\mix1.data_reg[63] ),
    .S(_03786_),
    .X(_03791_));
 sky130_fd_sc_hd__clkbuf_1 _15723_ (.A(_03791_),
    .X(_01808_));
 sky130_fd_sc_hd__mux2_1 _15724_ (.A0(\mix1.data_o[64] ),
    .A1(\mix1.data_reg[64] ),
    .S(_03786_),
    .X(_03792_));
 sky130_fd_sc_hd__clkbuf_1 _15725_ (.A(_03792_),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _15726_ (.A0(\mix1.data_o[65] ),
    .A1(net733),
    .S(_03786_),
    .X(_03793_));
 sky130_fd_sc_hd__clkbuf_1 _15727_ (.A(_03793_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _15728_ (.A0(\mix1.data_o[66] ),
    .A1(\mix1.data_reg[66] ),
    .S(_03786_),
    .X(_03794_));
 sky130_fd_sc_hd__clkbuf_1 _15729_ (.A(_03794_),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _15730_ (.A0(\mix1.data_o[67] ),
    .A1(\mix1.data_reg[67] ),
    .S(_03786_),
    .X(_03795_));
 sky130_fd_sc_hd__clkbuf_1 _15731_ (.A(_03795_),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _15732_ (.A0(\mix1.data_o[68] ),
    .A1(net839),
    .S(_03786_),
    .X(_03796_));
 sky130_fd_sc_hd__clkbuf_1 _15733_ (.A(_03796_),
    .X(_01813_));
 sky130_fd_sc_hd__buf_4 _15734_ (.A(_03741_),
    .X(_03797_));
 sky130_fd_sc_hd__mux2_1 _15735_ (.A0(\mix1.data_o[69] ),
    .A1(net750),
    .S(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__clkbuf_1 _15736_ (.A(_03798_),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _15737_ (.A0(\mix1.data_o[70] ),
    .A1(net697),
    .S(_03797_),
    .X(_03799_));
 sky130_fd_sc_hd__clkbuf_1 _15738_ (.A(_03799_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _15739_ (.A0(\mix1.data_o[71] ),
    .A1(net720),
    .S(_03797_),
    .X(_03800_));
 sky130_fd_sc_hd__clkbuf_1 _15740_ (.A(_03800_),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _15741_ (.A0(\mix1.data_o[72] ),
    .A1(net769),
    .S(_03797_),
    .X(_03801_));
 sky130_fd_sc_hd__clkbuf_1 _15742_ (.A(_03801_),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _15743_ (.A0(\mix1.data_o[73] ),
    .A1(net770),
    .S(_03797_),
    .X(_03802_));
 sky130_fd_sc_hd__clkbuf_1 _15744_ (.A(_03802_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _15745_ (.A0(\mix1.data_o[74] ),
    .A1(net727),
    .S(_03797_),
    .X(_03803_));
 sky130_fd_sc_hd__clkbuf_1 _15746_ (.A(_03803_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _15747_ (.A0(\mix1.data_o[75] ),
    .A1(net760),
    .S(_03797_),
    .X(_03804_));
 sky130_fd_sc_hd__clkbuf_1 _15748_ (.A(_03804_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _15749_ (.A0(\mix1.data_o[76] ),
    .A1(net777),
    .S(_03797_),
    .X(_03805_));
 sky130_fd_sc_hd__clkbuf_1 _15750_ (.A(_03805_),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _15751_ (.A0(\mix1.data_o[77] ),
    .A1(net780),
    .S(_03797_),
    .X(_03806_));
 sky130_fd_sc_hd__clkbuf_1 _15752_ (.A(_03806_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _15753_ (.A0(\mix1.data_o[78] ),
    .A1(net737),
    .S(_03797_),
    .X(_03807_));
 sky130_fd_sc_hd__clkbuf_1 _15754_ (.A(_03807_),
    .X(_01823_));
 sky130_fd_sc_hd__buf_4 _15755_ (.A(_03741_),
    .X(_03808_));
 sky130_fd_sc_hd__mux2_1 _15756_ (.A0(\mix1.data_o[79] ),
    .A1(net731),
    .S(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__clkbuf_1 _15757_ (.A(_03809_),
    .X(_01824_));
 sky130_fd_sc_hd__mux2_1 _15758_ (.A0(\mix1.data_o[80] ),
    .A1(net778),
    .S(_03808_),
    .X(_03810_));
 sky130_fd_sc_hd__clkbuf_1 _15759_ (.A(_03810_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _15760_ (.A0(\mix1.data_o[81] ),
    .A1(net755),
    .S(_03808_),
    .X(_03811_));
 sky130_fd_sc_hd__clkbuf_1 _15761_ (.A(_03811_),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _15762_ (.A0(\mix1.data_o[82] ),
    .A1(net748),
    .S(_03808_),
    .X(_03812_));
 sky130_fd_sc_hd__clkbuf_1 _15763_ (.A(_03812_),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _15764_ (.A0(\mix1.data_o[83] ),
    .A1(net786),
    .S(_03808_),
    .X(_03813_));
 sky130_fd_sc_hd__clkbuf_1 _15765_ (.A(_03813_),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _15766_ (.A0(\mix1.data_o[84] ),
    .A1(net783),
    .S(_03808_),
    .X(_03814_));
 sky130_fd_sc_hd__clkbuf_1 _15767_ (.A(_03814_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _15768_ (.A0(\mix1.data_o[85] ),
    .A1(net775),
    .S(_03808_),
    .X(_03815_));
 sky130_fd_sc_hd__clkbuf_1 _15769_ (.A(_03815_),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_1 _15770_ (.A0(\mix1.data_o[86] ),
    .A1(net792),
    .S(_03808_),
    .X(_03816_));
 sky130_fd_sc_hd__clkbuf_1 _15771_ (.A(_03816_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _15772_ (.A0(\mix1.data_o[87] ),
    .A1(net747),
    .S(_03808_),
    .X(_03817_));
 sky130_fd_sc_hd__clkbuf_1 _15773_ (.A(_03817_),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _15774_ (.A0(\mix1.data_o[88] ),
    .A1(net761),
    .S(_03808_),
    .X(_03818_));
 sky130_fd_sc_hd__clkbuf_1 _15775_ (.A(_03818_),
    .X(_01833_));
 sky130_fd_sc_hd__clkbuf_8 _15776_ (.A(_03741_),
    .X(_03819_));
 sky130_fd_sc_hd__mux2_1 _15777_ (.A0(\mix1.data_o[89] ),
    .A1(net785),
    .S(_03819_),
    .X(_03820_));
 sky130_fd_sc_hd__clkbuf_1 _15778_ (.A(_03820_),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_1 _15779_ (.A0(\mix1.data_o[90] ),
    .A1(net752),
    .S(_03819_),
    .X(_03821_));
 sky130_fd_sc_hd__clkbuf_1 _15780_ (.A(_03821_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _15781_ (.A0(\mix1.data_o[91] ),
    .A1(net736),
    .S(_03819_),
    .X(_03822_));
 sky130_fd_sc_hd__clkbuf_1 _15782_ (.A(_03822_),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _15783_ (.A0(\mix1.data_o[92] ),
    .A1(net782),
    .S(_03819_),
    .X(_03823_));
 sky130_fd_sc_hd__clkbuf_1 _15784_ (.A(_03823_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _15785_ (.A0(\mix1.data_o[93] ),
    .A1(net773),
    .S(_03819_),
    .X(_03824_));
 sky130_fd_sc_hd__clkbuf_1 _15786_ (.A(_03824_),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _15787_ (.A0(\mix1.data_o[94] ),
    .A1(net716),
    .S(_03819_),
    .X(_03825_));
 sky130_fd_sc_hd__clkbuf_1 _15788_ (.A(_03825_),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _15789_ (.A0(\mix1.data_o[95] ),
    .A1(net725),
    .S(_03819_),
    .X(_03826_));
 sky130_fd_sc_hd__clkbuf_1 _15790_ (.A(_03826_),
    .X(_01840_));
 sky130_fd_sc_hd__mux2_1 _15791_ (.A0(\mix1.data_o[96] ),
    .A1(net739),
    .S(_03819_),
    .X(_03827_));
 sky130_fd_sc_hd__clkbuf_1 _15792_ (.A(_03827_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _15793_ (.A0(\mix1.data_o[97] ),
    .A1(net759),
    .S(_03819_),
    .X(_03828_));
 sky130_fd_sc_hd__clkbuf_1 _15794_ (.A(_03828_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _15795_ (.A0(\mix1.data_o[98] ),
    .A1(net722),
    .S(_03819_),
    .X(_03829_));
 sky130_fd_sc_hd__clkbuf_1 _15796_ (.A(_03829_),
    .X(_01843_));
 sky130_fd_sc_hd__buf_4 _15797_ (.A(_03741_),
    .X(_03830_));
 sky130_fd_sc_hd__mux2_1 _15798_ (.A0(\mix1.data_o[99] ),
    .A1(net719),
    .S(_03830_),
    .X(_03831_));
 sky130_fd_sc_hd__clkbuf_1 _15799_ (.A(_03831_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _15800_ (.A0(\mix1.data_o[100] ),
    .A1(net709),
    .S(_03830_),
    .X(_03832_));
 sky130_fd_sc_hd__clkbuf_1 _15801_ (.A(_03832_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _15802_ (.A0(\mix1.data_o[101] ),
    .A1(net784),
    .S(_03830_),
    .X(_03833_));
 sky130_fd_sc_hd__clkbuf_1 _15803_ (.A(_03833_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _15804_ (.A0(\mix1.data_o[102] ),
    .A1(net717),
    .S(_03830_),
    .X(_03834_));
 sky130_fd_sc_hd__clkbuf_1 _15805_ (.A(_03834_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _15806_ (.A0(\mix1.data_o[103] ),
    .A1(net728),
    .S(_03830_),
    .X(_03835_));
 sky130_fd_sc_hd__clkbuf_1 _15807_ (.A(_03835_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _15808_ (.A0(\mix1.data_o[104] ),
    .A1(net781),
    .S(_03830_),
    .X(_03836_));
 sky130_fd_sc_hd__clkbuf_1 _15809_ (.A(_03836_),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _15810_ (.A0(\mix1.data_o[105] ),
    .A1(net687),
    .S(_03830_),
    .X(_03837_));
 sky130_fd_sc_hd__clkbuf_1 _15811_ (.A(_03837_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _15812_ (.A0(\mix1.data_o[106] ),
    .A1(net751),
    .S(_03830_),
    .X(_03838_));
 sky130_fd_sc_hd__clkbuf_1 _15813_ (.A(_03838_),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _15814_ (.A0(\mix1.data_o[107] ),
    .A1(net746),
    .S(_03830_),
    .X(_03839_));
 sky130_fd_sc_hd__clkbuf_1 _15815_ (.A(_03839_),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _15816_ (.A0(\mix1.data_o[108] ),
    .A1(net758),
    .S(_03830_),
    .X(_03840_));
 sky130_fd_sc_hd__clkbuf_1 _15817_ (.A(_03840_),
    .X(_01853_));
 sky130_fd_sc_hd__clkbuf_8 _15818_ (.A(_03741_),
    .X(_03841_));
 sky130_fd_sc_hd__mux2_1 _15819_ (.A0(\mix1.data_o[109] ),
    .A1(net787),
    .S(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__clkbuf_1 _15820_ (.A(_03842_),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _15821_ (.A0(\mix1.data_o[110] ),
    .A1(net711),
    .S(_03841_),
    .X(_03843_));
 sky130_fd_sc_hd__clkbuf_1 _15822_ (.A(_03843_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _15823_ (.A0(\mix1.data_o[111] ),
    .A1(net745),
    .S(_03841_),
    .X(_03844_));
 sky130_fd_sc_hd__clkbuf_1 _15824_ (.A(_03844_),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_1 _15825_ (.A0(\mix1.data_o[112] ),
    .A1(net771),
    .S(_03841_),
    .X(_03845_));
 sky130_fd_sc_hd__clkbuf_1 _15826_ (.A(_03845_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _15827_ (.A0(\mix1.data_o[113] ),
    .A1(net738),
    .S(_03841_),
    .X(_03846_));
 sky130_fd_sc_hd__clkbuf_1 _15828_ (.A(_03846_),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _15829_ (.A0(\mix1.data_o[114] ),
    .A1(net749),
    .S(_03841_),
    .X(_03847_));
 sky130_fd_sc_hd__clkbuf_1 _15830_ (.A(_03847_),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _15831_ (.A0(\mix1.data_o[115] ),
    .A1(net696),
    .S(_03841_),
    .X(_03848_));
 sky130_fd_sc_hd__clkbuf_1 _15832_ (.A(_03848_),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _15833_ (.A0(\mix1.data_o[116] ),
    .A1(net688),
    .S(_03841_),
    .X(_03849_));
 sky130_fd_sc_hd__clkbuf_1 _15834_ (.A(_03849_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _15835_ (.A0(\mix1.data_o[117] ),
    .A1(net776),
    .S(_03841_),
    .X(_03850_));
 sky130_fd_sc_hd__clkbuf_1 _15836_ (.A(_03850_),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _15837_ (.A0(\mix1.data_o[118] ),
    .A1(net779),
    .S(_03841_),
    .X(_03851_));
 sky130_fd_sc_hd__clkbuf_1 _15838_ (.A(_03851_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _15839_ (.A0(\mix1.data_o[119] ),
    .A1(net790),
    .S(_03729_),
    .X(_03852_));
 sky130_fd_sc_hd__clkbuf_1 _15840_ (.A(_03852_),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _15841_ (.A0(\mix1.data_o[120] ),
    .A1(net744),
    .S(_03729_),
    .X(_03853_));
 sky130_fd_sc_hd__clkbuf_1 _15842_ (.A(_03853_),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _15843_ (.A0(\mix1.data_o[121] ),
    .A1(net757),
    .S(_03729_),
    .X(_03854_));
 sky130_fd_sc_hd__clkbuf_1 _15844_ (.A(_03854_),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _15845_ (.A0(\mix1.data_o[122] ),
    .A1(net684),
    .S(_03729_),
    .X(_03855_));
 sky130_fd_sc_hd__clkbuf_1 _15846_ (.A(_03855_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _15847_ (.A0(\mix1.data_o[123] ),
    .A1(net774),
    .S(_03729_),
    .X(_03856_));
 sky130_fd_sc_hd__clkbuf_1 _15848_ (.A(_03856_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _15849_ (.A0(\mix1.data_o[124] ),
    .A1(net766),
    .S(_03729_),
    .X(_03857_));
 sky130_fd_sc_hd__clkbuf_1 _15850_ (.A(_03857_),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _15851_ (.A0(\mix1.data_o[125] ),
    .A1(net729),
    .S(_03729_),
    .X(_03858_));
 sky130_fd_sc_hd__clkbuf_1 _15852_ (.A(_03858_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _15853_ (.A0(\mix1.data_o[126] ),
    .A1(net765),
    .S(_03729_),
    .X(_03859_));
 sky130_fd_sc_hd__clkbuf_1 _15854_ (.A(_03859_),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _15855_ (.A0(\mix1.data_o[127] ),
    .A1(net706),
    .S(_03729_),
    .X(_03860_));
 sky130_fd_sc_hd__clkbuf_1 _15856_ (.A(_03860_),
    .X(_01872_));
 sky130_fd_sc_hd__or4_1 _15857_ (.A(_04362_),
    .B(_04363_),
    .C(_04364_),
    .D(_04365_),
    .X(_03861_));
 sky130_fd_sc_hd__or2_1 _15858_ (.A(\sub1.state[4] ),
    .B(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__o211a_1 _15859_ (.A1(_04652_),
    .A2(_03862_),
    .B1(_04673_),
    .C1(_05104_),
    .X(_01873_));
 sky130_fd_sc_hd__nand2_1 _15860_ (.A(_04705_),
    .B(_04680_),
    .Y(_01874_));
 sky130_fd_sc_hd__xnor2_1 _15861_ (.A(_04365_),
    .B(_04700_),
    .Y(_01875_));
 sky130_fd_sc_hd__a21boi_1 _15862_ (.A1(_04365_),
    .A2(_04687_),
    .B1_N(_04364_),
    .Y(_03863_));
 sky130_fd_sc_hd__or2_1 _15863_ (.A(_03709_),
    .B(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__clkbuf_1 _15864_ (.A(_03864_),
    .X(_01876_));
 sky130_fd_sc_hd__o21ai_1 _15865_ (.A1(net675),
    .A2(_03593_),
    .B1(_03861_),
    .Y(_03865_));
 sky130_fd_sc_hd__a21oi_1 _15866_ (.A1(net675),
    .A2(_03593_),
    .B1(_03865_),
    .Y(_01877_));
 sky130_fd_sc_hd__mux2_1 _15867_ (.A0(\sub1.data_o[88] ),
    .A1(_05547_),
    .S(_04888_),
    .X(_03866_));
 sky130_fd_sc_hd__clkbuf_1 _15868_ (.A(_03866_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _15869_ (.A0(\sub1.data_o[89] ),
    .A1(_05553_),
    .S(_04888_),
    .X(_03867_));
 sky130_fd_sc_hd__clkbuf_1 _15870_ (.A(_03867_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _15871_ (.A0(\sub1.data_o[90] ),
    .A1(_05559_),
    .S(_04888_),
    .X(_03868_));
 sky130_fd_sc_hd__clkbuf_1 _15872_ (.A(_03868_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _15873_ (.A0(\sub1.data_o[91] ),
    .A1(_05195_),
    .S(_04888_),
    .X(_03869_));
 sky130_fd_sc_hd__clkbuf_1 _15874_ (.A(_03869_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _15875_ (.A0(\sub1.data_o[92] ),
    .A1(_05218_),
    .S(_04888_),
    .X(_03870_));
 sky130_fd_sc_hd__clkbuf_1 _15876_ (.A(_03870_),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _15877_ (.A0(\sub1.data_o[93] ),
    .A1(_05227_),
    .S(_04888_),
    .X(_03871_));
 sky130_fd_sc_hd__clkbuf_1 _15878_ (.A(_03871_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _15879_ (.A0(\sub1.data_o[94] ),
    .A1(_05235_),
    .S(_04888_),
    .X(_03872_));
 sky130_fd_sc_hd__clkbuf_1 _15880_ (.A(_03872_),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _15881_ (.A0(\sub1.data_o[95] ),
    .A1(_05244_),
    .S(_04888_),
    .X(_03873_));
 sky130_fd_sc_hd__clkbuf_1 _15882_ (.A(_03873_),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _15883_ (.A0(_05547_),
    .A1(\sub1.data_o[64] ),
    .S(_05200_),
    .X(_03874_));
 sky130_fd_sc_hd__or2_1 _15884_ (.A(_04368_),
    .B(_04716_),
    .X(_03875_));
 sky130_fd_sc_hd__clkbuf_4 _15885_ (.A(_03875_),
    .X(_03876_));
 sky130_fd_sc_hd__mux2_1 _15886_ (.A0(\sub1.data_o[96] ),
    .A1(_03874_),
    .S(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__clkbuf_1 _15887_ (.A(_03877_),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _15888_ (.A0(_05553_),
    .A1(\sub1.data_o[65] ),
    .S(_05200_),
    .X(_03878_));
 sky130_fd_sc_hd__mux2_1 _15889_ (.A0(\sub1.data_o[97] ),
    .A1(_03878_),
    .S(_03876_),
    .X(_03879_));
 sky130_fd_sc_hd__clkbuf_1 _15890_ (.A(_03879_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _15891_ (.A0(_05559_),
    .A1(\sub1.data_o[66] ),
    .S(_05200_),
    .X(_03880_));
 sky130_fd_sc_hd__mux2_1 _15892_ (.A0(\sub1.data_o[98] ),
    .A1(_03880_),
    .S(_03876_),
    .X(_03881_));
 sky130_fd_sc_hd__clkbuf_1 _15893_ (.A(_03881_),
    .X(_01888_));
 sky130_fd_sc_hd__mux2_1 _15894_ (.A0(_05195_),
    .A1(\sub1.data_o[67] ),
    .S(_05200_),
    .X(_03882_));
 sky130_fd_sc_hd__mux2_1 _15895_ (.A0(\sub1.data_o[99] ),
    .A1(_03882_),
    .S(_03876_),
    .X(_03883_));
 sky130_fd_sc_hd__clkbuf_1 _15896_ (.A(_03883_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _15897_ (.A0(_05218_),
    .A1(\sub1.data_o[68] ),
    .S(_05200_),
    .X(_03884_));
 sky130_fd_sc_hd__mux2_1 _15898_ (.A0(\sub1.data_o[100] ),
    .A1(_03884_),
    .S(_03876_),
    .X(_03885_));
 sky130_fd_sc_hd__clkbuf_1 _15899_ (.A(_03885_),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _15900_ (.A0(_05227_),
    .A1(\sub1.data_o[69] ),
    .S(_05199_),
    .X(_03886_));
 sky130_fd_sc_hd__mux2_1 _15901_ (.A0(\sub1.data_o[101] ),
    .A1(_03886_),
    .S(_03876_),
    .X(_03887_));
 sky130_fd_sc_hd__clkbuf_1 _15902_ (.A(_03887_),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _15903_ (.A0(_05235_),
    .A1(\sub1.data_o[70] ),
    .S(_05199_),
    .X(_03888_));
 sky130_fd_sc_hd__mux2_1 _15904_ (.A0(\sub1.data_o[102] ),
    .A1(_03888_),
    .S(_03876_),
    .X(_03889_));
 sky130_fd_sc_hd__clkbuf_1 _15905_ (.A(_03889_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _15906_ (.A0(_05244_),
    .A1(\sub1.data_o[71] ),
    .S(_05199_),
    .X(_03890_));
 sky130_fd_sc_hd__mux2_1 _15907_ (.A0(\sub1.data_o[103] ),
    .A1(_03890_),
    .S(_03876_),
    .X(_03891_));
 sky130_fd_sc_hd__clkbuf_1 _15908_ (.A(_03891_),
    .X(_01893_));
 sky130_fd_sc_hd__nor2_2 _15909_ (.A(_04369_),
    .B(_04943_),
    .Y(_03892_));
 sky130_fd_sc_hd__a22o_1 _15910_ (.A1(\sub1.data_o[40] ),
    .A2(_03576_),
    .B1(_03892_),
    .B2(\sub1.data_o[104] ),
    .X(_03893_));
 sky130_fd_sc_hd__a31o_1 _15911_ (.A1(_03717_),
    .A2(_04943_),
    .A3(_05548_),
    .B1(_03893_),
    .X(_01894_));
 sky130_fd_sc_hd__a22o_1 _15912_ (.A1(\sub1.data_o[41] ),
    .A2(_03576_),
    .B1(_03892_),
    .B2(\sub1.data_o[105] ),
    .X(_03894_));
 sky130_fd_sc_hd__a31o_1 _15913_ (.A1(_03717_),
    .A2(_04943_),
    .A3(_05554_),
    .B1(_03894_),
    .X(_01895_));
 sky130_fd_sc_hd__a22o_1 _15914_ (.A1(\sub1.data_o[42] ),
    .A2(_03576_),
    .B1(_03892_),
    .B2(\sub1.data_o[106] ),
    .X(_03895_));
 sky130_fd_sc_hd__a31o_1 _15915_ (.A1(_03717_),
    .A2(_04943_),
    .A3(_05560_),
    .B1(_03895_),
    .X(_01896_));
 sky130_fd_sc_hd__a22o_1 _15916_ (.A1(\sub1.data_o[43] ),
    .A2(_03576_),
    .B1(_03892_),
    .B2(\sub1.data_o[107] ),
    .X(_03896_));
 sky130_fd_sc_hd__a31o_1 _15917_ (.A1(_03717_),
    .A2(_04943_),
    .A3(_05196_),
    .B1(_03896_),
    .X(_01897_));
 sky130_fd_sc_hd__a22o_1 _15918_ (.A1(\sub1.data_o[44] ),
    .A2(_03576_),
    .B1(_03892_),
    .B2(\sub1.data_o[108] ),
    .X(_03897_));
 sky130_fd_sc_hd__a31o_1 _15919_ (.A1(_03717_),
    .A2(_04943_),
    .A3(_05219_),
    .B1(_03897_),
    .X(_01898_));
 sky130_fd_sc_hd__a22o_1 _15920_ (.A1(\sub1.data_o[45] ),
    .A2(_03576_),
    .B1(_03892_),
    .B2(\sub1.data_o[109] ),
    .X(_03898_));
 sky130_fd_sc_hd__a31o_1 _15921_ (.A1(_03717_),
    .A2(_04943_),
    .A3(_05228_),
    .B1(_03898_),
    .X(_01899_));
 sky130_fd_sc_hd__a22o_1 _15922_ (.A1(\sub1.data_o[46] ),
    .A2(_03576_),
    .B1(_03892_),
    .B2(\sub1.data_o[110] ),
    .X(_03899_));
 sky130_fd_sc_hd__a31o_1 _15923_ (.A1(_03717_),
    .A2(_04943_),
    .A3(_05236_),
    .B1(_03899_),
    .X(_01900_));
 sky130_fd_sc_hd__a22o_1 _15924_ (.A1(\sub1.data_o[47] ),
    .A2(_03576_),
    .B1(_03892_),
    .B2(\sub1.data_o[111] ),
    .X(_03900_));
 sky130_fd_sc_hd__a31o_1 _15925_ (.A1(_03717_),
    .A2(_04943_),
    .A3(_05245_),
    .B1(_03900_),
    .X(_01901_));
 sky130_fd_sc_hd__clkbuf_4 _15926_ (.A(_04371_),
    .X(_03901_));
 sky130_fd_sc_hd__buf_4 _15927_ (.A(_04742_),
    .X(_03902_));
 sky130_fd_sc_hd__mux2_1 _15928_ (.A0(net253),
    .A1(\ks1.key_reg[96] ),
    .S(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__xor2_1 _15929_ (.A(\ks1.col[0] ),
    .B(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__buf_4 _15930_ (.A(_04742_),
    .X(_03905_));
 sky130_fd_sc_hd__buf_4 _15931_ (.A(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__buf_4 _15932_ (.A(_03906_),
    .X(_03907_));
 sky130_fd_sc_hd__mux2_1 _15933_ (.A0(net218),
    .A1(\ks1.key_reg[64] ),
    .S(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__xor2_1 _15934_ (.A(_03904_),
    .B(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__buf_4 _15935_ (.A(_03907_),
    .X(_03910_));
 sky130_fd_sc_hd__mux2_1 _15936_ (.A0(net183),
    .A1(\ks1.key_reg[32] ),
    .S(_03910_),
    .X(_03911_));
 sky130_fd_sc_hd__xor2_1 _15937_ (.A(_03909_),
    .B(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__or2_1 _15938_ (.A(_04920_),
    .B(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__buf_4 _15939_ (.A(_04371_),
    .X(_03914_));
 sky130_fd_sc_hd__a21oi_1 _15940_ (.A1(_04920_),
    .A2(_03912_),
    .B1(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__a22o_1 _15941_ (.A1(net704),
    .A2(_03901_),
    .B1(_03913_),
    .B2(_03915_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_2 _15942_ (.A0(net254),
    .A1(\ks1.key_reg[97] ),
    .S(_03902_),
    .X(_03916_));
 sky130_fd_sc_hd__xor2_4 _15943_ (.A(\ks1.col[1] ),
    .B(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__buf_4 _15944_ (.A(_03905_),
    .X(_03918_));
 sky130_fd_sc_hd__mux2_1 _15945_ (.A0(net219),
    .A1(\ks1.key_reg[65] ),
    .S(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__xor2_2 _15946_ (.A(_03917_),
    .B(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__mux2_1 _15947_ (.A0(net184),
    .A1(\ks1.key_reg[33] ),
    .S(_03910_),
    .X(_03921_));
 sky130_fd_sc_hd__xor2_2 _15948_ (.A(_03920_),
    .B(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__and2_1 _15949_ (.A(_04759_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__o21ai_1 _15950_ (.A1(_04759_),
    .A2(_03922_),
    .B1(_04373_),
    .Y(_03924_));
 sky130_fd_sc_hd__o22a_1 _15951_ (.A1(net703),
    .A2(\ks1.next_ready_o ),
    .B1(_03923_),
    .B2(_03924_),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_2 _15952_ (.A0(net255),
    .A1(\ks1.key_reg[98] ),
    .S(_03902_),
    .X(_03925_));
 sky130_fd_sc_hd__xor2_4 _15953_ (.A(\ks1.col[2] ),
    .B(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__mux2_1 _15954_ (.A0(net220),
    .A1(\ks1.key_reg[66] ),
    .S(_03907_),
    .X(_03927_));
 sky130_fd_sc_hd__xor2_1 _15955_ (.A(_03926_),
    .B(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__mux2_1 _15956_ (.A0(net185),
    .A1(\ks1.key_reg[34] ),
    .S(_03910_),
    .X(_03929_));
 sky130_fd_sc_hd__xor2_1 _15957_ (.A(_03928_),
    .B(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__or2_1 _15958_ (.A(_05050_),
    .B(_03930_),
    .X(_03931_));
 sky130_fd_sc_hd__a21oi_1 _15959_ (.A1(_05050_),
    .A2(_03930_),
    .B1(_03914_),
    .Y(_03932_));
 sky130_fd_sc_hd__a22o_1 _15960_ (.A1(net691),
    .A2(_03901_),
    .B1(_03931_),
    .B2(_03932_),
    .X(_01904_));
 sky130_fd_sc_hd__mux2_2 _15961_ (.A0(net256),
    .A1(\ks1.key_reg[99] ),
    .S(_03905_),
    .X(_03933_));
 sky130_fd_sc_hd__xor2_4 _15962_ (.A(\ks1.col[3] ),
    .B(_03933_),
    .X(_03934_));
 sky130_fd_sc_hd__mux2_1 _15963_ (.A0(net221),
    .A1(\ks1.key_reg[67] ),
    .S(_03918_),
    .X(_03935_));
 sky130_fd_sc_hd__xor2_2 _15964_ (.A(_03934_),
    .B(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__buf_4 _15965_ (.A(_03918_),
    .X(_03937_));
 sky130_fd_sc_hd__mux2_1 _15966_ (.A0(net186),
    .A1(\ks1.key_reg[35] ),
    .S(_03937_),
    .X(_03938_));
 sky130_fd_sc_hd__xor2_2 _15967_ (.A(_03936_),
    .B(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__xnor2_1 _15968_ (.A(_04800_),
    .B(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__mux2_1 _15969_ (.A0(\ks1.key_reg[3] ),
    .A1(_03940_),
    .S(_04373_),
    .X(_03941_));
 sky130_fd_sc_hd__clkbuf_1 _15970_ (.A(_03941_),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_2 _15971_ (.A0(net131),
    .A1(\ks1.key_reg[100] ),
    .S(_03905_),
    .X(_03942_));
 sky130_fd_sc_hd__xor2_4 _15972_ (.A(\ks1.col[4] ),
    .B(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__mux2_1 _15973_ (.A0(net222),
    .A1(\ks1.key_reg[68] ),
    .S(_03906_),
    .X(_03944_));
 sky130_fd_sc_hd__xor2_2 _15974_ (.A(_03943_),
    .B(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__mux2_1 _15975_ (.A0(net187),
    .A1(\ks1.key_reg[36] ),
    .S(_03937_),
    .X(_03946_));
 sky130_fd_sc_hd__xor2_2 _15976_ (.A(_03945_),
    .B(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__xnor2_1 _15977_ (.A(_04734_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__mux2_1 _15978_ (.A0(\ks1.key_reg[4] ),
    .A1(_03948_),
    .S(_04373_),
    .X(_03949_));
 sky130_fd_sc_hd__clkbuf_1 _15979_ (.A(_03949_),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_2 _15980_ (.A0(net132),
    .A1(\ks1.key_reg[101] ),
    .S(_03905_),
    .X(_03950_));
 sky130_fd_sc_hd__xor2_4 _15981_ (.A(\ks1.col[5] ),
    .B(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__mux2_2 _15982_ (.A0(net223),
    .A1(\ks1.key_reg[69] ),
    .S(_03906_),
    .X(_03952_));
 sky130_fd_sc_hd__xor2_4 _15983_ (.A(_03951_),
    .B(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__mux2_1 _15984_ (.A0(net188),
    .A1(\ks1.key_reg[37] ),
    .S(_03937_),
    .X(_03954_));
 sky130_fd_sc_hd__xor2_2 _15985_ (.A(_03953_),
    .B(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__xnor2_1 _15986_ (.A(_04961_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__buf_4 _15987_ (.A(_04372_),
    .X(_03957_));
 sky130_fd_sc_hd__buf_4 _15988_ (.A(_03957_),
    .X(_03958_));
 sky130_fd_sc_hd__mux2_1 _15989_ (.A0(\ks1.key_reg[5] ),
    .A1(_03956_),
    .S(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__clkbuf_1 _15990_ (.A(_03959_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_2 _15991_ (.A0(net133),
    .A1(\ks1.key_reg[102] ),
    .S(_03902_),
    .X(_03960_));
 sky130_fd_sc_hd__xor2_4 _15992_ (.A(\ks1.col[6] ),
    .B(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__mux2_2 _15993_ (.A0(net225),
    .A1(\ks1.key_reg[70] ),
    .S(_03907_),
    .X(_03962_));
 sky130_fd_sc_hd__xor2_4 _15994_ (.A(_03961_),
    .B(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__mux2_2 _15995_ (.A0(net189),
    .A1(\ks1.key_reg[38] ),
    .S(_03910_),
    .X(_03964_));
 sky130_fd_sc_hd__xor2_4 _15996_ (.A(_03963_),
    .B(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__or2_1 _15997_ (.A(_04865_),
    .B(_03965_),
    .X(_03966_));
 sky130_fd_sc_hd__a21oi_1 _15998_ (.A1(_04865_),
    .A2(_03965_),
    .B1(_03914_),
    .Y(_03967_));
 sky130_fd_sc_hd__a22o_1 _15999_ (.A1(net702),
    .A2(_03901_),
    .B1(_03966_),
    .B2(_03967_),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_2 _16000_ (.A0(net134),
    .A1(\ks1.key_reg[103] ),
    .S(_03902_),
    .X(_03968_));
 sky130_fd_sc_hd__xor2_4 _16001_ (.A(\ks1.col[7] ),
    .B(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__mux2_2 _16002_ (.A0(net226),
    .A1(\ks1.key_reg[71] ),
    .S(_03907_),
    .X(_03970_));
 sky130_fd_sc_hd__xor2_4 _16003_ (.A(_03969_),
    .B(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__mux2_1 _16004_ (.A0(net190),
    .A1(\ks1.key_reg[39] ),
    .S(_03910_),
    .X(_03972_));
 sky130_fd_sc_hd__xor2_2 _16005_ (.A(_03971_),
    .B(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__or2_1 _16006_ (.A(_05007_),
    .B(_03973_),
    .X(_03974_));
 sky130_fd_sc_hd__a21oi_1 _16007_ (.A1(_05007_),
    .A2(_03973_),
    .B1(_03914_),
    .Y(_03975_));
 sky130_fd_sc_hd__a22o_1 _16008_ (.A1(net713),
    .A2(_03901_),
    .B1(_03974_),
    .B2(_03975_),
    .X(_01909_));
 sky130_fd_sc_hd__buf_4 _16009_ (.A(_04742_),
    .X(_03976_));
 sky130_fd_sc_hd__mux2_1 _16010_ (.A0(net135),
    .A1(\ks1.key_reg[104] ),
    .S(_03976_),
    .X(_03977_));
 sky130_fd_sc_hd__xor2_2 _16011_ (.A(_05547_),
    .B(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__buf_4 _16012_ (.A(_03905_),
    .X(_03979_));
 sky130_fd_sc_hd__mux2_1 _16013_ (.A0(net227),
    .A1(\ks1.key_reg[72] ),
    .S(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__xor2_2 _16014_ (.A(_03978_),
    .B(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__buf_4 _16015_ (.A(_03918_),
    .X(_03982_));
 sky130_fd_sc_hd__mux2_1 _16016_ (.A0(net192),
    .A1(\ks1.key_reg[40] ),
    .S(_03982_),
    .X(_03983_));
 sky130_fd_sc_hd__xnor2_1 _16017_ (.A(_03981_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__xnor2_1 _16018_ (.A(_04913_),
    .B(_03984_),
    .Y(_03985_));
 sky130_fd_sc_hd__mux2_1 _16019_ (.A0(\ks1.key_reg[8] ),
    .A1(_03985_),
    .S(_03958_),
    .X(_03986_));
 sky130_fd_sc_hd__clkbuf_1 _16020_ (.A(_03986_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _16021_ (.A0(net228),
    .A1(\ks1.key_reg[73] ),
    .S(_03979_),
    .X(_03987_));
 sky130_fd_sc_hd__mux2_1 _16022_ (.A0(net136),
    .A1(\ks1.key_reg[105] ),
    .S(_03976_),
    .X(_03988_));
 sky130_fd_sc_hd__xnor2_2 _16023_ (.A(_05553_),
    .B(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__xnor2_2 _16024_ (.A(_03987_),
    .B(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__mux2_1 _16025_ (.A0(net193),
    .A1(\ks1.key_reg[41] ),
    .S(_03982_),
    .X(_03991_));
 sky130_fd_sc_hd__xnor2_2 _16026_ (.A(_03990_),
    .B(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__xor2_1 _16027_ (.A(_04757_),
    .B(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__mux2_1 _16028_ (.A0(\ks1.key_reg[9] ),
    .A1(_03993_),
    .S(_03958_),
    .X(_03994_));
 sky130_fd_sc_hd__clkbuf_1 _16029_ (.A(_03994_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _16030_ (.A0(net194),
    .A1(\ks1.key_reg[42] ),
    .S(_03910_),
    .X(_03995_));
 sky130_fd_sc_hd__mux2_1 _16031_ (.A0(net229),
    .A1(\ks1.key_reg[74] ),
    .S(_03907_),
    .X(_03996_));
 sky130_fd_sc_hd__mux2_1 _16032_ (.A0(net137),
    .A1(\ks1.key_reg[106] ),
    .S(_03979_),
    .X(_03997_));
 sky130_fd_sc_hd__xor2_2 _16033_ (.A(_05559_),
    .B(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__xor2_2 _16034_ (.A(_03996_),
    .B(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__xor2_2 _16035_ (.A(_03995_),
    .B(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__nor2_1 _16036_ (.A(_05048_),
    .B(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__a21o_1 _16037_ (.A1(_05048_),
    .A2(_04000_),
    .B1(_04371_),
    .X(_04002_));
 sky130_fd_sc_hd__o22a_1 _16038_ (.A1(net708),
    .A2(\ks1.next_ready_o ),
    .B1(_04001_),
    .B2(_04002_),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _16039_ (.A0(net195),
    .A1(\ks1.key_reg[43] ),
    .S(_03910_),
    .X(_04003_));
 sky130_fd_sc_hd__mux2_1 _16040_ (.A0(net230),
    .A1(\ks1.key_reg[75] ),
    .S(_03918_),
    .X(_04004_));
 sky130_fd_sc_hd__mux2_2 _16041_ (.A0(net138),
    .A1(\ks1.key_reg[107] ),
    .S(_03902_),
    .X(_04005_));
 sky130_fd_sc_hd__xor2_4 _16042_ (.A(_05195_),
    .B(_04005_),
    .X(_04006_));
 sky130_fd_sc_hd__xnor2_2 _16043_ (.A(_04004_),
    .B(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__xnor2_2 _16044_ (.A(_04003_),
    .B(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__or2_1 _16045_ (.A(_04798_),
    .B(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__a21oi_1 _16046_ (.A1(_04798_),
    .A2(_04008_),
    .B1(_03914_),
    .Y(_04010_));
 sky130_fd_sc_hd__a22o_1 _16047_ (.A1(net707),
    .A2(_03901_),
    .B1(_04009_),
    .B2(_04010_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _16048_ (.A0(net139),
    .A1(\ks1.key_reg[108] ),
    .S(_04742_),
    .X(_04011_));
 sky130_fd_sc_hd__xnor2_2 _16049_ (.A(_05218_),
    .B(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__mux2_1 _16050_ (.A0(net231),
    .A1(\ks1.key_reg[76] ),
    .S(_03979_),
    .X(_04013_));
 sky130_fd_sc_hd__xnor2_2 _16051_ (.A(_04012_),
    .B(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hd__mux2_1 _16052_ (.A0(net196),
    .A1(\ks1.key_reg[44] ),
    .S(_03907_),
    .X(_04015_));
 sky130_fd_sc_hd__xnor2_2 _16053_ (.A(_04014_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__xnor2_1 _16054_ (.A(_04736_),
    .B(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__mux2_1 _16055_ (.A0(\ks1.key_reg[12] ),
    .A1(_04017_),
    .S(_03958_),
    .X(_04018_));
 sky130_fd_sc_hd__clkbuf_1 _16056_ (.A(_04018_),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _16057_ (.A0(net197),
    .A1(\ks1.key_reg[45] ),
    .S(_03982_),
    .X(_04019_));
 sky130_fd_sc_hd__mux2_1 _16058_ (.A0(net232),
    .A1(\ks1.key_reg[77] ),
    .S(_03918_),
    .X(_04020_));
 sky130_fd_sc_hd__mux2_1 _16059_ (.A0(net140),
    .A1(\ks1.key_reg[109] ),
    .S(_03905_),
    .X(_04021_));
 sky130_fd_sc_hd__xnor2_2 _16060_ (.A(_05227_),
    .B(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__xnor2_2 _16061_ (.A(_04020_),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__xnor2_2 _16062_ (.A(_04019_),
    .B(_04023_),
    .Y(_04024_));
 sky130_fd_sc_hd__nor2_1 _16063_ (.A(_04959_),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__a21o_1 _16064_ (.A1(_04959_),
    .A2(_04024_),
    .B1(_04371_),
    .X(_04026_));
 sky130_fd_sc_hd__o22a_1 _16065_ (.A1(net695),
    .A2(\ks1.next_ready_o ),
    .B1(_04025_),
    .B2(_04026_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_2 _16066_ (.A0(net142),
    .A1(\ks1.key_reg[110] ),
    .S(_03979_),
    .X(_04027_));
 sky130_fd_sc_hd__xor2_4 _16067_ (.A(_05235_),
    .B(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__mux2_2 _16068_ (.A0(net233),
    .A1(\ks1.key_reg[78] ),
    .S(_03907_),
    .X(_04029_));
 sky130_fd_sc_hd__xor2_4 _16069_ (.A(_04028_),
    .B(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__mux2_2 _16070_ (.A0(net198),
    .A1(\ks1.key_reg[46] ),
    .S(_03910_),
    .X(_04031_));
 sky130_fd_sc_hd__xor2_4 _16071_ (.A(_04030_),
    .B(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__nor2_1 _16072_ (.A(_04862_),
    .B(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__a21o_1 _16073_ (.A1(_04862_),
    .A2(_04032_),
    .B1(_04371_),
    .X(_04034_));
 sky130_fd_sc_hd__o22a_1 _16074_ (.A1(net699),
    .A2(\ks1.next_ready_o ),
    .B1(_04033_),
    .B2(_04034_),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_1 _16075_ (.A0(net199),
    .A1(\ks1.key_reg[47] ),
    .S(_03982_),
    .X(_04035_));
 sky130_fd_sc_hd__mux2_1 _16076_ (.A0(net234),
    .A1(\ks1.key_reg[79] ),
    .S(_03979_),
    .X(_04036_));
 sky130_fd_sc_hd__mux2_1 _16077_ (.A0(net143),
    .A1(\ks1.key_reg[111] ),
    .S(_03905_),
    .X(_04037_));
 sky130_fd_sc_hd__xor2_2 _16078_ (.A(_05244_),
    .B(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__xnor2_2 _16079_ (.A(_04036_),
    .B(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__xnor2_2 _16080_ (.A(_04035_),
    .B(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__xnor2_1 _16081_ (.A(_05005_),
    .B(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__mux2_1 _16082_ (.A0(\ks1.key_reg[15] ),
    .A1(_04041_),
    .S(_03958_),
    .X(_04042_));
 sky130_fd_sc_hd__clkbuf_1 _16083_ (.A(_04042_),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _16084_ (.A0(net144),
    .A1(\ks1.key_reg[112] ),
    .S(_03902_),
    .X(_04043_));
 sky130_fd_sc_hd__xor2_2 _16085_ (.A(\ks1.col[16] ),
    .B(_04043_),
    .X(_04044_));
 sky130_fd_sc_hd__mux2_1 _16086_ (.A0(net236),
    .A1(\ks1.key_reg[80] ),
    .S(_03907_),
    .X(_04045_));
 sky130_fd_sc_hd__xor2_2 _16087_ (.A(_04044_),
    .B(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__mux2_1 _16088_ (.A0(net200),
    .A1(\ks1.key_reg[48] ),
    .S(_03910_),
    .X(_04047_));
 sky130_fd_sc_hd__xor2_2 _16089_ (.A(_04046_),
    .B(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__or2_1 _16090_ (.A(_04915_),
    .B(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__a21oi_1 _16091_ (.A1(_04915_),
    .A2(_04048_),
    .B1(_03914_),
    .Y(_04050_));
 sky130_fd_sc_hd__a22o_1 _16092_ (.A1(net701),
    .A2(_03901_),
    .B1(_04049_),
    .B2(_04050_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_2 _16093_ (.A0(net145),
    .A1(\ks1.key_reg[113] ),
    .S(_03905_),
    .X(_04051_));
 sky130_fd_sc_hd__xor2_4 _16094_ (.A(\ks1.col[17] ),
    .B(_04051_),
    .X(_04052_));
 sky130_fd_sc_hd__mux2_2 _16095_ (.A0(net237),
    .A1(\ks1.key_reg[81] ),
    .S(_03906_),
    .X(_04053_));
 sky130_fd_sc_hd__xor2_4 _16096_ (.A(_04052_),
    .B(_04053_),
    .X(_04054_));
 sky130_fd_sc_hd__mux2_1 _16097_ (.A0(net201),
    .A1(\ks1.key_reg[49] ),
    .S(_03937_),
    .X(_04055_));
 sky130_fd_sc_hd__xor2_2 _16098_ (.A(_04054_),
    .B(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__xnor2_1 _16099_ (.A(_04754_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__mux2_1 _16100_ (.A0(\ks1.key_reg[17] ),
    .A1(_04057_),
    .S(_03958_),
    .X(_04058_));
 sky130_fd_sc_hd__clkbuf_1 _16101_ (.A(_04058_),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_2 _16102_ (.A0(net146),
    .A1(\ks1.key_reg[114] ),
    .S(_03905_),
    .X(_04059_));
 sky130_fd_sc_hd__xor2_4 _16103_ (.A(\ks1.col[18] ),
    .B(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__mux2_2 _16104_ (.A0(net238),
    .A1(\ks1.key_reg[82] ),
    .S(_03906_),
    .X(_04061_));
 sky130_fd_sc_hd__xor2_4 _16105_ (.A(_04060_),
    .B(_04061_),
    .X(_04062_));
 sky130_fd_sc_hd__mux2_1 _16106_ (.A0(net203),
    .A1(\ks1.key_reg[50] ),
    .S(_03937_),
    .X(_04063_));
 sky130_fd_sc_hd__xor2_2 _16107_ (.A(_04062_),
    .B(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__xnor2_1 _16108_ (.A(_05052_),
    .B(_04064_),
    .Y(_04065_));
 sky130_fd_sc_hd__mux2_1 _16109_ (.A0(\ks1.key_reg[18] ),
    .A1(_04065_),
    .S(_03958_),
    .X(_04066_));
 sky130_fd_sc_hd__clkbuf_1 _16110_ (.A(_04066_),
    .X(_01920_));
 sky130_fd_sc_hd__mux2_2 _16111_ (.A0(net147),
    .A1(\ks1.key_reg[115] ),
    .S(_03976_),
    .X(_04067_));
 sky130_fd_sc_hd__xor2_4 _16112_ (.A(\ks1.col[19] ),
    .B(_04067_),
    .X(_04068_));
 sky130_fd_sc_hd__mux2_2 _16113_ (.A0(net239),
    .A1(\ks1.key_reg[83] ),
    .S(_03906_),
    .X(_04069_));
 sky130_fd_sc_hd__xor2_4 _16114_ (.A(_04068_),
    .B(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__mux2_1 _16115_ (.A0(net204),
    .A1(\ks1.key_reg[51] ),
    .S(_03937_),
    .X(_04071_));
 sky130_fd_sc_hd__xor2_2 _16116_ (.A(_04070_),
    .B(_04071_),
    .X(_04072_));
 sky130_fd_sc_hd__xnor2_1 _16117_ (.A(_04796_),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__mux2_1 _16118_ (.A0(\ks1.key_reg[19] ),
    .A1(_04073_),
    .S(_03958_),
    .X(_04074_));
 sky130_fd_sc_hd__clkbuf_1 _16119_ (.A(_04074_),
    .X(_01921_));
 sky130_fd_sc_hd__mux2_2 _16120_ (.A0(net148),
    .A1(\ks1.key_reg[116] ),
    .S(_03976_),
    .X(_04075_));
 sky130_fd_sc_hd__xor2_4 _16121_ (.A(\ks1.col[20] ),
    .B(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__mux2_2 _16122_ (.A0(net240),
    .A1(\ks1.key_reg[84] ),
    .S(_03906_),
    .X(_04077_));
 sky130_fd_sc_hd__xor2_4 _16123_ (.A(_04076_),
    .B(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__mux2_1 _16124_ (.A0(net205),
    .A1(\ks1.key_reg[52] ),
    .S(_03937_),
    .X(_04079_));
 sky130_fd_sc_hd__xor2_2 _16125_ (.A(_04078_),
    .B(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__xnor2_1 _16126_ (.A(_04744_),
    .B(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__mux2_1 _16127_ (.A0(\ks1.key_reg[20] ),
    .A1(_04081_),
    .S(_03958_),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _16128_ (.A(_04082_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _16129_ (.A0(net149),
    .A1(\ks1.key_reg[117] ),
    .S(_03902_),
    .X(_04083_));
 sky130_fd_sc_hd__xor2_2 _16130_ (.A(\ks1.col[21] ),
    .B(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__mux2_1 _16131_ (.A0(net241),
    .A1(\ks1.key_reg[85] ),
    .S(_03918_),
    .X(_04085_));
 sky130_fd_sc_hd__xor2_2 _16132_ (.A(_04084_),
    .B(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__mux2_1 _16133_ (.A0(net206),
    .A1(\ks1.key_reg[53] ),
    .S(_03910_),
    .X(_04087_));
 sky130_fd_sc_hd__xor2_2 _16134_ (.A(_04086_),
    .B(_04087_),
    .X(_04088_));
 sky130_fd_sc_hd__or2_1 _16135_ (.A(_04957_),
    .B(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__a21oi_1 _16136_ (.A1(_04957_),
    .A2(_04088_),
    .B1(_03914_),
    .Y(_04090_));
 sky130_fd_sc_hd__a22o_1 _16137_ (.A1(net698),
    .A2(_03901_),
    .B1(_04089_),
    .B2(_04090_),
    .X(_01923_));
 sky130_fd_sc_hd__mux2_1 _16138_ (.A0(net150),
    .A1(\ks1.key_reg[118] ),
    .S(_03976_),
    .X(_04091_));
 sky130_fd_sc_hd__xor2_2 _16139_ (.A(\ks1.col[22] ),
    .B(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__mux2_1 _16140_ (.A0(net242),
    .A1(\ks1.key_reg[86] ),
    .S(_03906_),
    .X(_04093_));
 sky130_fd_sc_hd__xor2_2 _16141_ (.A(_04092_),
    .B(_04093_),
    .X(_04094_));
 sky130_fd_sc_hd__mux2_1 _16142_ (.A0(net207),
    .A1(\ks1.key_reg[54] ),
    .S(_03982_),
    .X(_04095_));
 sky130_fd_sc_hd__xor2_1 _16143_ (.A(_04094_),
    .B(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__xnor2_1 _16144_ (.A(_04868_),
    .B(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__mux2_1 _16145_ (.A0(\ks1.key_reg[22] ),
    .A1(_04097_),
    .S(_03958_),
    .X(_04098_));
 sky130_fd_sc_hd__clkbuf_1 _16146_ (.A(_04098_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _16147_ (.A0(net151),
    .A1(\ks1.key_reg[119] ),
    .S(_03976_),
    .X(_04099_));
 sky130_fd_sc_hd__xor2_2 _16148_ (.A(\ks1.col[23] ),
    .B(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__mux2_1 _16149_ (.A0(net243),
    .A1(\ks1.key_reg[87] ),
    .S(_03906_),
    .X(_04101_));
 sky130_fd_sc_hd__xor2_2 _16150_ (.A(_04100_),
    .B(_04101_),
    .X(_04102_));
 sky130_fd_sc_hd__mux2_1 _16151_ (.A0(net208),
    .A1(\ks1.key_reg[55] ),
    .S(_03982_),
    .X(_04103_));
 sky130_fd_sc_hd__xor2_1 _16152_ (.A(_04102_),
    .B(_04103_),
    .X(_04104_));
 sky130_fd_sc_hd__xnor2_1 _16153_ (.A(_05000_),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__buf_4 _16154_ (.A(_03957_),
    .X(_04106_));
 sky130_fd_sc_hd__mux2_1 _16155_ (.A0(\ks1.key_reg[23] ),
    .A1(_04105_),
    .S(_04106_),
    .X(_04107_));
 sky130_fd_sc_hd__clkbuf_1 _16156_ (.A(_04107_),
    .X(_01925_));
 sky130_fd_sc_hd__inv_2 _16157_ (.A(\addroundkey_round[1] ),
    .Y(_04108_));
 sky130_fd_sc_hd__or2b_1 _16158_ (.A(_04727_),
    .B_N(_04638_),
    .X(_04109_));
 sky130_fd_sc_hd__nor2_1 _16159_ (.A(_04644_),
    .B(_05539_),
    .Y(_04110_));
 sky130_fd_sc_hd__a211o_2 _16160_ (.A1(_04108_),
    .A2(_04109_),
    .B1(_04110_),
    .C1(_04723_),
    .X(_04111_));
 sky130_fd_sc_hd__a31oi_4 _16161_ (.A1(\addroundkey_round[2] ),
    .A2(_04642_),
    .A3(_04644_),
    .B1(_05542_),
    .Y(_04112_));
 sky130_fd_sc_hd__a211o_2 _16162_ (.A1(\addroundkey_round[0] ),
    .A2(_04109_),
    .B1(_05538_),
    .C1(_04723_),
    .X(_04113_));
 sky130_fd_sc_hd__and3_1 _16163_ (.A(_04111_),
    .B(_04112_),
    .C(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__xnor2_2 _16164_ (.A(\ks1.col[24] ),
    .B(_04114_),
    .Y(_04115_));
 sky130_fd_sc_hd__mux2_1 _16165_ (.A0(net153),
    .A1(\ks1.key_reg[120] ),
    .S(_03976_),
    .X(_04116_));
 sky130_fd_sc_hd__xor2_2 _16166_ (.A(_04115_),
    .B(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__mux2_1 _16167_ (.A0(net244),
    .A1(\ks1.key_reg[88] ),
    .S(_03906_),
    .X(_04118_));
 sky130_fd_sc_hd__xnor2_2 _16168_ (.A(_04117_),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__mux2_1 _16169_ (.A0(net209),
    .A1(\ks1.key_reg[56] ),
    .S(_03982_),
    .X(_04120_));
 sky130_fd_sc_hd__xor2_1 _16170_ (.A(_04119_),
    .B(_04120_),
    .X(_04121_));
 sky130_fd_sc_hd__xnor2_1 _16171_ (.A(_04918_),
    .B(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__mux2_1 _16172_ (.A0(\ks1.key_reg[24] ),
    .A1(_04122_),
    .S(_04106_),
    .X(_04123_));
 sky130_fd_sc_hd__clkbuf_1 _16173_ (.A(_04123_),
    .X(_01926_));
 sky130_fd_sc_hd__xnor2_1 _16174_ (.A(_04111_),
    .B(_04113_),
    .Y(_04124_));
 sky130_fd_sc_hd__a31oi_4 _16175_ (.A1(\addroundkey_round[3] ),
    .A2(_04642_),
    .A3(_04644_),
    .B1(_05544_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _16176_ (.A(_04113_),
    .B(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__and3_1 _16177_ (.A(_04112_),
    .B(_04124_),
    .C(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__xor2_4 _16178_ (.A(\ks1.col[25] ),
    .B(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__mux2_2 _16179_ (.A0(net154),
    .A1(\ks1.key_reg[121] ),
    .S(_03902_),
    .X(_04129_));
 sky130_fd_sc_hd__xnor2_4 _16180_ (.A(_04128_),
    .B(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__mux2_2 _16181_ (.A0(net245),
    .A1(\ks1.key_reg[89] ),
    .S(_03918_),
    .X(_04131_));
 sky130_fd_sc_hd__xor2_4 _16182_ (.A(_04130_),
    .B(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__mux2_1 _16183_ (.A0(net210),
    .A1(\ks1.key_reg[57] ),
    .S(_03937_),
    .X(_04133_));
 sky130_fd_sc_hd__xor2_2 _16184_ (.A(_04132_),
    .B(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__xnor2_1 _16185_ (.A(_04761_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__buf_4 _16186_ (.A(_04371_),
    .X(_04136_));
 sky130_fd_sc_hd__nand2_1 _16187_ (.A(net712),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__o21ai_1 _16188_ (.A1(_03901_),
    .A2(_04135_),
    .B1(_04137_),
    .Y(_01927_));
 sky130_fd_sc_hd__inv_2 _16189_ (.A(_04112_),
    .Y(_04138_));
 sky130_fd_sc_hd__or2_1 _16190_ (.A(_04113_),
    .B(_04125_),
    .X(_04139_));
 sky130_fd_sc_hd__and2_1 _16191_ (.A(_04126_),
    .B(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__or3_2 _16192_ (.A(_04111_),
    .B(_04138_),
    .C(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__xnor2_4 _16193_ (.A(\ks1.col[26] ),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__mux2_2 _16194_ (.A0(net155),
    .A1(\ks1.key_reg[122] ),
    .S(_03902_),
    .X(_04143_));
 sky130_fd_sc_hd__xnor2_4 _16195_ (.A(_04142_),
    .B(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__mux2_1 _16196_ (.A0(net247),
    .A1(\ks1.key_reg[90] ),
    .S(_03918_),
    .X(_04145_));
 sky130_fd_sc_hd__xor2_2 _16197_ (.A(_04144_),
    .B(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__mux2_1 _16198_ (.A0(net211),
    .A1(\ks1.key_reg[58] ),
    .S(_03937_),
    .X(_04147_));
 sky130_fd_sc_hd__xor2_2 _16199_ (.A(_04146_),
    .B(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__xnor2_1 _16200_ (.A(_05046_),
    .B(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__nand2_1 _16201_ (.A(net714),
    .B(_04136_),
    .Y(_04150_));
 sky130_fd_sc_hd__o21ai_1 _16202_ (.A1(_03901_),
    .A2(_04149_),
    .B1(_04150_),
    .Y(_01928_));
 sky130_fd_sc_hd__xor2_1 _16203_ (.A(_04112_),
    .B(_04125_),
    .X(_04151_));
 sky130_fd_sc_hd__and3_2 _16204_ (.A(_04111_),
    .B(_04140_),
    .C(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__xnor2_4 _16205_ (.A(\ks1.col[27] ),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__mux2_2 _16206_ (.A0(net156),
    .A1(\ks1.key_reg[123] ),
    .S(_04742_),
    .X(_04154_));
 sky130_fd_sc_hd__xor2_4 _16207_ (.A(_04153_),
    .B(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__mux2_2 _16208_ (.A0(net248),
    .A1(\ks1.key_reg[91] ),
    .S(_03979_),
    .X(_04156_));
 sky130_fd_sc_hd__xnor2_4 _16209_ (.A(_04155_),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__mux2_1 _16210_ (.A0(net212),
    .A1(\ks1.key_reg[59] ),
    .S(_03907_),
    .X(_04158_));
 sky130_fd_sc_hd__xnor2_2 _16211_ (.A(_04157_),
    .B(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__xnor2_1 _16212_ (.A(_04831_),
    .B(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__mux2_1 _16213_ (.A0(net795),
    .A1(_04160_),
    .S(_04106_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _16214_ (.A(_04161_),
    .X(_01929_));
 sky130_fd_sc_hd__o211a_1 _16215_ (.A1(_04112_),
    .A2(_04113_),
    .B1(_04124_),
    .C1(_04151_),
    .X(_04162_));
 sky130_fd_sc_hd__xor2_4 _16216_ (.A(\ks1.col[28] ),
    .B(_04162_),
    .X(_04163_));
 sky130_fd_sc_hd__mux2_2 _16217_ (.A0(net157),
    .A1(\ks1.key_reg[124] ),
    .S(_03976_),
    .X(_04164_));
 sky130_fd_sc_hd__xnor2_4 _16218_ (.A(_04163_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__mux2_1 _16219_ (.A0(net249),
    .A1(\ks1.key_reg[92] ),
    .S(_03979_),
    .X(_04166_));
 sky130_fd_sc_hd__xor2_2 _16220_ (.A(_04165_),
    .B(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__mux2_1 _16221_ (.A0(net214),
    .A1(\ks1.key_reg[60] ),
    .S(_03982_),
    .X(_04168_));
 sky130_fd_sc_hd__xor2_2 _16222_ (.A(_04167_),
    .B(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__xnor2_1 _16223_ (.A(_04748_),
    .B(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__mux2_1 _16224_ (.A0(\ks1.key_reg[28] ),
    .A1(_04170_),
    .S(_04106_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _16225_ (.A(_04171_),
    .X(_01930_));
 sky130_fd_sc_hd__or3b_2 _16226_ (.A(_04111_),
    .B(_04113_),
    .C_N(_04151_),
    .X(_04172_));
 sky130_fd_sc_hd__xnor2_4 _16227_ (.A(\ks1.col[29] ),
    .B(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__mux2_2 _16228_ (.A0(net158),
    .A1(\ks1.key_reg[125] ),
    .S(_03976_),
    .X(_04174_));
 sky130_fd_sc_hd__xnor2_4 _16229_ (.A(_04173_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__mux2_1 _16230_ (.A0(net250),
    .A1(\ks1.key_reg[93] ),
    .S(_03979_),
    .X(_04176_));
 sky130_fd_sc_hd__xor2_2 _16231_ (.A(_04175_),
    .B(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__mux2_1 _16232_ (.A0(net215),
    .A1(\ks1.key_reg[61] ),
    .S(_03982_),
    .X(_04178_));
 sky130_fd_sc_hd__xor2_2 _16233_ (.A(_04177_),
    .B(_04178_),
    .X(_04179_));
 sky130_fd_sc_hd__xnor2_1 _16234_ (.A(_04963_),
    .B(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__mux2_1 _16235_ (.A0(\ks1.key_reg[29] ),
    .A1(_04180_),
    .S(_04106_),
    .X(_04181_));
 sky130_fd_sc_hd__clkbuf_1 _16236_ (.A(_04181_),
    .X(_01931_));
 sky130_fd_sc_hd__or3_2 _16237_ (.A(_04111_),
    .B(_04112_),
    .C(_04126_),
    .X(_04182_));
 sky130_fd_sc_hd__xnor2_4 _16238_ (.A(\ks1.col[30] ),
    .B(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__mux2_2 _16239_ (.A0(net159),
    .A1(\ks1.key_reg[126] ),
    .S(_03976_),
    .X(_04184_));
 sky130_fd_sc_hd__xnor2_4 _16240_ (.A(_04183_),
    .B(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__mux2_2 _16241_ (.A0(net251),
    .A1(\ks1.key_reg[94] ),
    .S(_03918_),
    .X(_04186_));
 sky130_fd_sc_hd__xor2_4 _16242_ (.A(_04185_),
    .B(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__mux2_1 _16243_ (.A0(net216),
    .A1(\ks1.key_reg[62] ),
    .S(_03937_),
    .X(_04188_));
 sky130_fd_sc_hd__xor2_2 _16244_ (.A(_04187_),
    .B(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__nor2_1 _16245_ (.A(_04869_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__a21o_1 _16246_ (.A1(_04869_),
    .A2(_04189_),
    .B1(_04371_),
    .X(_04191_));
 sky130_fd_sc_hd__o22a_1 _16247_ (.A1(net689),
    .A2(\ks1.next_ready_o ),
    .B1(_04190_),
    .B2(_04191_),
    .X(_01932_));
 sky130_fd_sc_hd__or4b_4 _16248_ (.A(_04138_),
    .B(_04113_),
    .C(_04125_),
    .D_N(_04111_),
    .X(_04192_));
 sky130_fd_sc_hd__xnor2_4 _16249_ (.A(\ks1.col[31] ),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__mux2_2 _16250_ (.A0(net160),
    .A1(\ks1.key_reg[127] ),
    .S(_04742_),
    .X(_04194_));
 sky130_fd_sc_hd__xnor2_4 _16251_ (.A(_04193_),
    .B(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__mux2_2 _16252_ (.A0(net252),
    .A1(\ks1.key_reg[95] ),
    .S(_03979_),
    .X(_04196_));
 sky130_fd_sc_hd__xor2_4 _16253_ (.A(_04195_),
    .B(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__mux2_1 _16254_ (.A0(net217),
    .A1(\ks1.key_reg[63] ),
    .S(_03982_),
    .X(_04198_));
 sky130_fd_sc_hd__xor2_2 _16255_ (.A(_04197_),
    .B(_04198_),
    .X(_04199_));
 sky130_fd_sc_hd__xnor2_1 _16256_ (.A(_05002_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__mux2_1 _16257_ (.A0(\ks1.key_reg[31] ),
    .A1(_04200_),
    .S(_04106_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _16258_ (.A(_04201_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _16259_ (.A0(net824),
    .A1(_03912_),
    .S(_04106_),
    .X(_04202_));
 sky130_fd_sc_hd__clkbuf_1 _16260_ (.A(_04202_),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_1 _16261_ (.A0(net813),
    .A1(_03922_),
    .S(_04106_),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_1 _16262_ (.A(_04203_),
    .X(_01935_));
 sky130_fd_sc_hd__mux2_1 _16263_ (.A0(net820),
    .A1(_03930_),
    .S(_04106_),
    .X(_04204_));
 sky130_fd_sc_hd__clkbuf_1 _16264_ (.A(_04204_),
    .X(_01936_));
 sky130_fd_sc_hd__mux2_1 _16265_ (.A0(\ks1.key_reg[35] ),
    .A1(_03939_),
    .S(_04106_),
    .X(_04205_));
 sky130_fd_sc_hd__clkbuf_1 _16266_ (.A(_04205_),
    .X(_01937_));
 sky130_fd_sc_hd__buf_4 _16267_ (.A(_03957_),
    .X(_04206_));
 sky130_fd_sc_hd__mux2_1 _16268_ (.A0(net825),
    .A1(_03947_),
    .S(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__clkbuf_1 _16269_ (.A(_04207_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_1 _16270_ (.A0(\ks1.key_reg[37] ),
    .A1(_03955_),
    .S(_04206_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_1 _16271_ (.A(_04208_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _16272_ (.A0(\ks1.key_reg[38] ),
    .A1(_03965_),
    .S(_04206_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _16273_ (.A(_04209_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _16274_ (.A0(\ks1.key_reg[39] ),
    .A1(_03973_),
    .S(_04206_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _16275_ (.A(_04210_),
    .X(_01941_));
 sky130_fd_sc_hd__nand2_1 _16276_ (.A(net677),
    .B(_04136_),
    .Y(_04211_));
 sky130_fd_sc_hd__o21ai_1 _16277_ (.A1(_03901_),
    .A2(_03984_),
    .B1(_04211_),
    .Y(_01942_));
 sky130_fd_sc_hd__nor2_1 _16278_ (.A(net683),
    .B(_04373_),
    .Y(_04212_));
 sky130_fd_sc_hd__a21oi_1 _16279_ (.A1(\ks1.next_ready_o ),
    .A2(_03992_),
    .B1(_04212_),
    .Y(_01943_));
 sky130_fd_sc_hd__mux2_1 _16280_ (.A0(\ks1.key_reg[42] ),
    .A1(_04000_),
    .S(_04206_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _16281_ (.A(_04213_),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _16282_ (.A0(\ks1.key_reg[43] ),
    .A1(_04008_),
    .S(_04206_),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_1 _16283_ (.A(_04214_),
    .X(_01945_));
 sky130_fd_sc_hd__buf_4 _16284_ (.A(_04371_),
    .X(_04215_));
 sky130_fd_sc_hd__nand2_1 _16285_ (.A(net679),
    .B(_04136_),
    .Y(_04216_));
 sky130_fd_sc_hd__o21ai_1 _16286_ (.A1(_04215_),
    .A2(_04016_),
    .B1(_04216_),
    .Y(_01946_));
 sky130_fd_sc_hd__inv_2 _16287_ (.A(_04024_),
    .Y(_04217_));
 sky130_fd_sc_hd__mux2_1 _16288_ (.A0(net818),
    .A1(_04217_),
    .S(_04206_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _16289_ (.A(_04218_),
    .X(_01947_));
 sky130_fd_sc_hd__mux2_1 _16290_ (.A0(net841),
    .A1(_04032_),
    .S(_04206_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _16291_ (.A(_04219_),
    .X(_01948_));
 sky130_fd_sc_hd__mux2_1 _16292_ (.A0(net830),
    .A1(_04040_),
    .S(_04206_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _16293_ (.A(_04220_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _16294_ (.A0(net811),
    .A1(_04048_),
    .S(_04206_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _16295_ (.A(_04221_),
    .X(_01950_));
 sky130_fd_sc_hd__buf_4 _16296_ (.A(_03957_),
    .X(_04222_));
 sky130_fd_sc_hd__mux2_1 _16297_ (.A0(net834),
    .A1(_04056_),
    .S(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__clkbuf_1 _16298_ (.A(_04223_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _16299_ (.A0(net833),
    .A1(_04064_),
    .S(_04222_),
    .X(_04224_));
 sky130_fd_sc_hd__clkbuf_1 _16300_ (.A(_04224_),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_1 _16301_ (.A0(net816),
    .A1(_04072_),
    .S(_04222_),
    .X(_04225_));
 sky130_fd_sc_hd__clkbuf_1 _16302_ (.A(_04225_),
    .X(_01953_));
 sky130_fd_sc_hd__mux2_1 _16303_ (.A0(\ks1.key_reg[52] ),
    .A1(_04080_),
    .S(_04222_),
    .X(_04226_));
 sky130_fd_sc_hd__clkbuf_1 _16304_ (.A(_04226_),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _16305_ (.A0(net810),
    .A1(_04088_),
    .S(_04222_),
    .X(_04227_));
 sky130_fd_sc_hd__clkbuf_1 _16306_ (.A(_04227_),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _16307_ (.A0(net821),
    .A1(_04096_),
    .S(_04222_),
    .X(_04228_));
 sky130_fd_sc_hd__clkbuf_1 _16308_ (.A(_04228_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _16309_ (.A0(net809),
    .A1(_04104_),
    .S(_04222_),
    .X(_04229_));
 sky130_fd_sc_hd__clkbuf_1 _16310_ (.A(_04229_),
    .X(_01957_));
 sky130_fd_sc_hd__mux2_1 _16311_ (.A0(net807),
    .A1(_04121_),
    .S(_04222_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _16312_ (.A(_04230_),
    .X(_01958_));
 sky130_fd_sc_hd__nand2_1 _16313_ (.A(net673),
    .B(_04136_),
    .Y(_04231_));
 sky130_fd_sc_hd__o21ai_1 _16314_ (.A1(_04215_),
    .A2(_04134_),
    .B1(_04231_),
    .Y(_01959_));
 sky130_fd_sc_hd__nand2_1 _16315_ (.A(net680),
    .B(_04136_),
    .Y(_04232_));
 sky130_fd_sc_hd__o21ai_1 _16316_ (.A1(_04215_),
    .A2(_04148_),
    .B1(_04232_),
    .Y(_01960_));
 sky130_fd_sc_hd__nor2_1 _16317_ (.A(net690),
    .B(_04373_),
    .Y(_04233_));
 sky130_fd_sc_hd__a21oi_1 _16318_ (.A1(\ks1.next_ready_o ),
    .A2(_04159_),
    .B1(_04233_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand2_1 _16319_ (.A(net676),
    .B(_04136_),
    .Y(_04234_));
 sky130_fd_sc_hd__o21ai_1 _16320_ (.A1(_04215_),
    .A2(_04169_),
    .B1(_04234_),
    .Y(_01962_));
 sky130_fd_sc_hd__nand2_1 _16321_ (.A(net672),
    .B(_04136_),
    .Y(_04235_));
 sky130_fd_sc_hd__o21ai_1 _16322_ (.A1(_04215_),
    .A2(_04179_),
    .B1(_04235_),
    .Y(_01963_));
 sky130_fd_sc_hd__inv_2 _16323_ (.A(_04189_),
    .Y(_04236_));
 sky130_fd_sc_hd__mux2_1 _16324_ (.A0(\ks1.key_reg[62] ),
    .A1(_04236_),
    .S(_04222_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_1 _16325_ (.A(_04237_),
    .X(_01964_));
 sky130_fd_sc_hd__nand2_1 _16326_ (.A(net674),
    .B(_04136_),
    .Y(_04238_));
 sky130_fd_sc_hd__o21ai_1 _16327_ (.A1(_04215_),
    .A2(_04199_),
    .B1(_04238_),
    .Y(_01965_));
 sky130_fd_sc_hd__mux2_1 _16328_ (.A0(net845),
    .A1(_03909_),
    .S(_04222_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _16329_ (.A(_04239_),
    .X(_01966_));
 sky130_fd_sc_hd__buf_4 _16330_ (.A(_04372_),
    .X(_04240_));
 sky130_fd_sc_hd__mux2_1 _16331_ (.A0(net838),
    .A1(_03920_),
    .S(_04240_),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_1 _16332_ (.A(_04241_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _16333_ (.A0(\ks1.key_reg[66] ),
    .A1(_03928_),
    .S(_04240_),
    .X(_04242_));
 sky130_fd_sc_hd__clkbuf_1 _16334_ (.A(_04242_),
    .X(_01968_));
 sky130_fd_sc_hd__mux2_1 _16335_ (.A0(net836),
    .A1(_03936_),
    .S(_04240_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _16336_ (.A(_04243_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _16337_ (.A0(net847),
    .A1(_03945_),
    .S(_04240_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _16338_ (.A(_04244_),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_1 _16339_ (.A0(net823),
    .A1(_03953_),
    .S(_04240_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _16340_ (.A(_04245_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_1 _16341_ (.A0(net802),
    .A1(_03963_),
    .S(_04240_),
    .X(_04246_));
 sky130_fd_sc_hd__clkbuf_1 _16342_ (.A(_04246_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _16343_ (.A0(net829),
    .A1(_03971_),
    .S(_04240_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_1 _16344_ (.A(_04247_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _16345_ (.A0(\ks1.key_reg[72] ),
    .A1(_03981_),
    .S(_04240_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_1 _16346_ (.A(_04248_),
    .X(_01974_));
 sky130_fd_sc_hd__mux2_1 _16347_ (.A0(\ks1.key_reg[73] ),
    .A1(_03990_),
    .S(_04240_),
    .X(_04249_));
 sky130_fd_sc_hd__clkbuf_1 _16348_ (.A(_04249_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _16349_ (.A0(net832),
    .A1(_03999_),
    .S(_04240_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _16350_ (.A(_04250_),
    .X(_01976_));
 sky130_fd_sc_hd__nor2_1 _16351_ (.A(net692),
    .B(_04373_),
    .Y(_04251_));
 sky130_fd_sc_hd__a21oi_1 _16352_ (.A1(\ks1.next_ready_o ),
    .A2(_04007_),
    .B1(_04251_),
    .Y(_01977_));
 sky130_fd_sc_hd__buf_4 _16353_ (.A(_04372_),
    .X(_04252_));
 sky130_fd_sc_hd__mux2_1 _16354_ (.A0(net796),
    .A1(_04014_),
    .S(_04252_),
    .X(_04253_));
 sky130_fd_sc_hd__clkbuf_1 _16355_ (.A(_04253_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _16356_ (.A0(\ks1.key_reg[77] ),
    .A1(_04023_),
    .S(_04252_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _16357_ (.A(_04254_),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_1 _16358_ (.A0(net817),
    .A1(_04030_),
    .S(_04252_),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_1 _16359_ (.A(_04255_),
    .X(_01980_));
 sky130_fd_sc_hd__nor2_1 _16360_ (.A(net685),
    .B(_04373_),
    .Y(_04256_));
 sky130_fd_sc_hd__a21oi_1 _16361_ (.A1(\ks1.next_ready_o ),
    .A2(_04039_),
    .B1(_04256_),
    .Y(_01981_));
 sky130_fd_sc_hd__mux2_1 _16362_ (.A0(net837),
    .A1(_04046_),
    .S(_04252_),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_1 _16363_ (.A(_04257_),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _16364_ (.A0(\ks1.key_reg[81] ),
    .A1(_04054_),
    .S(_04252_),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_1 _16365_ (.A(_04258_),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_1 _16366_ (.A0(net843),
    .A1(_04062_),
    .S(_04252_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _16367_ (.A(_04259_),
    .X(_01984_));
 sky130_fd_sc_hd__mux2_1 _16368_ (.A0(net808),
    .A1(_04070_),
    .S(_04252_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _16369_ (.A(_04260_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _16370_ (.A0(net803),
    .A1(_04078_),
    .S(_04252_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _16371_ (.A(_04261_),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_1 _16372_ (.A0(net800),
    .A1(_04086_),
    .S(_04252_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _16373_ (.A(_04262_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _16374_ (.A0(net805),
    .A1(_04094_),
    .S(_04252_),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _16375_ (.A(_04263_),
    .X(_01988_));
 sky130_fd_sc_hd__buf_4 _16376_ (.A(_04372_),
    .X(_04264_));
 sky130_fd_sc_hd__mux2_1 _16377_ (.A0(net831),
    .A1(_04102_),
    .S(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _16378_ (.A(_04265_),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_1 _16379_ (.A0(net822),
    .A1(_04119_),
    .S(_04264_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_1 _16380_ (.A(_04266_),
    .X(_01990_));
 sky130_fd_sc_hd__inv_2 _16381_ (.A(_04132_),
    .Y(_04267_));
 sky130_fd_sc_hd__mux2_1 _16382_ (.A0(net848),
    .A1(_04267_),
    .S(_04264_),
    .X(_04268_));
 sky130_fd_sc_hd__clkbuf_1 _16383_ (.A(_04268_),
    .X(_01991_));
 sky130_fd_sc_hd__inv_2 _16384_ (.A(_04146_),
    .Y(_04269_));
 sky130_fd_sc_hd__mux2_1 _16385_ (.A0(\ks1.key_reg[90] ),
    .A1(_04269_),
    .S(_04264_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _16386_ (.A(_04270_),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_1 _16387_ (.A0(net844),
    .A1(_04157_),
    .S(_04264_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _16388_ (.A(_04271_),
    .X(_01993_));
 sky130_fd_sc_hd__inv_2 _16389_ (.A(_04167_),
    .Y(_04272_));
 sky130_fd_sc_hd__mux2_1 _16390_ (.A0(\ks1.key_reg[92] ),
    .A1(_04272_),
    .S(_04264_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_1 _16391_ (.A(_04273_),
    .X(_01994_));
 sky130_fd_sc_hd__inv_2 _16392_ (.A(_04177_),
    .Y(_04274_));
 sky130_fd_sc_hd__mux2_1 _16393_ (.A0(\ks1.key_reg[93] ),
    .A1(_04274_),
    .S(_04264_),
    .X(_04275_));
 sky130_fd_sc_hd__clkbuf_1 _16394_ (.A(_04275_),
    .X(_01995_));
 sky130_fd_sc_hd__inv_2 _16395_ (.A(_04187_),
    .Y(_04276_));
 sky130_fd_sc_hd__mux2_1 _16396_ (.A0(\ks1.key_reg[94] ),
    .A1(_04276_),
    .S(_04264_),
    .X(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _16397_ (.A(_04277_),
    .X(_01996_));
 sky130_fd_sc_hd__inv_2 _16398_ (.A(_04197_),
    .Y(_04278_));
 sky130_fd_sc_hd__mux2_1 _16399_ (.A0(\ks1.key_reg[95] ),
    .A1(_04278_),
    .S(_04264_),
    .X(_04279_));
 sky130_fd_sc_hd__clkbuf_1 _16400_ (.A(_04279_),
    .X(_01997_));
 sky130_fd_sc_hd__mux2_1 _16401_ (.A0(\ks1.key_reg[96] ),
    .A1(_03904_),
    .S(_04264_),
    .X(_04280_));
 sky130_fd_sc_hd__clkbuf_1 _16402_ (.A(_04280_),
    .X(_01998_));
 sky130_fd_sc_hd__buf_4 _16403_ (.A(_04372_),
    .X(_04281_));
 sky130_fd_sc_hd__mux2_1 _16404_ (.A0(net827),
    .A1(_03917_),
    .S(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _16405_ (.A(_04282_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _16406_ (.A0(net828),
    .A1(_03926_),
    .S(_04281_),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _16407_ (.A(_04283_),
    .X(_02000_));
 sky130_fd_sc_hd__mux2_1 _16408_ (.A0(net799),
    .A1(_03934_),
    .S(_04281_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_1 _16409_ (.A(_04284_),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_1 _16410_ (.A0(\ks1.key_reg[100] ),
    .A1(_03943_),
    .S(_04281_),
    .X(_04285_));
 sky130_fd_sc_hd__clkbuf_1 _16411_ (.A(_04285_),
    .X(_02002_));
 sky130_fd_sc_hd__mux2_1 _16412_ (.A0(\ks1.key_reg[101] ),
    .A1(_03951_),
    .S(_04281_),
    .X(_04286_));
 sky130_fd_sc_hd__clkbuf_1 _16413_ (.A(_04286_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _16414_ (.A0(net804),
    .A1(_03961_),
    .S(_04281_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_1 _16415_ (.A(_04287_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _16416_ (.A0(net826),
    .A1(_03969_),
    .S(_04281_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_1 _16417_ (.A(_04288_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _16418_ (.A0(net812),
    .A1(_03978_),
    .S(_04281_),
    .X(_04289_));
 sky130_fd_sc_hd__clkbuf_1 _16419_ (.A(_04289_),
    .X(_02006_));
 sky130_fd_sc_hd__nand2_1 _16420_ (.A(net721),
    .B(_04136_),
    .Y(_04290_));
 sky130_fd_sc_hd__o21ai_1 _16421_ (.A1(_04215_),
    .A2(_03989_),
    .B1(_04290_),
    .Y(_02007_));
 sky130_fd_sc_hd__mux2_1 _16422_ (.A0(\ks1.key_reg[106] ),
    .A1(_03998_),
    .S(_04281_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _16423_ (.A(_04291_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _16424_ (.A0(net797),
    .A1(_04006_),
    .S(_04281_),
    .X(_04292_));
 sky130_fd_sc_hd__clkbuf_1 _16425_ (.A(_04292_),
    .X(_02009_));
 sky130_fd_sc_hd__nand2_1 _16426_ (.A(net678),
    .B(_03914_),
    .Y(_04293_));
 sky130_fd_sc_hd__o21ai_1 _16427_ (.A1(_04215_),
    .A2(_04012_),
    .B1(_04293_),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _16428_ (.A(net686),
    .B(_03914_),
    .Y(_04294_));
 sky130_fd_sc_hd__o21ai_1 _16429_ (.A1(_04215_),
    .A2(_04022_),
    .B1(_04294_),
    .Y(_02011_));
 sky130_fd_sc_hd__buf_4 _16430_ (.A(_04372_),
    .X(_04295_));
 sky130_fd_sc_hd__mux2_1 _16431_ (.A0(\ks1.key_reg[110] ),
    .A1(_04028_),
    .S(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _16432_ (.A(_04296_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _16433_ (.A0(\ks1.key_reg[111] ),
    .A1(_04038_),
    .S(_04295_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_1 _16434_ (.A(_04297_),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _16435_ (.A0(\ks1.key_reg[112] ),
    .A1(_04044_),
    .S(_04295_),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_1 _16436_ (.A(_04298_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _16437_ (.A0(net814),
    .A1(_04052_),
    .S(_04295_),
    .X(_04299_));
 sky130_fd_sc_hd__clkbuf_1 _16438_ (.A(_04299_),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _16439_ (.A0(net794),
    .A1(_04060_),
    .S(_04295_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _16440_ (.A(_04300_),
    .X(_02016_));
 sky130_fd_sc_hd__mux2_1 _16441_ (.A0(net793),
    .A1(_04068_),
    .S(_04295_),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _16442_ (.A(_04301_),
    .X(_02017_));
 sky130_fd_sc_hd__mux2_1 _16443_ (.A0(net842),
    .A1(_04076_),
    .S(_04295_),
    .X(_04302_));
 sky130_fd_sc_hd__clkbuf_1 _16444_ (.A(_04302_),
    .X(_02018_));
 sky130_fd_sc_hd__mux2_1 _16445_ (.A0(net846),
    .A1(_04084_),
    .S(_04295_),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_1 _16446_ (.A(_04303_),
    .X(_02019_));
 sky130_fd_sc_hd__mux2_1 _16447_ (.A0(net835),
    .A1(_04092_),
    .S(_04295_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _16448_ (.A(_04304_),
    .X(_02020_));
 sky130_fd_sc_hd__mux2_1 _16449_ (.A0(net801),
    .A1(_04100_),
    .S(_04295_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _16450_ (.A(_04305_),
    .X(_02021_));
 sky130_fd_sc_hd__nand2_1 _16451_ (.A(net681),
    .B(_03914_),
    .Y(_04306_));
 sky130_fd_sc_hd__o21ai_1 _16452_ (.A1(_04215_),
    .A2(_04117_),
    .B1(_04306_),
    .Y(_02022_));
 sky130_fd_sc_hd__inv_2 _16453_ (.A(_04130_),
    .Y(_04307_));
 sky130_fd_sc_hd__mux2_1 _16454_ (.A0(\ks1.key_reg[121] ),
    .A1(_04307_),
    .S(_03957_),
    .X(_04308_));
 sky130_fd_sc_hd__clkbuf_1 _16455_ (.A(_04308_),
    .X(_02023_));
 sky130_fd_sc_hd__inv_2 _16456_ (.A(_04144_),
    .Y(_04309_));
 sky130_fd_sc_hd__mux2_1 _16457_ (.A0(net815),
    .A1(_04309_),
    .S(_03957_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _16458_ (.A(_04310_),
    .X(_02024_));
 sky130_fd_sc_hd__nor2_1 _16459_ (.A(net682),
    .B(_04373_),
    .Y(_04311_));
 sky130_fd_sc_hd__a21oi_1 _16460_ (.A1(_04373_),
    .A2(_04155_),
    .B1(_04311_),
    .Y(_02025_));
 sky130_fd_sc_hd__inv_2 _16461_ (.A(_04165_),
    .Y(_04312_));
 sky130_fd_sc_hd__mux2_1 _16462_ (.A0(net819),
    .A1(_04312_),
    .S(_03957_),
    .X(_04313_));
 sky130_fd_sc_hd__clkbuf_1 _16463_ (.A(_04313_),
    .X(_02026_));
 sky130_fd_sc_hd__inv_2 _16464_ (.A(_04175_),
    .Y(_04314_));
 sky130_fd_sc_hd__mux2_1 _16465_ (.A0(net840),
    .A1(_04314_),
    .S(_03957_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _16466_ (.A(_04315_),
    .X(_02027_));
 sky130_fd_sc_hd__inv_2 _16467_ (.A(_04185_),
    .Y(_04316_));
 sky130_fd_sc_hd__mux2_1 _16468_ (.A0(\ks1.key_reg[126] ),
    .A1(_04316_),
    .S(_03957_),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_1 _16469_ (.A(_04317_),
    .X(_02028_));
 sky130_fd_sc_hd__inv_2 _16470_ (.A(_04195_),
    .Y(_04318_));
 sky130_fd_sc_hd__mux2_1 _16471_ (.A0(net849),
    .A1(_04318_),
    .S(_03957_),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _16472_ (.A(_04319_),
    .X(_02029_));
 sky130_fd_sc_hd__o21ai_1 _16473_ (.A1(net705),
    .A2(_03060_),
    .B1(_03053_),
    .Y(_02030_));
 sky130_fd_sc_hd__or2_1 _16474_ (.A(_03171_),
    .B(_03539_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_1 _16475_ (.A(_04320_),
    .X(_02031_));
 sky130_fd_sc_hd__buf_4 _16476_ (.A(_03143_),
    .X(_04321_));
 sky130_fd_sc_hd__mux2_1 _16477_ (.A0(net739),
    .A1(_03170_),
    .S(_04321_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _16478_ (.A(_04322_),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _16479_ (.A0(net759),
    .A1(_03236_),
    .S(_04321_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _16480_ (.A(_04323_),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_1 _16481_ (.A0(net722),
    .A1(_03283_),
    .S(_04321_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_1 _16482_ (.A(_04324_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _16483_ (.A0(net719),
    .A1(_03324_),
    .S(_04321_),
    .X(_04325_));
 sky130_fd_sc_hd__clkbuf_1 _16484_ (.A(_04325_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _16485_ (.A0(net709),
    .A1(_03363_),
    .S(_04321_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_1 _16486_ (.A(_04326_),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _16487_ (.A0(net784),
    .A1(_03382_),
    .S(_04321_),
    .X(_04327_));
 sky130_fd_sc_hd__clkbuf_1 _16488_ (.A(_04327_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _16489_ (.A0(net717),
    .A1(_03392_),
    .S(_04321_),
    .X(_04328_));
 sky130_fd_sc_hd__clkbuf_1 _16490_ (.A(_04328_),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _16491_ (.A0(net728),
    .A1(_03402_),
    .S(_04321_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _16492_ (.A(_04329_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _16493_ (.A0(net781),
    .A1(_03411_),
    .S(_04321_),
    .X(_04330_));
 sky130_fd_sc_hd__clkbuf_1 _16494_ (.A(_04330_),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _16495_ (.A0(net687),
    .A1(_03424_),
    .S(_04321_),
    .X(_04331_));
 sky130_fd_sc_hd__clkbuf_1 _16496_ (.A(_04331_),
    .X(_02041_));
 sky130_fd_sc_hd__buf_4 _16497_ (.A(_03143_),
    .X(_04332_));
 sky130_fd_sc_hd__mux2_1 _16498_ (.A0(net751),
    .A1(_03435_),
    .S(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__clkbuf_1 _16499_ (.A(_04333_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _16500_ (.A0(net746),
    .A1(_03446_),
    .S(_04332_),
    .X(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _16501_ (.A(_04334_),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _16502_ (.A0(net758),
    .A1(_03456_),
    .S(_04332_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _16503_ (.A(_04335_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _16504_ (.A0(net787),
    .A1(_03467_),
    .S(_04332_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _16505_ (.A(_04336_),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _16506_ (.A0(net711),
    .A1(_03477_),
    .S(_04332_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _16507_ (.A(_04337_),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_1 _16508_ (.A0(net745),
    .A1(_03484_),
    .S(_04332_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _16509_ (.A(_04338_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _16510_ (.A0(net771),
    .A1(_03487_),
    .S(_04332_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _16511_ (.A(_04339_),
    .X(_02048_));
 sky130_fd_sc_hd__mux2_1 _16512_ (.A0(net738),
    .A1(_03491_),
    .S(_04332_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _16513_ (.A(_04340_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _16514_ (.A0(net749),
    .A1(_03493_),
    .S(_04332_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _16515_ (.A(_04341_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _16516_ (.A0(net696),
    .A1(_03497_),
    .S(_04332_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _16517_ (.A(_04342_),
    .X(_02051_));
 sky130_fd_sc_hd__buf_4 _16518_ (.A(_03143_),
    .X(_04343_));
 sky130_fd_sc_hd__mux2_1 _16519_ (.A0(net688),
    .A1(_03502_),
    .S(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _16520_ (.A(_04344_),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _16521_ (.A0(net776),
    .A1(_03505_),
    .S(_04343_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_1 _16522_ (.A(_04345_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _16523_ (.A0(net779),
    .A1(_03507_),
    .S(_04343_),
    .X(_04346_));
 sky130_fd_sc_hd__clkbuf_1 _16524_ (.A(_04346_),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _16525_ (.A0(net790),
    .A1(_03510_),
    .S(_04343_),
    .X(_04347_));
 sky130_fd_sc_hd__clkbuf_1 _16526_ (.A(_04347_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _16527_ (.A0(net744),
    .A1(_03514_),
    .S(_04343_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _16528_ (.A(_04348_),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _16529_ (.A0(net757),
    .A1(_03516_),
    .S(_04343_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _16530_ (.A(_04349_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _16531_ (.A0(net684),
    .A1(_03521_),
    .S(_04343_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _16532_ (.A(_04350_),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _16533_ (.A0(net774),
    .A1(_03525_),
    .S(_04343_),
    .X(_04351_));
 sky130_fd_sc_hd__clkbuf_1 _16534_ (.A(_04351_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _16535_ (.A0(net766),
    .A1(_03527_),
    .S(_04343_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _16536_ (.A(_04352_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _16537_ (.A0(net729),
    .A1(_03529_),
    .S(_04343_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _16538_ (.A(_04353_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _16539_ (.A0(net765),
    .A1(_03533_),
    .S(_03143_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _16540_ (.A(_04354_),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _16541_ (.A0(net706),
    .A1(_03537_),
    .S(_03143_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _16542_ (.A(_04355_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _16543_ (.A0(\sub1.data_o[80] ),
    .A1(\sub1.data_o[16] ),
    .S(_03574_),
    .X(_04356_));
 sky130_fd_sc_hd__a22o_1 _16544_ (.A1(\sub1.data_o[112] ),
    .A2(_05197_),
    .B1(_04356_),
    .B2(_03594_),
    .X(_04357_));
 sky130_fd_sc_hd__a31o_1 _16545_ (.A1(_05103_),
    .A2(_04946_),
    .A3(_05548_),
    .B1(_04357_),
    .X(_02064_));
 sky130_fd_sc_hd__mux2_1 _16546_ (.A0(\sub1.data_o[81] ),
    .A1(\sub1.data_o[17] ),
    .S(_03574_),
    .X(_04358_));
 sky130_fd_sc_hd__a22o_1 _16547_ (.A1(\sub1.data_o[113] ),
    .A2(_05197_),
    .B1(_04358_),
    .B2(_03594_),
    .X(_04359_));
 sky130_fd_sc_hd__a31o_1 _16548_ (.A1(_05103_),
    .A2(_04946_),
    .A3(_05554_),
    .B1(_04359_),
    .X(_02065_));
 sky130_fd_sc_hd__mux2_1 _16549_ (.A0(\sub1.data_o[82] ),
    .A1(\sub1.data_o[18] ),
    .S(_03574_),
    .X(_04360_));
 sky130_fd_sc_hd__a22o_1 _16550_ (.A1(\sub1.data_o[114] ),
    .A2(_05197_),
    .B1(_04360_),
    .B2(_03594_),
    .X(_04361_));
 sky130_fd_sc_hd__a31o_1 _16551_ (.A1(_05103_),
    .A2(_04946_),
    .A3(_05560_),
    .B1(_04361_),
    .X(_02066_));
 sky130_fd_sc_hd__dfrtp_4 _16552_ (.CLK(clknet_leaf_28_clk),
    .D(_00000_),
    .RESET_B(net641),
    .Q(\sub1.data_o[115] ));
 sky130_fd_sc_hd__dfrtp_4 _16553_ (.CLK(clknet_leaf_21_clk),
    .D(_00001_),
    .RESET_B(net641),
    .Q(\sub1.data_o[116] ));
 sky130_fd_sc_hd__dfrtp_4 _16554_ (.CLK(clknet_leaf_28_clk),
    .D(_00002_),
    .RESET_B(net641),
    .Q(\sub1.data_o[117] ));
 sky130_fd_sc_hd__dfrtp_4 _16555_ (.CLK(clknet_leaf_28_clk),
    .D(_00003_),
    .RESET_B(net641),
    .Q(\sub1.data_o[118] ));
 sky130_fd_sc_hd__dfrtp_4 _16556_ (.CLK(clknet_leaf_28_clk),
    .D(_00004_),
    .RESET_B(net641),
    .Q(\sub1.data_o[119] ));
 sky130_fd_sc_hd__dfrtp_2 _16557_ (.CLK(clknet_leaf_54_clk),
    .D(_00005_),
    .RESET_B(net615),
    .Q(\ks1.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _16558_ (.CLK(clknet_leaf_54_clk),
    .D(_00006_),
    .RESET_B(net615),
    .Q(\ks1.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _16559_ (.CLK(clknet_leaf_49_clk),
    .D(_00007_),
    .RESET_B(net615),
    .Q(\ks1.state[2] ));
 sky130_fd_sc_hd__dfxtp_1 _16560_ (.CLK(net473),
    .D(_00008_),
    .Q(\fifo_bank_register.bank[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16561_ (.CLK(net490),
    .D(_00009_),
    .Q(\fifo_bank_register.bank[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16562_ (.CLK(net474),
    .D(_00010_),
    .Q(\fifo_bank_register.bank[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16563_ (.CLK(net473),
    .D(_00011_),
    .Q(\fifo_bank_register.bank[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16564_ (.CLK(net474),
    .D(_00012_),
    .Q(\fifo_bank_register.bank[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16565_ (.CLK(net473),
    .D(_00013_),
    .Q(\fifo_bank_register.bank[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16566_ (.CLK(net477),
    .D(_00014_),
    .Q(\fifo_bank_register.bank[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16567_ (.CLK(net477),
    .D(_00015_),
    .Q(\fifo_bank_register.bank[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16568_ (.CLK(net478),
    .D(_00016_),
    .Q(\fifo_bank_register.bank[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16569_ (.CLK(net478),
    .D(_00017_),
    .Q(\fifo_bank_register.bank[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16570_ (.CLK(net504),
    .D(_00018_),
    .Q(\fifo_bank_register.bank[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16571_ (.CLK(net533),
    .D(_00019_),
    .Q(\fifo_bank_register.bank[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16572_ (.CLK(net504),
    .D(_00020_),
    .Q(\fifo_bank_register.bank[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16573_ (.CLK(net505),
    .D(_00021_),
    .Q(\fifo_bank_register.bank[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16574_ (.CLK(net534),
    .D(_00022_),
    .Q(\fifo_bank_register.bank[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16575_ (.CLK(net534),
    .D(_00023_),
    .Q(\fifo_bank_register.bank[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16576_ (.CLK(net496),
    .D(_00024_),
    .Q(\fifo_bank_register.bank[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _16577_ (.CLK(net532),
    .D(_00025_),
    .Q(\fifo_bank_register.bank[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _16578_ (.CLK(net533),
    .D(_00026_),
    .Q(\fifo_bank_register.bank[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _16579_ (.CLK(net505),
    .D(_00027_),
    .Q(\fifo_bank_register.bank[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _16580_ (.CLK(net512),
    .D(_00028_),
    .Q(\fifo_bank_register.bank[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _16581_ (.CLK(net484),
    .D(_00029_),
    .Q(\fifo_bank_register.bank[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _16582_ (.CLK(net501),
    .D(_00030_),
    .Q(\fifo_bank_register.bank[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _16583_ (.CLK(net484),
    .D(_00031_),
    .Q(\fifo_bank_register.bank[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _16584_ (.CLK(net482),
    .D(_00032_),
    .Q(\fifo_bank_register.bank[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _16585_ (.CLK(net508),
    .D(_00033_),
    .Q(\fifo_bank_register.bank[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _16586_ (.CLK(net510),
    .D(_00034_),
    .Q(\fifo_bank_register.bank[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _16587_ (.CLK(net486),
    .D(_00035_),
    .Q(\fifo_bank_register.bank[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _16588_ (.CLK(net486),
    .D(_00036_),
    .Q(\fifo_bank_register.bank[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _16589_ (.CLK(net499),
    .D(_00037_),
    .Q(\fifo_bank_register.bank[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _16590_ (.CLK(net437),
    .D(_00038_),
    .Q(\fifo_bank_register.bank[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _16591_ (.CLK(net437),
    .D(_00039_),
    .Q(\fifo_bank_register.bank[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _16592_ (.CLK(net423),
    .D(_00040_),
    .Q(\fifo_bank_register.bank[9][32] ));
 sky130_fd_sc_hd__dfxtp_1 _16593_ (.CLK(net423),
    .D(_00041_),
    .Q(\fifo_bank_register.bank[9][33] ));
 sky130_fd_sc_hd__dfxtp_1 _16594_ (.CLK(net430),
    .D(_00042_),
    .Q(\fifo_bank_register.bank[9][34] ));
 sky130_fd_sc_hd__dfxtp_1 _16595_ (.CLK(net428),
    .D(_00043_),
    .Q(\fifo_bank_register.bank[9][35] ));
 sky130_fd_sc_hd__dfxtp_1 _16596_ (.CLK(net423),
    .D(_00044_),
    .Q(\fifo_bank_register.bank[9][36] ));
 sky130_fd_sc_hd__dfxtp_1 _16597_ (.CLK(net417),
    .D(_00045_),
    .Q(\fifo_bank_register.bank[9][37] ));
 sky130_fd_sc_hd__dfxtp_1 _16598_ (.CLK(net428),
    .D(_00046_),
    .Q(\fifo_bank_register.bank[9][38] ));
 sky130_fd_sc_hd__dfxtp_1 _16599_ (.CLK(net415),
    .D(_00047_),
    .Q(\fifo_bank_register.bank[9][39] ));
 sky130_fd_sc_hd__dfxtp_1 _16600_ (.CLK(net395),
    .D(_00048_),
    .Q(\fifo_bank_register.bank[9][40] ));
 sky130_fd_sc_hd__dfxtp_1 _16601_ (.CLK(net398),
    .D(_00049_),
    .Q(\fifo_bank_register.bank[9][41] ));
 sky130_fd_sc_hd__dfxtp_1 _16602_ (.CLK(net405),
    .D(_00050_),
    .Q(\fifo_bank_register.bank[9][42] ));
 sky130_fd_sc_hd__dfxtp_1 _16603_ (.CLK(net393),
    .D(_00051_),
    .Q(\fifo_bank_register.bank[9][43] ));
 sky130_fd_sc_hd__dfxtp_1 _16604_ (.CLK(net389),
    .D(_00052_),
    .Q(\fifo_bank_register.bank[9][44] ));
 sky130_fd_sc_hd__dfxtp_1 _16605_ (.CLK(net405),
    .D(_00053_),
    .Q(\fifo_bank_register.bank[9][45] ));
 sky130_fd_sc_hd__dfxtp_1 _16606_ (.CLK(net394),
    .D(_00054_),
    .Q(\fifo_bank_register.bank[9][46] ));
 sky130_fd_sc_hd__dfxtp_1 _16607_ (.CLK(net396),
    .D(_00055_),
    .Q(\fifo_bank_register.bank[9][47] ));
 sky130_fd_sc_hd__dfxtp_1 _16608_ (.CLK(net395),
    .D(_00056_),
    .Q(\fifo_bank_register.bank[9][48] ));
 sky130_fd_sc_hd__dfxtp_1 _16609_ (.CLK(net407),
    .D(_00057_),
    .Q(\fifo_bank_register.bank[9][49] ));
 sky130_fd_sc_hd__dfxtp_1 _16610_ (.CLK(net557),
    .D(_00058_),
    .Q(\fifo_bank_register.bank[9][50] ));
 sky130_fd_sc_hd__dfxtp_1 _16611_ (.CLK(net573),
    .D(_00059_),
    .Q(\fifo_bank_register.bank[9][51] ));
 sky130_fd_sc_hd__dfxtp_1 _16612_ (.CLK(net563),
    .D(_00060_),
    .Q(\fifo_bank_register.bank[9][52] ));
 sky130_fd_sc_hd__dfxtp_1 _16613_ (.CLK(net562),
    .D(_00061_),
    .Q(\fifo_bank_register.bank[9][53] ));
 sky130_fd_sc_hd__dfxtp_1 _16614_ (.CLK(net556),
    .D(_00062_),
    .Q(\fifo_bank_register.bank[9][54] ));
 sky130_fd_sc_hd__dfxtp_1 _16615_ (.CLK(net572),
    .D(_00063_),
    .Q(\fifo_bank_register.bank[9][55] ));
 sky130_fd_sc_hd__dfxtp_1 _16616_ (.CLK(net574),
    .D(_00064_),
    .Q(\fifo_bank_register.bank[9][56] ));
 sky130_fd_sc_hd__dfxtp_1 _16617_ (.CLK(net550),
    .D(_00065_),
    .Q(\fifo_bank_register.bank[9][57] ));
 sky130_fd_sc_hd__dfxtp_1 _16618_ (.CLK(net557),
    .D(_00066_),
    .Q(\fifo_bank_register.bank[9][58] ));
 sky130_fd_sc_hd__dfxtp_1 _16619_ (.CLK(net572),
    .D(_00067_),
    .Q(\fifo_bank_register.bank[9][59] ));
 sky130_fd_sc_hd__dfxtp_1 _16620_ (.CLK(net515),
    .D(_00068_),
    .Q(\fifo_bank_register.bank[9][60] ));
 sky130_fd_sc_hd__dfxtp_1 _16621_ (.CLK(net527),
    .D(_00069_),
    .Q(\fifo_bank_register.bank[9][61] ));
 sky130_fd_sc_hd__dfxtp_1 _16622_ (.CLK(net523),
    .D(_00070_),
    .Q(\fifo_bank_register.bank[9][62] ));
 sky130_fd_sc_hd__dfxtp_1 _16623_ (.CLK(net524),
    .D(_00071_),
    .Q(\fifo_bank_register.bank[9][63] ));
 sky130_fd_sc_hd__dfxtp_1 _16624_ (.CLK(net514),
    .D(_00072_),
    .Q(\fifo_bank_register.bank[9][64] ));
 sky130_fd_sc_hd__dfxtp_1 _16625_ (.CLK(net526),
    .D(_00073_),
    .Q(\fifo_bank_register.bank[9][65] ));
 sky130_fd_sc_hd__dfxtp_1 _16626_ (.CLK(net527),
    .D(_00074_),
    .Q(\fifo_bank_register.bank[9][66] ));
 sky130_fd_sc_hd__dfxtp_1 _16627_ (.CLK(net521),
    .D(_00075_),
    .Q(\fifo_bank_register.bank[9][67] ));
 sky130_fd_sc_hd__dfxtp_1 _16628_ (.CLK(net511),
    .D(_00076_),
    .Q(\fifo_bank_register.bank[9][68] ));
 sky130_fd_sc_hd__dfxtp_1 _16629_ (.CLK(net518),
    .D(_00077_),
    .Q(\fifo_bank_register.bank[9][69] ));
 sky130_fd_sc_hd__dfxtp_1 _16630_ (.CLK(net519),
    .D(_00078_),
    .Q(\fifo_bank_register.bank[9][70] ));
 sky130_fd_sc_hd__dfxtp_1 _16631_ (.CLK(net528),
    .D(_00079_),
    .Q(\fifo_bank_register.bank[9][71] ));
 sky130_fd_sc_hd__dfxtp_1 _16632_ (.CLK(net553),
    .D(_00080_),
    .Q(\fifo_bank_register.bank[9][72] ));
 sky130_fd_sc_hd__dfxtp_1 _16633_ (.CLK(net554),
    .D(_00081_),
    .Q(\fifo_bank_register.bank[9][73] ));
 sky130_fd_sc_hd__dfxtp_1 _16634_ (.CLK(net549),
    .D(_00082_),
    .Q(\fifo_bank_register.bank[9][74] ));
 sky130_fd_sc_hd__dfxtp_1 _16635_ (.CLK(net552),
    .D(_00083_),
    .Q(\fifo_bank_register.bank[9][75] ));
 sky130_fd_sc_hd__dfxtp_1 _16636_ (.CLK(net545),
    .D(_00084_),
    .Q(\fifo_bank_register.bank[9][76] ));
 sky130_fd_sc_hd__dfxtp_1 _16637_ (.CLK(net554),
    .D(_00085_),
    .Q(\fifo_bank_register.bank[9][77] ));
 sky130_fd_sc_hd__dfxtp_1 _16638_ (.CLK(net525),
    .D(_00086_),
    .Q(\fifo_bank_register.bank[9][78] ));
 sky130_fd_sc_hd__dfxtp_1 _16639_ (.CLK(net555),
    .D(_00087_),
    .Q(\fifo_bank_register.bank[9][79] ));
 sky130_fd_sc_hd__dfxtp_1 _16640_ (.CLK(net565),
    .D(_00088_),
    .Q(\fifo_bank_register.bank[9][80] ));
 sky130_fd_sc_hd__dfxtp_1 _16641_ (.CLK(net563),
    .D(_00089_),
    .Q(\fifo_bank_register.bank[9][81] ));
 sky130_fd_sc_hd__dfxtp_1 _16642_ (.CLK(net560),
    .D(_00090_),
    .Q(\fifo_bank_register.bank[9][82] ));
 sky130_fd_sc_hd__dfxtp_1 _16643_ (.CLK(net561),
    .D(_00091_),
    .Q(\fifo_bank_register.bank[9][83] ));
 sky130_fd_sc_hd__dfxtp_1 _16644_ (.CLK(net550),
    .D(_00092_),
    .Q(\fifo_bank_register.bank[9][84] ));
 sky130_fd_sc_hd__dfxtp_1 _16645_ (.CLK(net567),
    .D(_00093_),
    .Q(\fifo_bank_register.bank[9][85] ));
 sky130_fd_sc_hd__dfxtp_1 _16646_ (.CLK(net560),
    .D(_00094_),
    .Q(\fifo_bank_register.bank[9][86] ));
 sky130_fd_sc_hd__dfxtp_1 _16647_ (.CLK(net561),
    .D(_00095_),
    .Q(\fifo_bank_register.bank[9][87] ));
 sky130_fd_sc_hd__dfxtp_1 _16648_ (.CLK(net565),
    .D(_00096_),
    .Q(\fifo_bank_register.bank[9][88] ));
 sky130_fd_sc_hd__dfxtp_1 _16649_ (.CLK(net547),
    .D(_00097_),
    .Q(\fifo_bank_register.bank[9][89] ));
 sky130_fd_sc_hd__dfxtp_1 _16650_ (.CLK(net409),
    .D(_00098_),
    .Q(\fifo_bank_register.bank[9][90] ));
 sky130_fd_sc_hd__dfxtp_1 _16651_ (.CLK(net403),
    .D(_00099_),
    .Q(\fifo_bank_register.bank[9][91] ));
 sky130_fd_sc_hd__dfxtp_1 _16652_ (.CLK(net410),
    .D(_00100_),
    .Q(\fifo_bank_register.bank[9][92] ));
 sky130_fd_sc_hd__dfxtp_1 _16653_ (.CLK(net402),
    .D(_00101_),
    .Q(\fifo_bank_register.bank[9][93] ));
 sky130_fd_sc_hd__dfxtp_1 _16654_ (.CLK(net455),
    .D(_00102_),
    .Q(\fifo_bank_register.bank[9][94] ));
 sky130_fd_sc_hd__dfxtp_1 _16655_ (.CLK(net402),
    .D(_00103_),
    .Q(\fifo_bank_register.bank[9][95] ));
 sky130_fd_sc_hd__dfxtp_1 _16656_ (.CLK(net403),
    .D(_00104_),
    .Q(\fifo_bank_register.bank[9][96] ));
 sky130_fd_sc_hd__dfxtp_1 _16657_ (.CLK(net454),
    .D(_00105_),
    .Q(\fifo_bank_register.bank[9][97] ));
 sky130_fd_sc_hd__dfxtp_1 _16658_ (.CLK(net449),
    .D(_00106_),
    .Q(\fifo_bank_register.bank[9][98] ));
 sky130_fd_sc_hd__dfxtp_1 _16659_ (.CLK(net447),
    .D(_00107_),
    .Q(\fifo_bank_register.bank[9][99] ));
 sky130_fd_sc_hd__dfxtp_1 _16660_ (.CLK(net452),
    .D(_00108_),
    .Q(\fifo_bank_register.bank[9][100] ));
 sky130_fd_sc_hd__dfxtp_1 _16661_ (.CLK(net450),
    .D(_00109_),
    .Q(\fifo_bank_register.bank[9][101] ));
 sky130_fd_sc_hd__dfxtp_1 _16662_ (.CLK(net465),
    .D(_00110_),
    .Q(\fifo_bank_register.bank[9][102] ));
 sky130_fd_sc_hd__dfxtp_1 _16663_ (.CLK(net458),
    .D(_00111_),
    .Q(\fifo_bank_register.bank[9][103] ));
 sky130_fd_sc_hd__dfxtp_1 _16664_ (.CLK(net463),
    .D(_00112_),
    .Q(\fifo_bank_register.bank[9][104] ));
 sky130_fd_sc_hd__dfxtp_1 _16665_ (.CLK(net468),
    .D(_00113_),
    .Q(\fifo_bank_register.bank[9][105] ));
 sky130_fd_sc_hd__dfxtp_1 _16666_ (.CLK(net465),
    .D(_00114_),
    .Q(\fifo_bank_register.bank[9][106] ));
 sky130_fd_sc_hd__dfxtp_1 _16667_ (.CLK(net451),
    .D(_00115_),
    .Q(\fifo_bank_register.bank[9][107] ));
 sky130_fd_sc_hd__dfxtp_1 _16668_ (.CLK(net453),
    .D(_00116_),
    .Q(\fifo_bank_register.bank[9][108] ));
 sky130_fd_sc_hd__dfxtp_1 _16669_ (.CLK(net458),
    .D(_00117_),
    .Q(\fifo_bank_register.bank[9][109] ));
 sky130_fd_sc_hd__dfxtp_1 _16670_ (.CLK(net471),
    .D(_00118_),
    .Q(\fifo_bank_register.bank[9][110] ));
 sky130_fd_sc_hd__dfxtp_1 _16671_ (.CLK(net413),
    .D(_00119_),
    .Q(\fifo_bank_register.bank[9][111] ));
 sky130_fd_sc_hd__dfxtp_1 _16672_ (.CLK(net433),
    .D(_00120_),
    .Q(\fifo_bank_register.bank[9][112] ));
 sky130_fd_sc_hd__dfxtp_1 _16673_ (.CLK(net469),
    .D(_00121_),
    .Q(\fifo_bank_register.bank[9][113] ));
 sky130_fd_sc_hd__dfxtp_1 _16674_ (.CLK(net456),
    .D(_00122_),
    .Q(\fifo_bank_register.bank[9][114] ));
 sky130_fd_sc_hd__dfxtp_1 _16675_ (.CLK(net470),
    .D(_00123_),
    .Q(\fifo_bank_register.bank[9][115] ));
 sky130_fd_sc_hd__dfxtp_1 _16676_ (.CLK(net411),
    .D(_00124_),
    .Q(\fifo_bank_register.bank[9][116] ));
 sky130_fd_sc_hd__dfxtp_1 _16677_ (.CLK(net435),
    .D(_00125_),
    .Q(\fifo_bank_register.bank[9][117] ));
 sky130_fd_sc_hd__dfxtp_1 _16678_ (.CLK(net456),
    .D(_00126_),
    .Q(\fifo_bank_register.bank[9][118] ));
 sky130_fd_sc_hd__dfxtp_1 _16679_ (.CLK(net435),
    .D(_00127_),
    .Q(\fifo_bank_register.bank[9][119] ));
 sky130_fd_sc_hd__dfxtp_1 _16680_ (.CLK(net441),
    .D(_00128_),
    .Q(\fifo_bank_register.bank[9][120] ));
 sky130_fd_sc_hd__dfxtp_1 _16681_ (.CLK(net490),
    .D(_00129_),
    .Q(\fifo_bank_register.bank[9][121] ));
 sky130_fd_sc_hd__dfxtp_1 _16682_ (.CLK(net493),
    .D(_00130_),
    .Q(\fifo_bank_register.bank[9][122] ));
 sky130_fd_sc_hd__dfxtp_1 _16683_ (.CLK(net439),
    .D(_00131_),
    .Q(\fifo_bank_register.bank[9][123] ));
 sky130_fd_sc_hd__dfxtp_1 _16684_ (.CLK(net495),
    .D(_00132_),
    .Q(\fifo_bank_register.bank[9][124] ));
 sky130_fd_sc_hd__dfxtp_1 _16685_ (.CLK(net497),
    .D(_00133_),
    .Q(\fifo_bank_register.bank[9][125] ));
 sky130_fd_sc_hd__dfxtp_1 _16686_ (.CLK(net495),
    .D(_00134_),
    .Q(\fifo_bank_register.bank[9][126] ));
 sky130_fd_sc_hd__dfxtp_1 _16687_ (.CLK(net443),
    .D(_00135_),
    .Q(\fifo_bank_register.bank[9][127] ));
 sky130_fd_sc_hd__dfrtp_1 _16688_ (.CLK(clknet_leaf_49_clk),
    .D(\ks1.next_ready_o ),
    .RESET_B(net615),
    .Q(\ks1.ready_o ));
 sky130_fd_sc_hd__dfrtp_4 _16689_ (.CLK(clknet_leaf_50_clk),
    .D(_00136_),
    .RESET_B(net615),
    .Q(\addroundkey_round[0] ));
 sky130_fd_sc_hd__dfrtp_4 _16690_ (.CLK(clknet_leaf_54_clk),
    .D(_00137_),
    .RESET_B(net616),
    .Q(\addroundkey_round[1] ));
 sky130_fd_sc_hd__dfrtp_4 _16691_ (.CLK(clknet_leaf_50_clk),
    .D(_00138_),
    .RESET_B(net616),
    .Q(\addroundkey_round[2] ));
 sky130_fd_sc_hd__dfrtp_4 _16692_ (.CLK(clknet_leaf_50_clk),
    .D(_00139_),
    .RESET_B(net616),
    .Q(\addroundkey_round[3] ));
 sky130_fd_sc_hd__dfrtp_1 _16693_ (.CLK(clknet_leaf_5_clk),
    .D(_00140_),
    .RESET_B(net592),
    .Q(\sub1.data_o[120] ));
 sky130_fd_sc_hd__dfrtp_2 _16694_ (.CLK(clknet_leaf_72_clk),
    .D(_00141_),
    .RESET_B(net594),
    .Q(\sub1.data_o[121] ));
 sky130_fd_sc_hd__dfrtp_1 _16695_ (.CLK(clknet_leaf_5_clk),
    .D(_00142_),
    .RESET_B(net592),
    .Q(\sub1.data_o[122] ));
 sky130_fd_sc_hd__dfrtp_4 _16696_ (.CLK(clknet_leaf_72_clk),
    .D(_00143_),
    .RESET_B(net594),
    .Q(\sub1.data_o[123] ));
 sky130_fd_sc_hd__dfrtp_4 _16697_ (.CLK(clknet_leaf_71_clk),
    .D(_00144_),
    .RESET_B(net608),
    .Q(\sub1.data_o[124] ));
 sky130_fd_sc_hd__dfrtp_1 _16698_ (.CLK(clknet_leaf_71_clk),
    .D(_00145_),
    .RESET_B(net652),
    .Q(\sub1.data_o[125] ));
 sky130_fd_sc_hd__dfrtp_2 _16699_ (.CLK(clknet_leaf_72_clk),
    .D(_00146_),
    .RESET_B(net635),
    .Q(\sub1.data_o[126] ));
 sky130_fd_sc_hd__dfrtp_2 _16700_ (.CLK(clknet_leaf_71_clk),
    .D(_00147_),
    .RESET_B(net652),
    .Q(\sub1.data_o[127] ));
 sky130_fd_sc_hd__dfrtp_2 _16701_ (.CLK(clknet_leaf_44_clk),
    .D(next_state),
    .RESET_B(net653),
    .Q(state));
 sky130_fd_sc_hd__dfrtp_4 _16702_ (.CLK(clknet_leaf_40_clk),
    .D(_00148_),
    .RESET_B(net669),
    .Q(net388));
 sky130_fd_sc_hd__dfrtp_2 _16703_ (.CLK(clknet_leaf_40_clk),
    .D(_00149_),
    .RESET_B(net669),
    .Q(\round[0] ));
 sky130_fd_sc_hd__dfrtp_4 _16704_ (.CLK(clknet_leaf_40_clk),
    .D(_00150_),
    .RESET_B(net669),
    .Q(\round[1] ));
 sky130_fd_sc_hd__dfrtp_4 _16705_ (.CLK(clknet_leaf_40_clk),
    .D(_00151_),
    .RESET_B(net669),
    .Q(\round[2] ));
 sky130_fd_sc_hd__dfrtp_4 _16706_ (.CLK(clknet_leaf_40_clk),
    .D(_00152_),
    .RESET_B(net669),
    .Q(\round[3] ));
 sky130_fd_sc_hd__dfrtp_4 _16707_ (.CLK(clknet_leaf_44_clk),
    .D(next_addroundkey_ready_o),
    .RESET_B(net658),
    .Q(addroundkey_ready_o));
 sky130_fd_sc_hd__dfrtp_4 _16708_ (.CLK(clknet_leaf_44_clk),
    .D(next_addroundkey_start_i),
    .RESET_B(net658),
    .Q(addroundkey_start_i));
 sky130_fd_sc_hd__dfrtp_4 _16709_ (.CLK(clknet_leaf_50_clk),
    .D(_00153_),
    .RESET_B(net616),
    .Q(\addroundkey_data_o[0] ));
 sky130_fd_sc_hd__dfrtp_4 _16710_ (.CLK(clknet_leaf_41_clk),
    .D(_00154_),
    .RESET_B(net658),
    .Q(\addroundkey_data_o[1] ));
 sky130_fd_sc_hd__dfrtp_4 _16711_ (.CLK(clknet_leaf_51_clk),
    .D(_00155_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[2] ));
 sky130_fd_sc_hd__dfrtp_4 _16712_ (.CLK(clknet_leaf_51_clk),
    .D(_00156_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[3] ));
 sky130_fd_sc_hd__dfrtp_4 _16713_ (.CLK(clknet_leaf_51_clk),
    .D(_00157_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[4] ));
 sky130_fd_sc_hd__dfrtp_4 _16714_ (.CLK(clknet_leaf_41_clk),
    .D(_00158_),
    .RESET_B(net658),
    .Q(\addroundkey_data_o[5] ));
 sky130_fd_sc_hd__dfrtp_4 _16715_ (.CLK(clknet_leaf_51_clk),
    .D(_00159_),
    .RESET_B(net651),
    .Q(\addroundkey_data_o[6] ));
 sky130_fd_sc_hd__dfrtp_4 _16716_ (.CLK(clknet_leaf_49_clk),
    .D(_00160_),
    .RESET_B(net616),
    .Q(\addroundkey_data_o[7] ));
 sky130_fd_sc_hd__dfrtp_4 _16717_ (.CLK(clknet_leaf_51_clk),
    .D(_00161_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[8] ));
 sky130_fd_sc_hd__dfrtp_4 _16718_ (.CLK(clknet_leaf_43_clk),
    .D(_00162_),
    .RESET_B(net658),
    .Q(\addroundkey_data_o[9] ));
 sky130_fd_sc_hd__dfrtp_4 _16719_ (.CLK(clknet_leaf_51_clk),
    .D(_00163_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[10] ));
 sky130_fd_sc_hd__dfrtp_4 _16720_ (.CLK(clknet_leaf_52_clk),
    .D(_00164_),
    .RESET_B(net656),
    .Q(\addroundkey_data_o[11] ));
 sky130_fd_sc_hd__dfrtp_4 _16721_ (.CLK(clknet_leaf_52_clk),
    .D(_00165_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[12] ));
 sky130_fd_sc_hd__dfrtp_4 _16722_ (.CLK(clknet_leaf_42_clk),
    .D(_00166_),
    .RESET_B(net659),
    .Q(\addroundkey_data_o[13] ));
 sky130_fd_sc_hd__dfrtp_4 _16723_ (.CLK(clknet_leaf_43_clk),
    .D(_00167_),
    .RESET_B(net655),
    .Q(\addroundkey_data_o[14] ));
 sky130_fd_sc_hd__dfrtp_4 _16724_ (.CLK(clknet_leaf_42_clk),
    .D(_00168_),
    .RESET_B(net659),
    .Q(\addroundkey_data_o[15] ));
 sky130_fd_sc_hd__dfrtp_4 _16725_ (.CLK(clknet_leaf_41_clk),
    .D(_00169_),
    .RESET_B(net658),
    .Q(\addroundkey_data_o[16] ));
 sky130_fd_sc_hd__dfrtp_4 _16726_ (.CLK(clknet_leaf_41_clk),
    .D(_00170_),
    .RESET_B(net658),
    .Q(\addroundkey_data_o[17] ));
 sky130_fd_sc_hd__dfrtp_4 _16727_ (.CLK(clknet_leaf_40_clk),
    .D(_00171_),
    .RESET_B(net659),
    .Q(\addroundkey_data_o[18] ));
 sky130_fd_sc_hd__dfrtp_4 _16728_ (.CLK(clknet_leaf_41_clk),
    .D(_00172_),
    .RESET_B(net659),
    .Q(\addroundkey_data_o[19] ));
 sky130_fd_sc_hd__dfrtp_4 _16729_ (.CLK(clknet_leaf_43_clk),
    .D(_00173_),
    .RESET_B(net658),
    .Q(\addroundkey_data_o[20] ));
 sky130_fd_sc_hd__dfrtp_4 _16730_ (.CLK(clknet_leaf_41_clk),
    .D(_00174_),
    .RESET_B(net659),
    .Q(\addroundkey_data_o[21] ));
 sky130_fd_sc_hd__dfrtp_4 _16731_ (.CLK(clknet_leaf_42_clk),
    .D(_00175_),
    .RESET_B(net659),
    .Q(\addroundkey_data_o[22] ));
 sky130_fd_sc_hd__dfrtp_4 _16732_ (.CLK(clknet_leaf_43_clk),
    .D(_00176_),
    .RESET_B(net658),
    .Q(\addroundkey_data_o[23] ));
 sky130_fd_sc_hd__dfrtp_4 _16733_ (.CLK(clknet_leaf_51_clk),
    .D(_00177_),
    .RESET_B(net616),
    .Q(\addroundkey_data_o[24] ));
 sky130_fd_sc_hd__dfrtp_4 _16734_ (.CLK(clknet_leaf_50_clk),
    .D(_00178_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[25] ));
 sky130_fd_sc_hd__dfrtp_4 _16735_ (.CLK(clknet_leaf_52_clk),
    .D(_00179_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[26] ));
 sky130_fd_sc_hd__dfrtp_2 _16736_ (.CLK(clknet_leaf_43_clk),
    .D(_00180_),
    .RESET_B(net655),
    .Q(\addroundkey_data_o[27] ));
 sky130_fd_sc_hd__dfrtp_4 _16737_ (.CLK(clknet_leaf_52_clk),
    .D(_00181_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[28] ));
 sky130_fd_sc_hd__dfrtp_4 _16738_ (.CLK(clknet_leaf_51_clk),
    .D(_00182_),
    .RESET_B(net654),
    .Q(\addroundkey_data_o[29] ));
 sky130_fd_sc_hd__dfrtp_4 _16739_ (.CLK(clknet_leaf_47_clk),
    .D(_00183_),
    .RESET_B(net653),
    .Q(\addroundkey_data_o[30] ));
 sky130_fd_sc_hd__dfrtp_4 _16740_ (.CLK(clknet_leaf_47_clk),
    .D(_00184_),
    .RESET_B(net651),
    .Q(\addroundkey_data_o[31] ));
 sky130_fd_sc_hd__dfrtp_4 _16741_ (.CLK(clknet_leaf_47_clk),
    .D(_00185_),
    .RESET_B(net651),
    .Q(\addroundkey_data_o[32] ));
 sky130_fd_sc_hd__dfrtp_4 _16742_ (.CLK(clknet_leaf_47_clk),
    .D(_00186_),
    .RESET_B(net611),
    .Q(\addroundkey_data_o[33] ));
 sky130_fd_sc_hd__dfrtp_4 _16743_ (.CLK(clknet_leaf_48_clk),
    .D(_00187_),
    .RESET_B(net611),
    .Q(\addroundkey_data_o[34] ));
 sky130_fd_sc_hd__dfrtp_2 _16744_ (.CLK(clknet_leaf_45_clk),
    .D(_00188_),
    .RESET_B(net653),
    .Q(\addroundkey_data_o[35] ));
 sky130_fd_sc_hd__dfrtp_4 _16745_ (.CLK(clknet_leaf_48_clk),
    .D(_00189_),
    .RESET_B(net611),
    .Q(\addroundkey_data_o[36] ));
 sky130_fd_sc_hd__dfrtp_4 _16746_ (.CLK(clknet_leaf_45_clk),
    .D(_00190_),
    .RESET_B(net653),
    .Q(\addroundkey_data_o[37] ));
 sky130_fd_sc_hd__dfrtp_4 _16747_ (.CLK(clknet_leaf_45_clk),
    .D(_00191_),
    .RESET_B(net653),
    .Q(\addroundkey_data_o[38] ));
 sky130_fd_sc_hd__dfrtp_4 _16748_ (.CLK(clknet_leaf_65_clk),
    .D(_00192_),
    .RESET_B(net604),
    .Q(\addroundkey_data_o[39] ));
 sky130_fd_sc_hd__dfrtp_4 _16749_ (.CLK(clknet_leaf_68_clk),
    .D(_00193_),
    .RESET_B(net608),
    .Q(\addroundkey_data_o[40] ));
 sky130_fd_sc_hd__dfrtp_4 _16750_ (.CLK(clknet_leaf_70_clk),
    .D(_00194_),
    .RESET_B(net609),
    .Q(\addroundkey_data_o[41] ));
 sky130_fd_sc_hd__dfrtp_4 _16751_ (.CLK(clknet_leaf_70_clk),
    .D(_00195_),
    .RESET_B(net608),
    .Q(\addroundkey_data_o[42] ));
 sky130_fd_sc_hd__dfrtp_2 _16752_ (.CLK(clknet_leaf_70_clk),
    .D(_00196_),
    .RESET_B(net609),
    .Q(\addroundkey_data_o[43] ));
 sky130_fd_sc_hd__dfrtp_4 _16753_ (.CLK(clknet_leaf_65_clk),
    .D(_00197_),
    .RESET_B(net603),
    .Q(\addroundkey_data_o[44] ));
 sky130_fd_sc_hd__dfrtp_4 _16754_ (.CLK(clknet_leaf_64_clk),
    .D(_00198_),
    .RESET_B(net603),
    .Q(\addroundkey_data_o[45] ));
 sky130_fd_sc_hd__dfrtp_4 _16755_ (.CLK(clknet_leaf_66_clk),
    .D(_00199_),
    .RESET_B(net603),
    .Q(\addroundkey_data_o[46] ));
 sky130_fd_sc_hd__dfrtp_4 _16756_ (.CLK(clknet_leaf_66_clk),
    .D(_00200_),
    .RESET_B(net604),
    .Q(\addroundkey_data_o[47] ));
 sky130_fd_sc_hd__dfrtp_4 _16757_ (.CLK(clknet_leaf_66_clk),
    .D(_00201_),
    .RESET_B(net603),
    .Q(\addroundkey_data_o[48] ));
 sky130_fd_sc_hd__dfrtp_4 _16758_ (.CLK(clknet_leaf_39_clk),
    .D(_00202_),
    .RESET_B(net668),
    .Q(\addroundkey_data_o[49] ));
 sky130_fd_sc_hd__dfrtp_4 _16759_ (.CLK(clknet_leaf_39_clk),
    .D(_00203_),
    .RESET_B(net663),
    .Q(\addroundkey_data_o[50] ));
 sky130_fd_sc_hd__dfrtp_4 _16760_ (.CLK(clknet_leaf_39_clk),
    .D(_00204_),
    .RESET_B(net663),
    .Q(\addroundkey_data_o[51] ));
 sky130_fd_sc_hd__dfrtp_4 _16761_ (.CLK(clknet_leaf_68_clk),
    .D(_00205_),
    .RESET_B(net609),
    .Q(\addroundkey_data_o[52] ));
 sky130_fd_sc_hd__dfrtp_2 _16762_ (.CLK(clknet_leaf_38_clk),
    .D(_00206_),
    .RESET_B(net668),
    .Q(\addroundkey_data_o[53] ));
 sky130_fd_sc_hd__dfrtp_4 _16763_ (.CLK(clknet_leaf_70_clk),
    .D(_00207_),
    .RESET_B(net608),
    .Q(\addroundkey_data_o[54] ));
 sky130_fd_sc_hd__dfrtp_4 _16764_ (.CLK(clknet_leaf_39_clk),
    .D(_00208_),
    .RESET_B(net668),
    .Q(\addroundkey_data_o[55] ));
 sky130_fd_sc_hd__dfrtp_4 _16765_ (.CLK(clknet_leaf_48_clk),
    .D(_00209_),
    .RESET_B(net611),
    .Q(\addroundkey_data_o[56] ));
 sky130_fd_sc_hd__dfrtp_4 _16766_ (.CLK(clknet_leaf_48_clk),
    .D(_00210_),
    .RESET_B(net610),
    .Q(\addroundkey_data_o[57] ));
 sky130_fd_sc_hd__dfrtp_4 _16767_ (.CLK(clknet_leaf_68_clk),
    .D(_00211_),
    .RESET_B(net611),
    .Q(\addroundkey_data_o[58] ));
 sky130_fd_sc_hd__dfrtp_2 _16768_ (.CLK(clknet_leaf_47_clk),
    .D(_00212_),
    .RESET_B(net651),
    .Q(\addroundkey_data_o[59] ));
 sky130_fd_sc_hd__dfrtp_4 _16769_ (.CLK(clknet_leaf_48_clk),
    .D(_00213_),
    .RESET_B(net611),
    .Q(\addroundkey_data_o[60] ));
 sky130_fd_sc_hd__dfrtp_4 _16770_ (.CLK(clknet_leaf_48_clk),
    .D(_00214_),
    .RESET_B(net610),
    .Q(\addroundkey_data_o[61] ));
 sky130_fd_sc_hd__dfrtp_4 _16771_ (.CLK(clknet_leaf_48_clk),
    .D(_00215_),
    .RESET_B(net611),
    .Q(\addroundkey_data_o[62] ));
 sky130_fd_sc_hd__dfrtp_4 _16772_ (.CLK(clknet_leaf_47_clk),
    .D(_00216_),
    .RESET_B(net651),
    .Q(\addroundkey_data_o[63] ));
 sky130_fd_sc_hd__dfrtp_4 _16773_ (.CLK(clknet_leaf_67_clk),
    .D(_00217_),
    .RESET_B(net610),
    .Q(\addroundkey_data_o[64] ));
 sky130_fd_sc_hd__dfrtp_4 _16774_ (.CLK(clknet_leaf_47_clk),
    .D(_00218_),
    .RESET_B(net651),
    .Q(\addroundkey_data_o[65] ));
 sky130_fd_sc_hd__dfrtp_4 _16775_ (.CLK(clknet_leaf_67_clk),
    .D(_00219_),
    .RESET_B(net610),
    .Q(\addroundkey_data_o[66] ));
 sky130_fd_sc_hd__dfrtp_4 _16776_ (.CLK(clknet_leaf_48_clk),
    .D(_00220_),
    .RESET_B(net610),
    .Q(\addroundkey_data_o[67] ));
 sky130_fd_sc_hd__dfrtp_4 _16777_ (.CLK(clknet_leaf_48_clk),
    .D(_00221_),
    .RESET_B(net611),
    .Q(\addroundkey_data_o[68] ));
 sky130_fd_sc_hd__dfrtp_4 _16778_ (.CLK(clknet_leaf_79_clk),
    .D(_00222_),
    .RESET_B(net579),
    .Q(\addroundkey_data_o[69] ));
 sky130_fd_sc_hd__dfrtp_4 _16779_ (.CLK(clknet_leaf_79_clk),
    .D(_00223_),
    .RESET_B(net579),
    .Q(\addroundkey_data_o[70] ));
 sky130_fd_sc_hd__dfrtp_4 _16780_ (.CLK(clknet_leaf_79_clk),
    .D(_00224_),
    .RESET_B(net579),
    .Q(\addroundkey_data_o[71] ));
 sky130_fd_sc_hd__dfrtp_4 _16781_ (.CLK(clknet_leaf_77_clk),
    .D(_00225_),
    .RESET_B(net590),
    .Q(\addroundkey_data_o[72] ));
 sky130_fd_sc_hd__dfrtp_4 _16782_ (.CLK(clknet_leaf_73_clk),
    .D(_00226_),
    .RESET_B(net593),
    .Q(\addroundkey_data_o[73] ));
 sky130_fd_sc_hd__dfrtp_1 _16783_ (.CLK(clknet_leaf_74_clk),
    .D(_00227_),
    .RESET_B(net591),
    .Q(\addroundkey_data_o[74] ));
 sky130_fd_sc_hd__dfrtp_4 _16784_ (.CLK(clknet_leaf_73_clk),
    .D(_00228_),
    .RESET_B(net593),
    .Q(\addroundkey_data_o[75] ));
 sky130_fd_sc_hd__dfrtp_4 _16785_ (.CLK(clknet_leaf_80_clk),
    .D(_00229_),
    .RESET_B(net578),
    .Q(\addroundkey_data_o[76] ));
 sky130_fd_sc_hd__dfrtp_4 _16786_ (.CLK(clknet_leaf_73_clk),
    .D(_00230_),
    .RESET_B(net590),
    .Q(\addroundkey_data_o[77] ));
 sky130_fd_sc_hd__dfrtp_4 _16787_ (.CLK(clknet_leaf_80_clk),
    .D(_00231_),
    .RESET_B(net579),
    .Q(\addroundkey_data_o[78] ));
 sky130_fd_sc_hd__dfrtp_4 _16788_ (.CLK(clknet_3_1__leaf_clk),
    .D(_00232_),
    .RESET_B(net594),
    .Q(\addroundkey_data_o[79] ));
 sky130_fd_sc_hd__dfrtp_2 _16789_ (.CLK(clknet_leaf_36_clk),
    .D(_00233_),
    .RESET_B(net649),
    .Q(\addroundkey_data_o[80] ));
 sky130_fd_sc_hd__dfrtp_4 _16790_ (.CLK(clknet_leaf_26_clk),
    .D(_00234_),
    .RESET_B(net649),
    .Q(\addroundkey_data_o[81] ));
 sky130_fd_sc_hd__dfrtp_4 _16791_ (.CLK(clknet_leaf_24_clk),
    .D(_00235_),
    .RESET_B(net649),
    .Q(\addroundkey_data_o[82] ));
 sky130_fd_sc_hd__dfrtp_4 _16792_ (.CLK(clknet_leaf_26_clk),
    .D(_00236_),
    .RESET_B(net649),
    .Q(\addroundkey_data_o[83] ));
 sky130_fd_sc_hd__dfrtp_4 _16793_ (.CLK(clknet_leaf_73_clk),
    .D(_00237_),
    .RESET_B(net593),
    .Q(\addroundkey_data_o[84] ));
 sky130_fd_sc_hd__dfrtp_4 _16794_ (.CLK(clknet_leaf_39_clk),
    .D(_00238_),
    .RESET_B(net663),
    .Q(\addroundkey_data_o[85] ));
 sky130_fd_sc_hd__dfrtp_4 _16795_ (.CLK(clknet_leaf_73_clk),
    .D(_00239_),
    .RESET_B(net590),
    .Q(\addroundkey_data_o[86] ));
 sky130_fd_sc_hd__dfrtp_1 _16796_ (.CLK(clknet_leaf_26_clk),
    .D(_00240_),
    .RESET_B(net649),
    .Q(\addroundkey_data_o[87] ));
 sky130_fd_sc_hd__dfrtp_2 _16797_ (.CLK(clknet_leaf_73_clk),
    .D(_00241_),
    .RESET_B(net593),
    .Q(\addroundkey_data_o[88] ));
 sky130_fd_sc_hd__dfrtp_4 _16798_ (.CLK(clknet_leaf_79_clk),
    .D(_00242_),
    .RESET_B(net579),
    .Q(\addroundkey_data_o[89] ));
 sky130_fd_sc_hd__dfrtp_4 _16799_ (.CLK(clknet_leaf_63_clk),
    .D(_00243_),
    .RESET_B(net598),
    .Q(\addroundkey_data_o[90] ));
 sky130_fd_sc_hd__dfrtp_4 _16800_ (.CLK(clknet_leaf_63_clk),
    .D(_00244_),
    .RESET_B(net598),
    .Q(\addroundkey_data_o[91] ));
 sky130_fd_sc_hd__dfrtp_2 _16801_ (.CLK(clknet_leaf_69_clk),
    .D(_00245_),
    .RESET_B(net593),
    .Q(\addroundkey_data_o[92] ));
 sky130_fd_sc_hd__dfrtp_4 _16802_ (.CLK(clknet_leaf_79_clk),
    .D(_00246_),
    .RESET_B(net579),
    .Q(\addroundkey_data_o[93] ));
 sky130_fd_sc_hd__dfrtp_2 _16803_ (.CLK(clknet_leaf_73_clk),
    .D(_00247_),
    .RESET_B(net593),
    .Q(\addroundkey_data_o[94] ));
 sky130_fd_sc_hd__dfrtp_4 _16804_ (.CLK(clknet_leaf_79_clk),
    .D(_00248_),
    .RESET_B(net578),
    .Q(\addroundkey_data_o[95] ));
 sky130_fd_sc_hd__dfrtp_4 _16805_ (.CLK(clknet_leaf_80_clk),
    .D(_00249_),
    .RESET_B(net578),
    .Q(\addroundkey_data_o[96] ));
 sky130_fd_sc_hd__dfrtp_4 _16806_ (.CLK(clknet_leaf_80_clk),
    .D(_00250_),
    .RESET_B(net578),
    .Q(\addroundkey_data_o[97] ));
 sky130_fd_sc_hd__dfrtp_4 _16807_ (.CLK(clknet_leaf_74_clk),
    .D(_00251_),
    .RESET_B(net591),
    .Q(\addroundkey_data_o[98] ));
 sky130_fd_sc_hd__dfrtp_4 _16808_ (.CLK(clknet_leaf_4_clk),
    .D(_00252_),
    .RESET_B(net591),
    .Q(\addroundkey_data_o[99] ));
 sky130_fd_sc_hd__dfrtp_4 _16809_ (.CLK(clknet_leaf_81_clk),
    .D(_00253_),
    .RESET_B(net586),
    .Q(\addroundkey_data_o[100] ));
 sky130_fd_sc_hd__dfrtp_4 _16810_ (.CLK(clknet_leaf_81_clk),
    .D(_00254_),
    .RESET_B(net586),
    .Q(\addroundkey_data_o[101] ));
 sky130_fd_sc_hd__dfrtp_4 _16811_ (.CLK(clknet_leaf_74_clk),
    .D(_00255_),
    .RESET_B(net591),
    .Q(\addroundkey_data_o[102] ));
 sky130_fd_sc_hd__dfrtp_4 _16812_ (.CLK(clknet_leaf_75_clk),
    .D(_00256_),
    .RESET_B(net586),
    .Q(\addroundkey_data_o[103] ));
 sky130_fd_sc_hd__dfrtp_2 _16813_ (.CLK(clknet_leaf_74_clk),
    .D(_00257_),
    .RESET_B(net591),
    .Q(\addroundkey_data_o[104] ));
 sky130_fd_sc_hd__dfrtp_4 _16814_ (.CLK(clknet_leaf_74_clk),
    .D(_00258_),
    .RESET_B(net591),
    .Q(\addroundkey_data_o[105] ));
 sky130_fd_sc_hd__dfrtp_4 _16815_ (.CLK(clknet_leaf_4_clk),
    .D(_00259_),
    .RESET_B(net584),
    .Q(\addroundkey_data_o[106] ));
 sky130_fd_sc_hd__dfrtp_4 _16816_ (.CLK(clknet_leaf_82_clk),
    .D(_00260_),
    .RESET_B(net585),
    .Q(\addroundkey_data_o[107] ));
 sky130_fd_sc_hd__dfrtp_4 _16817_ (.CLK(clknet_leaf_82_clk),
    .D(_00261_),
    .RESET_B(net585),
    .Q(\addroundkey_data_o[108] ));
 sky130_fd_sc_hd__dfrtp_4 _16818_ (.CLK(clknet_leaf_4_clk),
    .D(_00262_),
    .RESET_B(net591),
    .Q(\addroundkey_data_o[109] ));
 sky130_fd_sc_hd__dfrtp_4 _16819_ (.CLK(clknet_leaf_4_clk),
    .D(_00263_),
    .RESET_B(net591),
    .Q(\addroundkey_data_o[110] ));
 sky130_fd_sc_hd__dfrtp_2 _16820_ (.CLK(clknet_leaf_4_clk),
    .D(_00264_),
    .RESET_B(net584),
    .Q(\addroundkey_data_o[111] ));
 sky130_fd_sc_hd__dfrtp_4 _16821_ (.CLK(clknet_leaf_81_clk),
    .D(_00265_),
    .RESET_B(net586),
    .Q(\addroundkey_data_o[112] ));
 sky130_fd_sc_hd__dfrtp_4 _16822_ (.CLK(clknet_leaf_75_clk),
    .D(_00266_),
    .RESET_B(net587),
    .Q(\addroundkey_data_o[113] ));
 sky130_fd_sc_hd__dfrtp_1 _16823_ (.CLK(clknet_leaf_8_clk),
    .D(_00267_),
    .RESET_B(net633),
    .Q(\addroundkey_data_o[114] ));
 sky130_fd_sc_hd__dfrtp_1 _16824_ (.CLK(clknet_leaf_29_clk),
    .D(_00268_),
    .RESET_B(net635),
    .Q(\addroundkey_data_o[115] ));
 sky130_fd_sc_hd__dfrtp_2 _16825_ (.CLK(clknet_leaf_8_clk),
    .D(_00269_),
    .RESET_B(net632),
    .Q(\addroundkey_data_o[116] ));
 sky130_fd_sc_hd__dfrtp_4 _16826_ (.CLK(clknet_leaf_76_clk),
    .D(_00270_),
    .RESET_B(net586),
    .Q(\addroundkey_data_o[117] ));
 sky130_fd_sc_hd__dfrtp_1 _16827_ (.CLK(clknet_leaf_8_clk),
    .D(_00271_),
    .RESET_B(net633),
    .Q(\addroundkey_data_o[118] ));
 sky130_fd_sc_hd__dfrtp_4 _16828_ (.CLK(clknet_leaf_73_clk),
    .D(_00272_),
    .RESET_B(net590),
    .Q(\addroundkey_data_o[119] ));
 sky130_fd_sc_hd__dfrtp_1 _16829_ (.CLK(clknet_leaf_74_clk),
    .D(_00273_),
    .RESET_B(net591),
    .Q(\addroundkey_data_o[120] ));
 sky130_fd_sc_hd__dfrtp_4 _16830_ (.CLK(clknet_leaf_73_clk),
    .D(_00274_),
    .RESET_B(net593),
    .Q(\addroundkey_data_o[121] ));
 sky130_fd_sc_hd__dfrtp_4 _16831_ (.CLK(clknet_leaf_74_clk),
    .D(_00275_),
    .RESET_B(net587),
    .Q(\addroundkey_data_o[122] ));
 sky130_fd_sc_hd__dfrtp_4 _16832_ (.CLK(clknet_leaf_69_clk),
    .D(_00276_),
    .RESET_B(net604),
    .Q(\addroundkey_data_o[123] ));
 sky130_fd_sc_hd__dfrtp_2 _16833_ (.CLK(clknet_leaf_47_clk),
    .D(_00277_),
    .RESET_B(net612),
    .Q(\addroundkey_data_o[124] ));
 sky130_fd_sc_hd__dfrtp_2 _16834_ (.CLK(clknet_leaf_47_clk),
    .D(_00278_),
    .RESET_B(net651),
    .Q(\addroundkey_data_o[125] ));
 sky130_fd_sc_hd__dfrtp_4 _16835_ (.CLK(clknet_leaf_68_clk),
    .D(_00279_),
    .RESET_B(net608),
    .Q(\addroundkey_data_o[126] ));
 sky130_fd_sc_hd__dfrtp_2 _16836_ (.CLK(clknet_leaf_69_clk),
    .D(_00280_),
    .RESET_B(net608),
    .Q(\addroundkey_data_o[127] ));
 sky130_fd_sc_hd__dfrtp_1 _16837_ (.CLK(clknet_leaf_44_clk),
    .D(next_first_round_reg),
    .RESET_B(net663),
    .Q(first_round_reg));
 sky130_fd_sc_hd__dfxtp_1 _16838_ (.CLK(net421),
    .D(_00281_),
    .Q(\fifo_bank_register.bank[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16839_ (.CLK(net439),
    .D(_00282_),
    .Q(\fifo_bank_register.bank[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16840_ (.CLK(net420),
    .D(_00283_),
    .Q(\fifo_bank_register.bank[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16841_ (.CLK(net420),
    .D(_00284_),
    .Q(\fifo_bank_register.bank[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16842_ (.CLK(net420),
    .D(_00285_),
    .Q(\fifo_bank_register.bank[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16843_ (.CLK(net421),
    .D(_00286_),
    .Q(\fifo_bank_register.bank[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16844_ (.CLK(net425),
    .D(_00287_),
    .Q(\fifo_bank_register.bank[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16845_ (.CLK(net425),
    .D(_00288_),
    .Q(\fifo_bank_register.bank[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16846_ (.CLK(net425),
    .D(_00289_),
    .Q(\fifo_bank_register.bank[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16847_ (.CLK(net426),
    .D(_00290_),
    .Q(\fifo_bank_register.bank[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16848_ (.CLK(net503),
    .D(_00291_),
    .Q(\fifo_bank_register.bank[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16849_ (.CLK(net533),
    .D(_00292_),
    .Q(\fifo_bank_register.bank[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16850_ (.CLK(net504),
    .D(_00293_),
    .Q(\fifo_bank_register.bank[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16851_ (.CLK(net517),
    .D(_00294_),
    .Q(\fifo_bank_register.bank[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16852_ (.CLK(net534),
    .D(_00295_),
    .Q(\fifo_bank_register.bank[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16853_ (.CLK(net505),
    .D(_00296_),
    .Q(\fifo_bank_register.bank[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16854_ (.CLK(net497),
    .D(_00297_),
    .Q(\fifo_bank_register.bank[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _16855_ (.CLK(net532),
    .D(_00298_),
    .Q(\fifo_bank_register.bank[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _16856_ (.CLK(net532),
    .D(_00299_),
    .Q(\fifo_bank_register.bank[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _16857_ (.CLK(net505),
    .D(_00300_),
    .Q(\fifo_bank_register.bank[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _16858_ (.CLK(net501),
    .D(_00301_),
    .Q(\fifo_bank_register.bank[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _16859_ (.CLK(net484),
    .D(_00302_),
    .Q(\fifo_bank_register.bank[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _16860_ (.CLK(net501),
    .D(_00303_),
    .Q(\fifo_bank_register.bank[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _16861_ (.CLK(net483),
    .D(_00304_),
    .Q(\fifo_bank_register.bank[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _16862_ (.CLK(net482),
    .D(_00305_),
    .Q(\fifo_bank_register.bank[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _16863_ (.CLK(net488),
    .D(_00306_),
    .Q(\fifo_bank_register.bank[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _16864_ (.CLK(net483),
    .D(_00307_),
    .Q(\fifo_bank_register.bank[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _16865_ (.CLK(net479),
    .D(_00308_),
    .Q(\fifo_bank_register.bank[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _16866_ (.CLK(net486),
    .D(_00309_),
    .Q(\fifo_bank_register.bank[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _16867_ (.CLK(net499),
    .D(_00310_),
    .Q(\fifo_bank_register.bank[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _16868_ (.CLK(net430),
    .D(_00311_),
    .Q(\fifo_bank_register.bank[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _16869_ (.CLK(net437),
    .D(_00312_),
    .Q(\fifo_bank_register.bank[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _16870_ (.CLK(net417),
    .D(_00313_),
    .Q(\fifo_bank_register.bank[8][32] ));
 sky130_fd_sc_hd__dfxtp_1 _16871_ (.CLK(net423),
    .D(_00314_),
    .Q(\fifo_bank_register.bank[8][33] ));
 sky130_fd_sc_hd__dfxtp_1 _16872_ (.CLK(net430),
    .D(_00315_),
    .Q(\fifo_bank_register.bank[8][34] ));
 sky130_fd_sc_hd__dfxtp_1 _16873_ (.CLK(net428),
    .D(_00316_),
    .Q(\fifo_bank_register.bank[8][35] ));
 sky130_fd_sc_hd__dfxtp_1 _16874_ (.CLK(net423),
    .D(_00317_),
    .Q(\fifo_bank_register.bank[8][36] ));
 sky130_fd_sc_hd__dfxtp_1 _16875_ (.CLK(net417),
    .D(_00318_),
    .Q(\fifo_bank_register.bank[8][37] ));
 sky130_fd_sc_hd__dfxtp_1 _16876_ (.CLK(net416),
    .D(_00319_),
    .Q(\fifo_bank_register.bank[8][38] ));
 sky130_fd_sc_hd__dfxtp_1 _16877_ (.CLK(net415),
    .D(_00320_),
    .Q(\fifo_bank_register.bank[8][39] ));
 sky130_fd_sc_hd__dfxtp_1 _16878_ (.CLK(net393),
    .D(_00321_),
    .Q(\fifo_bank_register.bank[8][40] ));
 sky130_fd_sc_hd__dfxtp_1 _16879_ (.CLK(net398),
    .D(_00322_),
    .Q(\fifo_bank_register.bank[8][41] ));
 sky130_fd_sc_hd__dfxtp_1 _16880_ (.CLK(net405),
    .D(_00323_),
    .Q(\fifo_bank_register.bank[8][42] ));
 sky130_fd_sc_hd__dfxtp_1 _16881_ (.CLK(net393),
    .D(_00324_),
    .Q(\fifo_bank_register.bank[8][43] ));
 sky130_fd_sc_hd__dfxtp_1 _16882_ (.CLK(net389),
    .D(_00325_),
    .Q(\fifo_bank_register.bank[8][44] ));
 sky130_fd_sc_hd__dfxtp_1 _16883_ (.CLK(net405),
    .D(_00326_),
    .Q(\fifo_bank_register.bank[8][45] ));
 sky130_fd_sc_hd__dfxtp_1 _16884_ (.CLK(net394),
    .D(_00327_),
    .Q(\fifo_bank_register.bank[8][46] ));
 sky130_fd_sc_hd__dfxtp_1 _16885_ (.CLK(net394),
    .D(_00328_),
    .Q(\fifo_bank_register.bank[8][47] ));
 sky130_fd_sc_hd__dfxtp_1 _16886_ (.CLK(net393),
    .D(_00329_),
    .Q(\fifo_bank_register.bank[8][48] ));
 sky130_fd_sc_hd__dfxtp_1 _16887_ (.CLK(net405),
    .D(_00330_),
    .Q(\fifo_bank_register.bank[8][49] ));
 sky130_fd_sc_hd__dfxtp_1 _16888_ (.CLK(net558),
    .D(_00331_),
    .Q(\fifo_bank_register.bank[8][50] ));
 sky130_fd_sc_hd__dfxtp_1 _16889_ (.CLK(net572),
    .D(_00332_),
    .Q(\fifo_bank_register.bank[8][51] ));
 sky130_fd_sc_hd__dfxtp_1 _16890_ (.CLK(net562),
    .D(_00333_),
    .Q(\fifo_bank_register.bank[8][52] ));
 sky130_fd_sc_hd__dfxtp_1 _16891_ (.CLK(net563),
    .D(_00334_),
    .Q(\fifo_bank_register.bank[8][53] ));
 sky130_fd_sc_hd__dfxtp_1 _16892_ (.CLK(net570),
    .D(_00335_),
    .Q(\fifo_bank_register.bank[8][54] ));
 sky130_fd_sc_hd__dfxtp_1 _16893_ (.CLK(net571),
    .D(_00336_),
    .Q(\fifo_bank_register.bank[8][55] ));
 sky130_fd_sc_hd__dfxtp_1 _16894_ (.CLK(net571),
    .D(_00337_),
    .Q(\fifo_bank_register.bank[8][56] ));
 sky130_fd_sc_hd__dfxtp_1 _16895_ (.CLK(net550),
    .D(_00338_),
    .Q(\fifo_bank_register.bank[8][57] ));
 sky130_fd_sc_hd__dfxtp_1 _16896_ (.CLK(net558),
    .D(_00339_),
    .Q(\fifo_bank_register.bank[8][58] ));
 sky130_fd_sc_hd__dfxtp_1 _16897_ (.CLK(net572),
    .D(_00340_),
    .Q(\fifo_bank_register.bank[8][59] ));
 sky130_fd_sc_hd__dfxtp_1 _16898_ (.CLK(net514),
    .D(_00341_),
    .Q(\fifo_bank_register.bank[8][60] ));
 sky130_fd_sc_hd__dfxtp_1 _16899_ (.CLK(net527),
    .D(_00342_),
    .Q(\fifo_bank_register.bank[8][61] ));
 sky130_fd_sc_hd__dfxtp_1 _16900_ (.CLK(net511),
    .D(_00343_),
    .Q(\fifo_bank_register.bank[8][62] ));
 sky130_fd_sc_hd__dfxtp_1 _16901_ (.CLK(net524),
    .D(_00344_),
    .Q(\fifo_bank_register.bank[8][63] ));
 sky130_fd_sc_hd__dfxtp_1 _16902_ (.CLK(net509),
    .D(_00345_),
    .Q(\fifo_bank_register.bank[8][64] ));
 sky130_fd_sc_hd__dfxtp_1 _16903_ (.CLK(net518),
    .D(_00346_),
    .Q(\fifo_bank_register.bank[8][65] ));
 sky130_fd_sc_hd__dfxtp_1 _16904_ (.CLK(net526),
    .D(_00347_),
    .Q(\fifo_bank_register.bank[8][66] ));
 sky130_fd_sc_hd__dfxtp_1 _16905_ (.CLK(net509),
    .D(_00348_),
    .Q(\fifo_bank_register.bank[8][67] ));
 sky130_fd_sc_hd__dfxtp_1 _16906_ (.CLK(net511),
    .D(_00349_),
    .Q(\fifo_bank_register.bank[8][68] ));
 sky130_fd_sc_hd__dfxtp_1 _16907_ (.CLK(net518),
    .D(_00350_),
    .Q(\fifo_bank_register.bank[8][69] ));
 sky130_fd_sc_hd__dfxtp_1 _16908_ (.CLK(net519),
    .D(_00351_),
    .Q(\fifo_bank_register.bank[8][70] ));
 sky130_fd_sc_hd__dfxtp_1 _16909_ (.CLK(net525),
    .D(_00352_),
    .Q(\fifo_bank_register.bank[8][71] ));
 sky130_fd_sc_hd__dfxtp_1 _16910_ (.CLK(net555),
    .D(_00353_),
    .Q(\fifo_bank_register.bank[8][72] ));
 sky130_fd_sc_hd__dfxtp_1 _16911_ (.CLK(net552),
    .D(_00354_),
    .Q(\fifo_bank_register.bank[8][73] ));
 sky130_fd_sc_hd__dfxtp_1 _16912_ (.CLK(net545),
    .D(_00355_),
    .Q(\fifo_bank_register.bank[8][74] ));
 sky130_fd_sc_hd__dfxtp_1 _16913_ (.CLK(net545),
    .D(_00356_),
    .Q(\fifo_bank_register.bank[8][75] ));
 sky130_fd_sc_hd__dfxtp_1 _16914_ (.CLK(net545),
    .D(_00357_),
    .Q(\fifo_bank_register.bank[8][76] ));
 sky130_fd_sc_hd__dfxtp_1 _16915_ (.CLK(net553),
    .D(_00358_),
    .Q(\fifo_bank_register.bank[8][77] ));
 sky130_fd_sc_hd__dfxtp_1 _16916_ (.CLK(net525),
    .D(_00359_),
    .Q(\fifo_bank_register.bank[8][78] ));
 sky130_fd_sc_hd__dfxtp_1 _16917_ (.CLK(net549),
    .D(_00360_),
    .Q(\fifo_bank_register.bank[8][79] ));
 sky130_fd_sc_hd__dfxtp_1 _16918_ (.CLK(net566),
    .D(_00361_),
    .Q(\fifo_bank_register.bank[8][80] ));
 sky130_fd_sc_hd__dfxtp_1 _16919_ (.CLK(net565),
    .D(_00362_),
    .Q(\fifo_bank_register.bank[8][81] ));
 sky130_fd_sc_hd__dfxtp_1 _16920_ (.CLK(net560),
    .D(_00363_),
    .Q(\fifo_bank_register.bank[8][82] ));
 sky130_fd_sc_hd__dfxtp_1 _16921_ (.CLK(net561),
    .D(_00364_),
    .Q(\fifo_bank_register.bank[8][83] ));
 sky130_fd_sc_hd__dfxtp_1 _16922_ (.CLK(net548),
    .D(_00365_),
    .Q(\fifo_bank_register.bank[8][84] ));
 sky130_fd_sc_hd__dfxtp_1 _16923_ (.CLK(net566),
    .D(_00366_),
    .Q(\fifo_bank_register.bank[8][85] ));
 sky130_fd_sc_hd__dfxtp_1 _16924_ (.CLK(net547),
    .D(_00367_),
    .Q(\fifo_bank_register.bank[8][86] ));
 sky130_fd_sc_hd__dfxtp_1 _16925_ (.CLK(net561),
    .D(_00368_),
    .Q(\fifo_bank_register.bank[8][87] ));
 sky130_fd_sc_hd__dfxtp_1 _16926_ (.CLK(net566),
    .D(_00369_),
    .Q(\fifo_bank_register.bank[8][88] ));
 sky130_fd_sc_hd__dfxtp_1 _16927_ (.CLK(net548),
    .D(_00370_),
    .Q(\fifo_bank_register.bank[8][89] ));
 sky130_fd_sc_hd__dfxtp_1 _16928_ (.CLK(net409),
    .D(_00371_),
    .Q(\fifo_bank_register.bank[8][90] ));
 sky130_fd_sc_hd__dfxtp_1 _16929_ (.CLK(net401),
    .D(_00372_),
    .Q(\fifo_bank_register.bank[8][91] ));
 sky130_fd_sc_hd__dfxtp_1 _16930_ (.CLK(net410),
    .D(_00373_),
    .Q(\fifo_bank_register.bank[8][92] ));
 sky130_fd_sc_hd__dfxtp_1 _16931_ (.CLK(net400),
    .D(_00374_),
    .Q(\fifo_bank_register.bank[8][93] ));
 sky130_fd_sc_hd__dfxtp_1 _16932_ (.CLK(net454),
    .D(_00375_),
    .Q(\fifo_bank_register.bank[8][94] ));
 sky130_fd_sc_hd__dfxtp_1 _16933_ (.CLK(net402),
    .D(_00376_),
    .Q(\fifo_bank_register.bank[8][95] ));
 sky130_fd_sc_hd__dfxtp_1 _16934_ (.CLK(net445),
    .D(_00377_),
    .Q(\fifo_bank_register.bank[8][96] ));
 sky130_fd_sc_hd__dfxtp_1 _16935_ (.CLK(net454),
    .D(_00378_),
    .Q(\fifo_bank_register.bank[8][97] ));
 sky130_fd_sc_hd__dfxtp_1 _16936_ (.CLK(net448),
    .D(_00379_),
    .Q(\fifo_bank_register.bank[8][98] ));
 sky130_fd_sc_hd__dfxtp_1 _16937_ (.CLK(net445),
    .D(_00380_),
    .Q(\fifo_bank_register.bank[8][99] ));
 sky130_fd_sc_hd__dfxtp_1 _16938_ (.CLK(net452),
    .D(_00381_),
    .Q(\fifo_bank_register.bank[8][100] ));
 sky130_fd_sc_hd__dfxtp_1 _16939_ (.CLK(net450),
    .D(_00382_),
    .Q(\fifo_bank_register.bank[8][101] ));
 sky130_fd_sc_hd__dfxtp_1 _16940_ (.CLK(net465),
    .D(_00383_),
    .Q(\fifo_bank_register.bank[8][102] ));
 sky130_fd_sc_hd__dfxtp_1 _16941_ (.CLK(net467),
    .D(_00384_),
    .Q(\fifo_bank_register.bank[8][103] ));
 sky130_fd_sc_hd__dfxtp_1 _16942_ (.CLK(net463),
    .D(_00385_),
    .Q(\fifo_bank_register.bank[8][104] ));
 sky130_fd_sc_hd__dfxtp_1 _16943_ (.CLK(net468),
    .D(_00386_),
    .Q(\fifo_bank_register.bank[8][105] ));
 sky130_fd_sc_hd__dfxtp_1 _16944_ (.CLK(net463),
    .D(_00387_),
    .Q(\fifo_bank_register.bank[8][106] ));
 sky130_fd_sc_hd__dfxtp_1 _16945_ (.CLK(net451),
    .D(_00388_),
    .Q(\fifo_bank_register.bank[8][107] ));
 sky130_fd_sc_hd__dfxtp_1 _16946_ (.CLK(net452),
    .D(_00389_),
    .Q(\fifo_bank_register.bank[8][108] ));
 sky130_fd_sc_hd__dfxtp_1 _16947_ (.CLK(net459),
    .D(_00390_),
    .Q(\fifo_bank_register.bank[8][109] ));
 sky130_fd_sc_hd__dfxtp_1 _16948_ (.CLK(net432),
    .D(_00391_),
    .Q(\fifo_bank_register.bank[8][110] ));
 sky130_fd_sc_hd__dfxtp_1 _16949_ (.CLK(net411),
    .D(_00392_),
    .Q(\fifo_bank_register.bank[8][111] ));
 sky130_fd_sc_hd__dfxtp_1 _16950_ (.CLK(net411),
    .D(_00393_),
    .Q(\fifo_bank_register.bank[8][112] ));
 sky130_fd_sc_hd__dfxtp_1 _16951_ (.CLK(net470),
    .D(_00394_),
    .Q(\fifo_bank_register.bank[8][113] ));
 sky130_fd_sc_hd__dfxtp_1 _16952_ (.CLK(net456),
    .D(_00395_),
    .Q(\fifo_bank_register.bank[8][114] ));
 sky130_fd_sc_hd__dfxtp_1 _16953_ (.CLK(net469),
    .D(_00396_),
    .Q(\fifo_bank_register.bank[8][115] ));
 sky130_fd_sc_hd__dfxtp_1 _16954_ (.CLK(net456),
    .D(_00397_),
    .Q(\fifo_bank_register.bank[8][116] ));
 sky130_fd_sc_hd__dfxtp_1 _16955_ (.CLK(net432),
    .D(_00398_),
    .Q(\fifo_bank_register.bank[8][117] ));
 sky130_fd_sc_hd__dfxtp_1 _16956_ (.CLK(net457),
    .D(_00399_),
    .Q(\fifo_bank_register.bank[8][118] ));
 sky130_fd_sc_hd__dfxtp_1 _16957_ (.CLK(net469),
    .D(_00400_),
    .Q(\fifo_bank_register.bank[8][119] ));
 sky130_fd_sc_hd__dfxtp_1 _16958_ (.CLK(net442),
    .D(_00401_),
    .Q(\fifo_bank_register.bank[8][120] ));
 sky130_fd_sc_hd__dfxtp_1 _16959_ (.CLK(net490),
    .D(_00402_),
    .Q(\fifo_bank_register.bank[8][121] ));
 sky130_fd_sc_hd__dfxtp_1 _16960_ (.CLK(net491),
    .D(_00403_),
    .Q(\fifo_bank_register.bank[8][122] ));
 sky130_fd_sc_hd__dfxtp_1 _16961_ (.CLK(net437),
    .D(_00404_),
    .Q(\fifo_bank_register.bank[8][123] ));
 sky130_fd_sc_hd__dfxtp_1 _16962_ (.CLK(net471),
    .D(_00405_),
    .Q(\fifo_bank_register.bank[8][124] ));
 sky130_fd_sc_hd__dfxtp_1 _16963_ (.CLK(net495),
    .D(_00406_),
    .Q(\fifo_bank_register.bank[8][125] ));
 sky130_fd_sc_hd__dfxtp_1 _16964_ (.CLK(net531),
    .D(_00407_),
    .Q(\fifo_bank_register.bank[8][126] ));
 sky130_fd_sc_hd__dfxtp_1 _16965_ (.CLK(net471),
    .D(_00408_),
    .Q(\fifo_bank_register.bank[8][127] ));
 sky130_fd_sc_hd__dfxtp_1 _16966_ (.CLK(net475),
    .D(_00409_),
    .Q(\fifo_bank_register.bank[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _16967_ (.CLK(net492),
    .D(_00410_),
    .Q(\fifo_bank_register.bank[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _16968_ (.CLK(net476),
    .D(_00411_),
    .Q(\fifo_bank_register.bank[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _16969_ (.CLK(net475),
    .D(_00412_),
    .Q(\fifo_bank_register.bank[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _16970_ (.CLK(net476),
    .D(_00413_),
    .Q(\fifo_bank_register.bank[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _16971_ (.CLK(net476),
    .D(_00414_),
    .Q(\fifo_bank_register.bank[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _16972_ (.CLK(net479),
    .D(_00415_),
    .Q(\fifo_bank_register.bank[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _16973_ (.CLK(net479),
    .D(_00416_),
    .Q(\fifo_bank_register.bank[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _16974_ (.CLK(net480),
    .D(_00417_),
    .Q(\fifo_bank_register.bank[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _16975_ (.CLK(net480),
    .D(_00418_),
    .Q(\fifo_bank_register.bank[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _16976_ (.CLK(net500),
    .D(_00419_),
    .Q(\fifo_bank_register.bank[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _16977_ (.CLK(net503),
    .D(_00420_),
    .Q(\fifo_bank_register.bank[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _16978_ (.CLK(net500),
    .D(_00421_),
    .Q(\fifo_bank_register.bank[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _16979_ (.CLK(net506),
    .D(_00422_),
    .Q(\fifo_bank_register.bank[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _16980_ (.CLK(net506),
    .D(_00423_),
    .Q(\fifo_bank_register.bank[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _16981_ (.CLK(net505),
    .D(_00424_),
    .Q(\fifo_bank_register.bank[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _16982_ (.CLK(net496),
    .D(_00425_),
    .Q(\fifo_bank_register.bank[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _16983_ (.CLK(net497),
    .D(_00426_),
    .Q(\fifo_bank_register.bank[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _16984_ (.CLK(net503),
    .D(_00427_),
    .Q(\fifo_bank_register.bank[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _16985_ (.CLK(net502),
    .D(_00428_),
    .Q(\fifo_bank_register.bank[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _16986_ (.CLK(net508),
    .D(_00429_),
    .Q(\fifo_bank_register.bank[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _16987_ (.CLK(net483),
    .D(_00430_),
    .Q(\fifo_bank_register.bank[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _16988_ (.CLK(net501),
    .D(_00431_),
    .Q(\fifo_bank_register.bank[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _16989_ (.CLK(net487),
    .D(_00432_),
    .Q(\fifo_bank_register.bank[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _16990_ (.CLK(net482),
    .D(_00433_),
    .Q(\fifo_bank_register.bank[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _16991_ (.CLK(net508),
    .D(_00434_),
    .Q(\fifo_bank_register.bank[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _16992_ (.CLK(net508),
    .D(_00435_),
    .Q(\fifo_bank_register.bank[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _16993_ (.CLK(net486),
    .D(_00436_),
    .Q(\fifo_bank_register.bank[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _16994_ (.CLK(net486),
    .D(_00437_),
    .Q(\fifo_bank_register.bank[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _16995_ (.CLK(net499),
    .D(_00438_),
    .Q(\fifo_bank_register.bank[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _16996_ (.CLK(net424),
    .D(_00439_),
    .Q(\fifo_bank_register.bank[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _16997_ (.CLK(net423),
    .D(_00440_),
    .Q(\fifo_bank_register.bank[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _16998_ (.CLK(net414),
    .D(_00441_),
    .Q(\fifo_bank_register.bank[7][32] ));
 sky130_fd_sc_hd__dfxtp_1 _16999_ (.CLK(net424),
    .D(_00442_),
    .Q(\fifo_bank_register.bank[7][33] ));
 sky130_fd_sc_hd__dfxtp_1 _17000_ (.CLK(net417),
    .D(_00443_),
    .Q(\fifo_bank_register.bank[7][34] ));
 sky130_fd_sc_hd__dfxtp_1 _17001_ (.CLK(net416),
    .D(_00444_),
    .Q(\fifo_bank_register.bank[7][35] ));
 sky130_fd_sc_hd__dfxtp_1 _17002_ (.CLK(net422),
    .D(_00445_),
    .Q(\fifo_bank_register.bank[7][36] ));
 sky130_fd_sc_hd__dfxtp_1 _17003_ (.CLK(net414),
    .D(_00446_),
    .Q(\fifo_bank_register.bank[7][37] ));
 sky130_fd_sc_hd__dfxtp_1 _17004_ (.CLK(net418),
    .D(_00447_),
    .Q(\fifo_bank_register.bank[7][38] ));
 sky130_fd_sc_hd__dfxtp_1 _17005_ (.CLK(net414),
    .D(_00448_),
    .Q(\fifo_bank_register.bank[7][39] ));
 sky130_fd_sc_hd__dfxtp_1 _17006_ (.CLK(net392),
    .D(_00449_),
    .Q(\fifo_bank_register.bank[7][40] ));
 sky130_fd_sc_hd__dfxtp_1 _17007_ (.CLK(net389),
    .D(_00450_),
    .Q(\fifo_bank_register.bank[7][41] ));
 sky130_fd_sc_hd__dfxtp_1 _17008_ (.CLK(net394),
    .D(_00451_),
    .Q(\fifo_bank_register.bank[7][42] ));
 sky130_fd_sc_hd__dfxtp_1 _17009_ (.CLK(net392),
    .D(_00452_),
    .Q(\fifo_bank_register.bank[7][43] ));
 sky130_fd_sc_hd__dfxtp_1 _17010_ (.CLK(net392),
    .D(_00453_),
    .Q(\fifo_bank_register.bank[7][44] ));
 sky130_fd_sc_hd__dfxtp_1 _17011_ (.CLK(net405),
    .D(_00454_),
    .Q(\fifo_bank_register.bank[7][45] ));
 sky130_fd_sc_hd__dfxtp_1 _17012_ (.CLK(net392),
    .D(_00455_),
    .Q(\fifo_bank_register.bank[7][46] ));
 sky130_fd_sc_hd__dfxtp_1 _17013_ (.CLK(net396),
    .D(_00456_),
    .Q(\fifo_bank_register.bank[7][47] ));
 sky130_fd_sc_hd__dfxtp_1 _17014_ (.CLK(net397),
    .D(_00457_),
    .Q(\fifo_bank_register.bank[7][48] ));
 sky130_fd_sc_hd__dfxtp_1 _17015_ (.CLK(net407),
    .D(_00458_),
    .Q(\fifo_bank_register.bank[7][49] ));
 sky130_fd_sc_hd__dfxtp_1 _17016_ (.CLK(net558),
    .D(_00459_),
    .Q(\fifo_bank_register.bank[7][50] ));
 sky130_fd_sc_hd__dfxtp_1 _17017_ (.CLK(net573),
    .D(_00460_),
    .Q(\fifo_bank_register.bank[7][51] ));
 sky130_fd_sc_hd__dfxtp_1 _17018_ (.CLK(net563),
    .D(_00461_),
    .Q(\fifo_bank_register.bank[7][52] ));
 sky130_fd_sc_hd__dfxtp_1 _17019_ (.CLK(net562),
    .D(_00462_),
    .Q(\fifo_bank_register.bank[7][53] ));
 sky130_fd_sc_hd__dfxtp_1 _17020_ (.CLK(net556),
    .D(_00463_),
    .Q(\fifo_bank_register.bank[7][54] ));
 sky130_fd_sc_hd__dfxtp_1 _17021_ (.CLK(net570),
    .D(_00464_),
    .Q(\fifo_bank_register.bank[7][55] ));
 sky130_fd_sc_hd__dfxtp_1 _17022_ (.CLK(net571),
    .D(_00465_),
    .Q(\fifo_bank_register.bank[7][56] ));
 sky130_fd_sc_hd__dfxtp_1 _17023_ (.CLK(net550),
    .D(_00466_),
    .Q(\fifo_bank_register.bank[7][57] ));
 sky130_fd_sc_hd__dfxtp_1 _17024_ (.CLK(net557),
    .D(_00467_),
    .Q(\fifo_bank_register.bank[7][58] ));
 sky130_fd_sc_hd__dfxtp_1 _17025_ (.CLK(net572),
    .D(_00468_),
    .Q(\fifo_bank_register.bank[7][59] ));
 sky130_fd_sc_hd__dfxtp_1 _17026_ (.CLK(net515),
    .D(_00469_),
    .Q(\fifo_bank_register.bank[7][60] ));
 sky130_fd_sc_hd__dfxtp_1 _17027_ (.CLK(net525),
    .D(_00470_),
    .Q(\fifo_bank_register.bank[7][61] ));
 sky130_fd_sc_hd__dfxtp_1 _17028_ (.CLK(net523),
    .D(_00471_),
    .Q(\fifo_bank_register.bank[7][62] ));
 sky130_fd_sc_hd__dfxtp_1 _17029_ (.CLK(net524),
    .D(_00472_),
    .Q(\fifo_bank_register.bank[7][63] ));
 sky130_fd_sc_hd__dfxtp_1 _17030_ (.CLK(net514),
    .D(_00473_),
    .Q(\fifo_bank_register.bank[7][64] ));
 sky130_fd_sc_hd__dfxtp_1 _17031_ (.CLK(net526),
    .D(_00474_),
    .Q(\fifo_bank_register.bank[7][65] ));
 sky130_fd_sc_hd__dfxtp_1 _17032_ (.CLK(net526),
    .D(_00475_),
    .Q(\fifo_bank_register.bank[7][66] ));
 sky130_fd_sc_hd__dfxtp_1 _17033_ (.CLK(net515),
    .D(_00476_),
    .Q(\fifo_bank_register.bank[7][67] ));
 sky130_fd_sc_hd__dfxtp_1 _17034_ (.CLK(net521),
    .D(_00477_),
    .Q(\fifo_bank_register.bank[7][68] ));
 sky130_fd_sc_hd__dfxtp_1 _17035_ (.CLK(net516),
    .D(_00478_),
    .Q(\fifo_bank_register.bank[7][69] ));
 sky130_fd_sc_hd__dfxtp_1 _17036_ (.CLK(net518),
    .D(_00479_),
    .Q(\fifo_bank_register.bank[7][70] ));
 sky130_fd_sc_hd__dfxtp_1 _17037_ (.CLK(net519),
    .D(_00480_),
    .Q(\fifo_bank_register.bank[7][71] ));
 sky130_fd_sc_hd__dfxtp_1 _17038_ (.CLK(net546),
    .D(_00481_),
    .Q(\fifo_bank_register.bank[7][72] ));
 sky130_fd_sc_hd__dfxtp_1 _17039_ (.CLK(net545),
    .D(_00482_),
    .Q(\fifo_bank_register.bank[7][73] ));
 sky130_fd_sc_hd__dfxtp_1 _17040_ (.CLK(net546),
    .D(_00483_),
    .Q(\fifo_bank_register.bank[7][74] ));
 sky130_fd_sc_hd__dfxtp_1 _17041_ (.CLK(net543),
    .D(_00484_),
    .Q(\fifo_bank_register.bank[7][75] ));
 sky130_fd_sc_hd__dfxtp_1 _17042_ (.CLK(net545),
    .D(_00485_),
    .Q(\fifo_bank_register.bank[7][76] ));
 sky130_fd_sc_hd__dfxtp_1 _17043_ (.CLK(net546),
    .D(_00486_),
    .Q(\fifo_bank_register.bank[7][77] ));
 sky130_fd_sc_hd__dfxtp_1 _17044_ (.CLK(net516),
    .D(_00487_),
    .Q(\fifo_bank_register.bank[7][78] ));
 sky130_fd_sc_hd__dfxtp_1 _17045_ (.CLK(net547),
    .D(_00488_),
    .Q(\fifo_bank_register.bank[7][79] ));
 sky130_fd_sc_hd__dfxtp_1 _17046_ (.CLK(net541),
    .D(_00489_),
    .Q(\fifo_bank_register.bank[7][80] ));
 sky130_fd_sc_hd__dfxtp_1 _17047_ (.CLK(net540),
    .D(_00490_),
    .Q(\fifo_bank_register.bank[7][81] ));
 sky130_fd_sc_hd__dfxtp_1 _17048_ (.CLK(net538),
    .D(_00491_),
    .Q(\fifo_bank_register.bank[7][82] ));
 sky130_fd_sc_hd__dfxtp_1 _17049_ (.CLK(net539),
    .D(_00492_),
    .Q(\fifo_bank_register.bank[7][83] ));
 sky130_fd_sc_hd__dfxtp_1 _17050_ (.CLK(net536),
    .D(_00493_),
    .Q(\fifo_bank_register.bank[7][84] ));
 sky130_fd_sc_hd__dfxtp_1 _17051_ (.CLK(net540),
    .D(_00494_),
    .Q(\fifo_bank_register.bank[7][85] ));
 sky130_fd_sc_hd__dfxtp_1 _17052_ (.CLK(net536),
    .D(_00495_),
    .Q(\fifo_bank_register.bank[7][86] ));
 sky130_fd_sc_hd__dfxtp_1 _17053_ (.CLK(net538),
    .D(_00496_),
    .Q(\fifo_bank_register.bank[7][87] ));
 sky130_fd_sc_hd__dfxtp_1 _17054_ (.CLK(net541),
    .D(_00497_),
    .Q(\fifo_bank_register.bank[7][88] ));
 sky130_fd_sc_hd__dfxtp_1 _17055_ (.CLK(net536),
    .D(_00498_),
    .Q(\fifo_bank_register.bank[7][89] ));
 sky130_fd_sc_hd__dfxtp_1 _17056_ (.CLK(net409),
    .D(_00499_),
    .Q(\fifo_bank_register.bank[7][90] ));
 sky130_fd_sc_hd__dfxtp_1 _17057_ (.CLK(net401),
    .D(_00500_),
    .Q(\fifo_bank_register.bank[7][91] ));
 sky130_fd_sc_hd__dfxtp_1 _17058_ (.CLK(net410),
    .D(_00501_),
    .Q(\fifo_bank_register.bank[7][92] ));
 sky130_fd_sc_hd__dfxtp_1 _17059_ (.CLK(net400),
    .D(_00502_),
    .Q(\fifo_bank_register.bank[7][93] ));
 sky130_fd_sc_hd__dfxtp_1 _17060_ (.CLK(net447),
    .D(_00503_),
    .Q(\fifo_bank_register.bank[7][94] ));
 sky130_fd_sc_hd__dfxtp_1 _17061_ (.CLK(net400),
    .D(_00504_),
    .Q(\fifo_bank_register.bank[7][95] ));
 sky130_fd_sc_hd__dfxtp_1 _17062_ (.CLK(net401),
    .D(_00505_),
    .Q(\fifo_bank_register.bank[7][96] ));
 sky130_fd_sc_hd__dfxtp_1 _17063_ (.CLK(net402),
    .D(_00506_),
    .Q(\fifo_bank_register.bank[7][97] ));
 sky130_fd_sc_hd__dfxtp_1 _17064_ (.CLK(net446),
    .D(_00507_),
    .Q(\fifo_bank_register.bank[7][98] ));
 sky130_fd_sc_hd__dfxtp_1 _17065_ (.CLK(net446),
    .D(_00508_),
    .Q(\fifo_bank_register.bank[7][99] ));
 sky130_fd_sc_hd__dfxtp_1 _17066_ (.CLK(net447),
    .D(_00509_),
    .Q(\fifo_bank_register.bank[7][100] ));
 sky130_fd_sc_hd__dfxtp_1 _17067_ (.CLK(net446),
    .D(_00510_),
    .Q(\fifo_bank_register.bank[7][101] ));
 sky130_fd_sc_hd__dfxtp_1 _17068_ (.CLK(net464),
    .D(_00511_),
    .Q(\fifo_bank_register.bank[7][102] ));
 sky130_fd_sc_hd__dfxtp_1 _17069_ (.CLK(net458),
    .D(_00512_),
    .Q(\fifo_bank_register.bank[7][103] ));
 sky130_fd_sc_hd__dfxtp_1 _17070_ (.CLK(net462),
    .D(_00513_),
    .Q(\fifo_bank_register.bank[7][104] ));
 sky130_fd_sc_hd__dfxtp_1 _17071_ (.CLK(net467),
    .D(_00514_),
    .Q(\fifo_bank_register.bank[7][105] ));
 sky130_fd_sc_hd__dfxtp_1 _17072_ (.CLK(net464),
    .D(_00515_),
    .Q(\fifo_bank_register.bank[7][106] ));
 sky130_fd_sc_hd__dfxtp_1 _17073_ (.CLK(net462),
    .D(_00516_),
    .Q(\fifo_bank_register.bank[7][107] ));
 sky130_fd_sc_hd__dfxtp_1 _17074_ (.CLK(net452),
    .D(_00517_),
    .Q(\fifo_bank_register.bank[7][108] ));
 sky130_fd_sc_hd__dfxtp_1 _17075_ (.CLK(net455),
    .D(_00518_),
    .Q(\fifo_bank_register.bank[7][109] ));
 sky130_fd_sc_hd__dfxtp_1 _17076_ (.CLK(net434),
    .D(_00519_),
    .Q(\fifo_bank_register.bank[7][110] ));
 sky130_fd_sc_hd__dfxtp_1 _17077_ (.CLK(net412),
    .D(_00520_),
    .Q(\fifo_bank_register.bank[7][111] ));
 sky130_fd_sc_hd__dfxtp_1 _17078_ (.CLK(net432),
    .D(_00521_),
    .Q(\fifo_bank_register.bank[7][112] ));
 sky130_fd_sc_hd__dfxtp_1 _17079_ (.CLK(net428),
    .D(_00522_),
    .Q(\fifo_bank_register.bank[7][113] ));
 sky130_fd_sc_hd__dfxtp_1 _17080_ (.CLK(net407),
    .D(_00523_),
    .Q(\fifo_bank_register.bank[7][114] ));
 sky130_fd_sc_hd__dfxtp_1 _17081_ (.CLK(net434),
    .D(_00524_),
    .Q(\fifo_bank_register.bank[7][115] ));
 sky130_fd_sc_hd__dfxtp_1 _17082_ (.CLK(net412),
    .D(_00525_),
    .Q(\fifo_bank_register.bank[7][116] ));
 sky130_fd_sc_hd__dfxtp_1 _17083_ (.CLK(net434),
    .D(_00526_),
    .Q(\fifo_bank_register.bank[7][117] ));
 sky130_fd_sc_hd__dfxtp_1 _17084_ (.CLK(net412),
    .D(_00527_),
    .Q(\fifo_bank_register.bank[7][118] ));
 sky130_fd_sc_hd__dfxtp_1 _17085_ (.CLK(net430),
    .D(_00528_),
    .Q(\fifo_bank_register.bank[7][119] ));
 sky130_fd_sc_hd__dfxtp_1 _17086_ (.CLK(net441),
    .D(_00529_),
    .Q(\fifo_bank_register.bank[7][120] ));
 sky130_fd_sc_hd__dfxtp_1 _17087_ (.CLK(net491),
    .D(_00530_),
    .Q(\fifo_bank_register.bank[7][121] ));
 sky130_fd_sc_hd__dfxtp_1 _17088_ (.CLK(net493),
    .D(_00531_),
    .Q(\fifo_bank_register.bank[7][122] ));
 sky130_fd_sc_hd__dfxtp_1 _17089_ (.CLK(net440),
    .D(_00532_),
    .Q(\fifo_bank_register.bank[7][123] ));
 sky130_fd_sc_hd__dfxtp_1 _17090_ (.CLK(net494),
    .D(_00533_),
    .Q(\fifo_bank_register.bank[7][124] ));
 sky130_fd_sc_hd__dfxtp_1 _17091_ (.CLK(net496),
    .D(_00534_),
    .Q(\fifo_bank_register.bank[7][125] ));
 sky130_fd_sc_hd__dfxtp_1 _17092_ (.CLK(net494),
    .D(_00535_),
    .Q(\fifo_bank_register.bank[7][126] ));
 sky130_fd_sc_hd__dfxtp_1 _17093_ (.CLK(net441),
    .D(_00536_),
    .Q(\fifo_bank_register.bank[7][127] ));
 sky130_fd_sc_hd__dfxtp_1 _17094_ (.CLK(net481),
    .D(_00537_),
    .Q(\fifo_bank_register.bank[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17095_ (.CLK(net490),
    .D(_00538_),
    .Q(\fifo_bank_register.bank[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17096_ (.CLK(net474),
    .D(_00539_),
    .Q(\fifo_bank_register.bank[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17097_ (.CLK(net473),
    .D(_00540_),
    .Q(\fifo_bank_register.bank[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17098_ (.CLK(net474),
    .D(_00541_),
    .Q(\fifo_bank_register.bank[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17099_ (.CLK(net473),
    .D(_00542_),
    .Q(\fifo_bank_register.bank[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17100_ (.CLK(net477),
    .D(_00543_),
    .Q(\fifo_bank_register.bank[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17101_ (.CLK(net477),
    .D(_00544_),
    .Q(\fifo_bank_register.bank[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17102_ (.CLK(net478),
    .D(_00545_),
    .Q(\fifo_bank_register.bank[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17103_ (.CLK(net478),
    .D(_00546_),
    .Q(\fifo_bank_register.bank[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17104_ (.CLK(net504),
    .D(_00547_),
    .Q(\fifo_bank_register.bank[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17105_ (.CLK(net535),
    .D(_00548_),
    .Q(\fifo_bank_register.bank[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17106_ (.CLK(net504),
    .D(_00549_),
    .Q(\fifo_bank_register.bank[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17107_ (.CLK(net505),
    .D(_00550_),
    .Q(\fifo_bank_register.bank[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17108_ (.CLK(net534),
    .D(_00551_),
    .Q(\fifo_bank_register.bank[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17109_ (.CLK(net534),
    .D(_00552_),
    .Q(\fifo_bank_register.bank[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17110_ (.CLK(net496),
    .D(_00553_),
    .Q(\fifo_bank_register.bank[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17111_ (.CLK(net532),
    .D(_00554_),
    .Q(\fifo_bank_register.bank[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17112_ (.CLK(net533),
    .D(_00555_),
    .Q(\fifo_bank_register.bank[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17113_ (.CLK(net505),
    .D(_00556_),
    .Q(\fifo_bank_register.bank[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17114_ (.CLK(net512),
    .D(_00557_),
    .Q(\fifo_bank_register.bank[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17115_ (.CLK(net484),
    .D(_00558_),
    .Q(\fifo_bank_register.bank[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17116_ (.CLK(net502),
    .D(_00559_),
    .Q(\fifo_bank_register.bank[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17117_ (.CLK(net483),
    .D(_00560_),
    .Q(\fifo_bank_register.bank[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17118_ (.CLK(net485),
    .D(_00561_),
    .Q(\fifo_bank_register.bank[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17119_ (.CLK(net508),
    .D(_00562_),
    .Q(\fifo_bank_register.bank[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17120_ (.CLK(net510),
    .D(_00563_),
    .Q(\fifo_bank_register.bank[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17121_ (.CLK(net499),
    .D(_00564_),
    .Q(\fifo_bank_register.bank[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17122_ (.CLK(net485),
    .D(_00565_),
    .Q(\fifo_bank_register.bank[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17123_ (.CLK(net499),
    .D(_00566_),
    .Q(\fifo_bank_register.bank[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17124_ (.CLK(net430),
    .D(_00567_),
    .Q(\fifo_bank_register.bank[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17125_ (.CLK(net437),
    .D(_00568_),
    .Q(\fifo_bank_register.bank[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17126_ (.CLK(net422),
    .D(_00569_),
    .Q(\fifo_bank_register.bank[6][32] ));
 sky130_fd_sc_hd__dfxtp_1 _17127_ (.CLK(net423),
    .D(_00570_),
    .Q(\fifo_bank_register.bank[6][33] ));
 sky130_fd_sc_hd__dfxtp_1 _17128_ (.CLK(net431),
    .D(_00571_),
    .Q(\fifo_bank_register.bank[6][34] ));
 sky130_fd_sc_hd__dfxtp_1 _17129_ (.CLK(net429),
    .D(_00572_),
    .Q(\fifo_bank_register.bank[6][35] ));
 sky130_fd_sc_hd__dfxtp_1 _17130_ (.CLK(net422),
    .D(_00573_),
    .Q(\fifo_bank_register.bank[6][36] ));
 sky130_fd_sc_hd__dfxtp_1 _17131_ (.CLK(net414),
    .D(_00574_),
    .Q(\fifo_bank_register.bank[6][37] ));
 sky130_fd_sc_hd__dfxtp_1 _17132_ (.CLK(net417),
    .D(_00575_),
    .Q(\fifo_bank_register.bank[6][38] ));
 sky130_fd_sc_hd__dfxtp_1 _17133_ (.CLK(net415),
    .D(_00576_),
    .Q(\fifo_bank_register.bank[6][39] ));
 sky130_fd_sc_hd__dfxtp_1 _17134_ (.CLK(net395),
    .D(_00577_),
    .Q(\fifo_bank_register.bank[6][40] ));
 sky130_fd_sc_hd__dfxtp_1 _17135_ (.CLK(net399),
    .D(_00578_),
    .Q(\fifo_bank_register.bank[6][41] ));
 sky130_fd_sc_hd__dfxtp_1 _17136_ (.CLK(net406),
    .D(_00579_),
    .Q(\fifo_bank_register.bank[6][42] ));
 sky130_fd_sc_hd__dfxtp_1 _17137_ (.CLK(net393),
    .D(_00580_),
    .Q(\fifo_bank_register.bank[6][43] ));
 sky130_fd_sc_hd__dfxtp_1 _17138_ (.CLK(net389),
    .D(_00581_),
    .Q(\fifo_bank_register.bank[6][44] ));
 sky130_fd_sc_hd__dfxtp_1 _17139_ (.CLK(net406),
    .D(_00582_),
    .Q(\fifo_bank_register.bank[6][45] ));
 sky130_fd_sc_hd__dfxtp_1 _17140_ (.CLK(net390),
    .D(_00583_),
    .Q(\fifo_bank_register.bank[6][46] ));
 sky130_fd_sc_hd__dfxtp_1 _17141_ (.CLK(net396),
    .D(_00584_),
    .Q(\fifo_bank_register.bank[6][47] ));
 sky130_fd_sc_hd__dfxtp_1 _17142_ (.CLK(net395),
    .D(_00585_),
    .Q(\fifo_bank_register.bank[6][48] ));
 sky130_fd_sc_hd__dfxtp_1 _17143_ (.CLK(net407),
    .D(_00586_),
    .Q(\fifo_bank_register.bank[6][49] ));
 sky130_fd_sc_hd__dfxtp_1 _17144_ (.CLK(net572),
    .D(_00587_),
    .Q(\fifo_bank_register.bank[6][50] ));
 sky130_fd_sc_hd__dfxtp_1 _17145_ (.CLK(net575),
    .D(_00588_),
    .Q(\fifo_bank_register.bank[6][51] ));
 sky130_fd_sc_hd__dfxtp_1 _17146_ (.CLK(net567),
    .D(_00589_),
    .Q(\fifo_bank_register.bank[6][52] ));
 sky130_fd_sc_hd__dfxtp_1 _17147_ (.CLK(net567),
    .D(_00590_),
    .Q(\fifo_bank_register.bank[6][53] ));
 sky130_fd_sc_hd__dfxtp_1 _17148_ (.CLK(net556),
    .D(_00591_),
    .Q(\fifo_bank_register.bank[6][54] ));
 sky130_fd_sc_hd__dfxtp_1 _17149_ (.CLK(net574),
    .D(_00592_),
    .Q(\fifo_bank_register.bank[6][55] ));
 sky130_fd_sc_hd__dfxtp_1 _17150_ (.CLK(net574),
    .D(_00593_),
    .Q(\fifo_bank_register.bank[6][56] ));
 sky130_fd_sc_hd__dfxtp_1 _17151_ (.CLK(net549),
    .D(_00594_),
    .Q(\fifo_bank_register.bank[6][57] ));
 sky130_fd_sc_hd__dfxtp_1 _17152_ (.CLK(net558),
    .D(_00595_),
    .Q(\fifo_bank_register.bank[6][58] ));
 sky130_fd_sc_hd__dfxtp_1 _17153_ (.CLK(net573),
    .D(_00596_),
    .Q(\fifo_bank_register.bank[6][59] ));
 sky130_fd_sc_hd__dfxtp_1 _17154_ (.CLK(net515),
    .D(_00597_),
    .Q(\fifo_bank_register.bank[6][60] ));
 sky130_fd_sc_hd__dfxtp_1 _17155_ (.CLK(net527),
    .D(_00598_),
    .Q(\fifo_bank_register.bank[6][61] ));
 sky130_fd_sc_hd__dfxtp_1 _17156_ (.CLK(net523),
    .D(_00599_),
    .Q(\fifo_bank_register.bank[6][62] ));
 sky130_fd_sc_hd__dfxtp_1 _17157_ (.CLK(net523),
    .D(_00600_),
    .Q(\fifo_bank_register.bank[6][63] ));
 sky130_fd_sc_hd__dfxtp_1 _17158_ (.CLK(net514),
    .D(_00601_),
    .Q(\fifo_bank_register.bank[6][64] ));
 sky130_fd_sc_hd__dfxtp_1 _17159_ (.CLK(net518),
    .D(_00602_),
    .Q(\fifo_bank_register.bank[6][65] ));
 sky130_fd_sc_hd__dfxtp_1 _17160_ (.CLK(net523),
    .D(_00603_),
    .Q(\fifo_bank_register.bank[6][66] ));
 sky130_fd_sc_hd__dfxtp_1 _17161_ (.CLK(net514),
    .D(_00604_),
    .Q(\fifo_bank_register.bank[6][67] ));
 sky130_fd_sc_hd__dfxtp_1 _17162_ (.CLK(net521),
    .D(_00605_),
    .Q(\fifo_bank_register.bank[6][68] ));
 sky130_fd_sc_hd__dfxtp_1 _17163_ (.CLK(net514),
    .D(_00606_),
    .Q(\fifo_bank_register.bank[6][69] ));
 sky130_fd_sc_hd__dfxtp_1 _17164_ (.CLK(net518),
    .D(_00607_),
    .Q(\fifo_bank_register.bank[6][70] ));
 sky130_fd_sc_hd__dfxtp_1 _17165_ (.CLK(net527),
    .D(_00608_),
    .Q(\fifo_bank_register.bank[6][71] ));
 sky130_fd_sc_hd__dfxtp_1 _17166_ (.CLK(net554),
    .D(_00609_),
    .Q(\fifo_bank_register.bank[6][72] ));
 sky130_fd_sc_hd__dfxtp_1 _17167_ (.CLK(net554),
    .D(_00610_),
    .Q(\fifo_bank_register.bank[6][73] ));
 sky130_fd_sc_hd__dfxtp_1 _17168_ (.CLK(net546),
    .D(_00611_),
    .Q(\fifo_bank_register.bank[6][74] ));
 sky130_fd_sc_hd__dfxtp_1 _17169_ (.CLK(net552),
    .D(_00612_),
    .Q(\fifo_bank_register.bank[6][75] ));
 sky130_fd_sc_hd__dfxtp_1 _17170_ (.CLK(net545),
    .D(_00613_),
    .Q(\fifo_bank_register.bank[6][76] ));
 sky130_fd_sc_hd__dfxtp_1 _17171_ (.CLK(net554),
    .D(_00614_),
    .Q(\fifo_bank_register.bank[6][77] ));
 sky130_fd_sc_hd__dfxtp_1 _17172_ (.CLK(net525),
    .D(_00615_),
    .Q(\fifo_bank_register.bank[6][78] ));
 sky130_fd_sc_hd__dfxtp_1 _17173_ (.CLK(net553),
    .D(_00616_),
    .Q(\fifo_bank_register.bank[6][79] ));
 sky130_fd_sc_hd__dfxtp_1 _17174_ (.CLK(net565),
    .D(_00617_),
    .Q(\fifo_bank_register.bank[6][80] ));
 sky130_fd_sc_hd__dfxtp_1 _17175_ (.CLK(net564),
    .D(_00618_),
    .Q(\fifo_bank_register.bank[6][81] ));
 sky130_fd_sc_hd__dfxtp_1 _17176_ (.CLK(net550),
    .D(_00619_),
    .Q(\fifo_bank_register.bank[6][82] ));
 sky130_fd_sc_hd__dfxtp_1 _17177_ (.CLK(net561),
    .D(_00620_),
    .Q(\fifo_bank_register.bank[6][83] ));
 sky130_fd_sc_hd__dfxtp_1 _17178_ (.CLK(net547),
    .D(_00621_),
    .Q(\fifo_bank_register.bank[6][84] ));
 sky130_fd_sc_hd__dfxtp_1 _17179_ (.CLK(net567),
    .D(_00622_),
    .Q(\fifo_bank_register.bank[6][85] ));
 sky130_fd_sc_hd__dfxtp_1 _17180_ (.CLK(net561),
    .D(_00623_),
    .Q(\fifo_bank_register.bank[6][86] ));
 sky130_fd_sc_hd__dfxtp_1 _17181_ (.CLK(net560),
    .D(_00624_),
    .Q(\fifo_bank_register.bank[6][87] ));
 sky130_fd_sc_hd__dfxtp_1 _17182_ (.CLK(net565),
    .D(_00625_),
    .Q(\fifo_bank_register.bank[6][88] ));
 sky130_fd_sc_hd__dfxtp_1 _17183_ (.CLK(net548),
    .D(_00626_),
    .Q(\fifo_bank_register.bank[6][89] ));
 sky130_fd_sc_hd__dfxtp_1 _17184_ (.CLK(net409),
    .D(_00627_),
    .Q(\fifo_bank_register.bank[6][90] ));
 sky130_fd_sc_hd__dfxtp_1 _17185_ (.CLK(net401),
    .D(_00628_),
    .Q(\fifo_bank_register.bank[6][91] ));
 sky130_fd_sc_hd__dfxtp_1 _17186_ (.CLK(net410),
    .D(_00629_),
    .Q(\fifo_bank_register.bank[6][92] ));
 sky130_fd_sc_hd__dfxtp_1 _17187_ (.CLK(net402),
    .D(_00630_),
    .Q(\fifo_bank_register.bank[6][93] ));
 sky130_fd_sc_hd__dfxtp_1 _17188_ (.CLK(net455),
    .D(_00631_),
    .Q(\fifo_bank_register.bank[6][94] ));
 sky130_fd_sc_hd__dfxtp_1 _17189_ (.CLK(net402),
    .D(_00632_),
    .Q(\fifo_bank_register.bank[6][95] ));
 sky130_fd_sc_hd__dfxtp_1 _17190_ (.CLK(net448),
    .D(_00633_),
    .Q(\fifo_bank_register.bank[6][96] ));
 sky130_fd_sc_hd__dfxtp_1 _17191_ (.CLK(net454),
    .D(_00634_),
    .Q(\fifo_bank_register.bank[6][97] ));
 sky130_fd_sc_hd__dfxtp_1 _17192_ (.CLK(net447),
    .D(_00635_),
    .Q(\fifo_bank_register.bank[6][98] ));
 sky130_fd_sc_hd__dfxtp_1 _17193_ (.CLK(net446),
    .D(_00636_),
    .Q(\fifo_bank_register.bank[6][99] ));
 sky130_fd_sc_hd__dfxtp_1 _17194_ (.CLK(net453),
    .D(_00637_),
    .Q(\fifo_bank_register.bank[6][100] ));
 sky130_fd_sc_hd__dfxtp_1 _17195_ (.CLK(net450),
    .D(_00638_),
    .Q(\fifo_bank_register.bank[6][101] ));
 sky130_fd_sc_hd__dfxtp_1 _17196_ (.CLK(net465),
    .D(_00639_),
    .Q(\fifo_bank_register.bank[6][102] ));
 sky130_fd_sc_hd__dfxtp_1 _17197_ (.CLK(net467),
    .D(_00640_),
    .Q(\fifo_bank_register.bank[6][103] ));
 sky130_fd_sc_hd__dfxtp_1 _17198_ (.CLK(net463),
    .D(_00641_),
    .Q(\fifo_bank_register.bank[6][104] ));
 sky130_fd_sc_hd__dfxtp_1 _17199_ (.CLK(net467),
    .D(_00642_),
    .Q(\fifo_bank_register.bank[6][105] ));
 sky130_fd_sc_hd__dfxtp_1 _17200_ (.CLK(net465),
    .D(_00643_),
    .Q(\fifo_bank_register.bank[6][106] ));
 sky130_fd_sc_hd__dfxtp_1 _17201_ (.CLK(net451),
    .D(_00644_),
    .Q(\fifo_bank_register.bank[6][107] ));
 sky130_fd_sc_hd__dfxtp_1 _17202_ (.CLK(net453),
    .D(_00645_),
    .Q(\fifo_bank_register.bank[6][108] ));
 sky130_fd_sc_hd__dfxtp_1 _17203_ (.CLK(net459),
    .D(_00646_),
    .Q(\fifo_bank_register.bank[6][109] ));
 sky130_fd_sc_hd__dfxtp_1 _17204_ (.CLK(net471),
    .D(_00647_),
    .Q(\fifo_bank_register.bank[6][110] ));
 sky130_fd_sc_hd__dfxtp_1 _17205_ (.CLK(net411),
    .D(_00648_),
    .Q(\fifo_bank_register.bank[6][111] ));
 sky130_fd_sc_hd__dfxtp_1 _17206_ (.CLK(net433),
    .D(_00649_),
    .Q(\fifo_bank_register.bank[6][112] ));
 sky130_fd_sc_hd__dfxtp_1 _17207_ (.CLK(net469),
    .D(_00650_),
    .Q(\fifo_bank_register.bank[6][113] ));
 sky130_fd_sc_hd__dfxtp_1 _17208_ (.CLK(net456),
    .D(_00651_),
    .Q(\fifo_bank_register.bank[6][114] ));
 sky130_fd_sc_hd__dfxtp_1 _17209_ (.CLK(net470),
    .D(_00652_),
    .Q(\fifo_bank_register.bank[6][115] ));
 sky130_fd_sc_hd__dfxtp_1 _17210_ (.CLK(net411),
    .D(_00653_),
    .Q(\fifo_bank_register.bank[6][116] ));
 sky130_fd_sc_hd__dfxtp_1 _17211_ (.CLK(net435),
    .D(_00654_),
    .Q(\fifo_bank_register.bank[6][117] ));
 sky130_fd_sc_hd__dfxtp_1 _17212_ (.CLK(net469),
    .D(_00655_),
    .Q(\fifo_bank_register.bank[6][118] ));
 sky130_fd_sc_hd__dfxtp_1 _17213_ (.CLK(net435),
    .D(_00656_),
    .Q(\fifo_bank_register.bank[6][119] ));
 sky130_fd_sc_hd__dfxtp_1 _17214_ (.CLK(net441),
    .D(_00657_),
    .Q(\fifo_bank_register.bank[6][120] ));
 sky130_fd_sc_hd__dfxtp_1 _17215_ (.CLK(net440),
    .D(_00658_),
    .Q(\fifo_bank_register.bank[6][121] ));
 sky130_fd_sc_hd__dfxtp_1 _17216_ (.CLK(net490),
    .D(_00659_),
    .Q(\fifo_bank_register.bank[6][122] ));
 sky130_fd_sc_hd__dfxtp_1 _17217_ (.CLK(net439),
    .D(_00660_),
    .Q(\fifo_bank_register.bank[6][123] ));
 sky130_fd_sc_hd__dfxtp_1 _17218_ (.CLK(net495),
    .D(_00661_),
    .Q(\fifo_bank_register.bank[6][124] ));
 sky130_fd_sc_hd__dfxtp_1 _17219_ (.CLK(net496),
    .D(_00662_),
    .Q(\fifo_bank_register.bank[6][125] ));
 sky130_fd_sc_hd__dfxtp_1 _17220_ (.CLK(net495),
    .D(_00663_),
    .Q(\fifo_bank_register.bank[6][126] ));
 sky130_fd_sc_hd__dfxtp_1 _17221_ (.CLK(net441),
    .D(_00664_),
    .Q(\fifo_bank_register.bank[6][127] ));
 sky130_fd_sc_hd__dfxtp_1 _17222_ (.CLK(net475),
    .D(_00665_),
    .Q(\fifo_bank_register.bank[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17223_ (.CLK(net492),
    .D(_00666_),
    .Q(\fifo_bank_register.bank[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17224_ (.CLK(net476),
    .D(_00667_),
    .Q(\fifo_bank_register.bank[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17225_ (.CLK(net475),
    .D(_00668_),
    .Q(\fifo_bank_register.bank[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17226_ (.CLK(net476),
    .D(_00669_),
    .Q(\fifo_bank_register.bank[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17227_ (.CLK(net476),
    .D(_00670_),
    .Q(\fifo_bank_register.bank[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17228_ (.CLK(net479),
    .D(_00671_),
    .Q(\fifo_bank_register.bank[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17229_ (.CLK(net479),
    .D(_00672_),
    .Q(\fifo_bank_register.bank[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17230_ (.CLK(net492),
    .D(_00673_),
    .Q(\fifo_bank_register.bank[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17231_ (.CLK(net479),
    .D(_00674_),
    .Q(\fifo_bank_register.bank[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17232_ (.CLK(net493),
    .D(_00675_),
    .Q(\fifo_bank_register.bank[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17233_ (.CLK(net504),
    .D(_00676_),
    .Q(\fifo_bank_register.bank[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17234_ (.CLK(net500),
    .D(_00677_),
    .Q(\fifo_bank_register.bank[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17235_ (.CLK(net504),
    .D(_00678_),
    .Q(\fifo_bank_register.bank[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17236_ (.CLK(net506),
    .D(_00679_),
    .Q(\fifo_bank_register.bank[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17237_ (.CLK(net506),
    .D(_00680_),
    .Q(\fifo_bank_register.bank[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17238_ (.CLK(net493),
    .D(_00681_),
    .Q(\fifo_bank_register.bank[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17239_ (.CLK(net497),
    .D(_00682_),
    .Q(\fifo_bank_register.bank[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17240_ (.CLK(net503),
    .D(_00683_),
    .Q(\fifo_bank_register.bank[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17241_ (.CLK(net502),
    .D(_00684_),
    .Q(\fifo_bank_register.bank[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17242_ (.CLK(net487),
    .D(_00685_),
    .Q(\fifo_bank_register.bank[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17243_ (.CLK(net487),
    .D(_00686_),
    .Q(\fifo_bank_register.bank[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17244_ (.CLK(net488),
    .D(_00687_),
    .Q(\fifo_bank_register.bank[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17245_ (.CLK(net487),
    .D(_00688_),
    .Q(\fifo_bank_register.bank[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17246_ (.CLK(net485),
    .D(_00689_),
    .Q(\fifo_bank_register.bank[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17247_ (.CLK(net487),
    .D(_00690_),
    .Q(\fifo_bank_register.bank[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17248_ (.CLK(net508),
    .D(_00691_),
    .Q(\fifo_bank_register.bank[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17249_ (.CLK(net488),
    .D(_00692_),
    .Q(\fifo_bank_register.bank[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17250_ (.CLK(net488),
    .D(_00693_),
    .Q(\fifo_bank_register.bank[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17251_ (.CLK(net499),
    .D(_00694_),
    .Q(\fifo_bank_register.bank[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17252_ (.CLK(net418),
    .D(_00695_),
    .Q(\fifo_bank_register.bank[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17253_ (.CLK(net424),
    .D(_00696_),
    .Q(\fifo_bank_register.bank[5][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17254_ (.CLK(net419),
    .D(_00697_),
    .Q(\fifo_bank_register.bank[5][32] ));
 sky130_fd_sc_hd__dfxtp_1 _17255_ (.CLK(net424),
    .D(_00698_),
    .Q(\fifo_bank_register.bank[5][33] ));
 sky130_fd_sc_hd__dfxtp_1 _17256_ (.CLK(net418),
    .D(_00699_),
    .Q(\fifo_bank_register.bank[5][34] ));
 sky130_fd_sc_hd__dfxtp_1 _17257_ (.CLK(net416),
    .D(_00700_),
    .Q(\fifo_bank_register.bank[5][35] ));
 sky130_fd_sc_hd__dfxtp_1 _17258_ (.CLK(net422),
    .D(_00701_),
    .Q(\fifo_bank_register.bank[5][36] ));
 sky130_fd_sc_hd__dfxtp_1 _17259_ (.CLK(net414),
    .D(_00702_),
    .Q(\fifo_bank_register.bank[5][37] ));
 sky130_fd_sc_hd__dfxtp_1 _17260_ (.CLK(net416),
    .D(_00703_),
    .Q(\fifo_bank_register.bank[5][38] ));
 sky130_fd_sc_hd__dfxtp_1 _17261_ (.CLK(net414),
    .D(_00704_),
    .Q(\fifo_bank_register.bank[5][39] ));
 sky130_fd_sc_hd__dfxtp_1 _17262_ (.CLK(net392),
    .D(_00705_),
    .Q(\fifo_bank_register.bank[5][40] ));
 sky130_fd_sc_hd__dfxtp_1 _17263_ (.CLK(net398),
    .D(_00706_),
    .Q(\fifo_bank_register.bank[5][41] ));
 sky130_fd_sc_hd__dfxtp_1 _17264_ (.CLK(net390),
    .D(_00707_),
    .Q(\fifo_bank_register.bank[5][42] ));
 sky130_fd_sc_hd__dfxtp_1 _17265_ (.CLK(net392),
    .D(_00708_),
    .Q(\fifo_bank_register.bank[5][43] ));
 sky130_fd_sc_hd__dfxtp_1 _17266_ (.CLK(net391),
    .D(_00709_),
    .Q(\fifo_bank_register.bank[5][44] ));
 sky130_fd_sc_hd__dfxtp_1 _17267_ (.CLK(net394),
    .D(_00710_),
    .Q(\fifo_bank_register.bank[5][45] ));
 sky130_fd_sc_hd__dfxtp_1 _17268_ (.CLK(net391),
    .D(_00711_),
    .Q(\fifo_bank_register.bank[5][46] ));
 sky130_fd_sc_hd__dfxtp_1 _17269_ (.CLK(net396),
    .D(_00712_),
    .Q(\fifo_bank_register.bank[5][47] ));
 sky130_fd_sc_hd__dfxtp_1 _17270_ (.CLK(net397),
    .D(_00713_),
    .Q(\fifo_bank_register.bank[5][48] ));
 sky130_fd_sc_hd__dfxtp_1 _17271_ (.CLK(net407),
    .D(_00714_),
    .Q(\fifo_bank_register.bank[5][49] ));
 sky130_fd_sc_hd__dfxtp_1 _17272_ (.CLK(net555),
    .D(_00715_),
    .Q(\fifo_bank_register.bank[5][50] ));
 sky130_fd_sc_hd__dfxtp_1 _17273_ (.CLK(net572),
    .D(_00716_),
    .Q(\fifo_bank_register.bank[5][51] ));
 sky130_fd_sc_hd__dfxtp_1 _17274_ (.CLK(net562),
    .D(_00717_),
    .Q(\fifo_bank_register.bank[5][52] ));
 sky130_fd_sc_hd__dfxtp_1 _17275_ (.CLK(net562),
    .D(_00718_),
    .Q(\fifo_bank_register.bank[5][53] ));
 sky130_fd_sc_hd__dfxtp_1 _17276_ (.CLK(net555),
    .D(_00719_),
    .Q(\fifo_bank_register.bank[5][54] ));
 sky130_fd_sc_hd__dfxtp_1 _17277_ (.CLK(net570),
    .D(_00720_),
    .Q(\fifo_bank_register.bank[5][55] ));
 sky130_fd_sc_hd__dfxtp_1 _17278_ (.CLK(net570),
    .D(_00721_),
    .Q(\fifo_bank_register.bank[5][56] ));
 sky130_fd_sc_hd__dfxtp_1 _17279_ (.CLK(net549),
    .D(_00722_),
    .Q(\fifo_bank_register.bank[5][57] ));
 sky130_fd_sc_hd__dfxtp_1 _17280_ (.CLK(net555),
    .D(_00723_),
    .Q(\fifo_bank_register.bank[5][58] ));
 sky130_fd_sc_hd__dfxtp_1 _17281_ (.CLK(net570),
    .D(_00724_),
    .Q(\fifo_bank_register.bank[5][59] ));
 sky130_fd_sc_hd__dfxtp_1 _17282_ (.CLK(net512),
    .D(_00725_),
    .Q(\fifo_bank_register.bank[5][60] ));
 sky130_fd_sc_hd__dfxtp_1 _17283_ (.CLK(net526),
    .D(_00726_),
    .Q(\fifo_bank_register.bank[5][61] ));
 sky130_fd_sc_hd__dfxtp_1 _17284_ (.CLK(net521),
    .D(_00727_),
    .Q(\fifo_bank_register.bank[5][62] ));
 sky130_fd_sc_hd__dfxtp_1 _17285_ (.CLK(net522),
    .D(_00728_),
    .Q(\fifo_bank_register.bank[5][63] ));
 sky130_fd_sc_hd__dfxtp_1 _17286_ (.CLK(net512),
    .D(_00729_),
    .Q(\fifo_bank_register.bank[5][64] ));
 sky130_fd_sc_hd__dfxtp_1 _17287_ (.CLK(net521),
    .D(_00730_),
    .Q(\fifo_bank_register.bank[5][65] ));
 sky130_fd_sc_hd__dfxtp_1 _17288_ (.CLK(net522),
    .D(_00731_),
    .Q(\fifo_bank_register.bank[5][66] ));
 sky130_fd_sc_hd__dfxtp_1 _17289_ (.CLK(net522),
    .D(_00732_),
    .Q(\fifo_bank_register.bank[5][67] ));
 sky130_fd_sc_hd__dfxtp_1 _17290_ (.CLK(net522),
    .D(_00733_),
    .Q(\fifo_bank_register.bank[5][68] ));
 sky130_fd_sc_hd__dfxtp_1 _17291_ (.CLK(net512),
    .D(_00734_),
    .Q(\fifo_bank_register.bank[5][69] ));
 sky130_fd_sc_hd__dfxtp_1 _17292_ (.CLK(net517),
    .D(_00735_),
    .Q(\fifo_bank_register.bank[5][70] ));
 sky130_fd_sc_hd__dfxtp_1 _17293_ (.CLK(net517),
    .D(_00736_),
    .Q(\fifo_bank_register.bank[5][71] ));
 sky130_fd_sc_hd__dfxtp_1 _17294_ (.CLK(net544),
    .D(_00737_),
    .Q(\fifo_bank_register.bank[5][72] ));
 sky130_fd_sc_hd__dfxtp_1 _17295_ (.CLK(net543),
    .D(_00738_),
    .Q(\fifo_bank_register.bank[5][73] ));
 sky130_fd_sc_hd__dfxtp_1 _17296_ (.CLK(net544),
    .D(_00739_),
    .Q(\fifo_bank_register.bank[5][74] ));
 sky130_fd_sc_hd__dfxtp_1 _17297_ (.CLK(net543),
    .D(_00740_),
    .Q(\fifo_bank_register.bank[5][75] ));
 sky130_fd_sc_hd__dfxtp_1 _17298_ (.CLK(net543),
    .D(_00741_),
    .Q(\fifo_bank_register.bank[5][76] ));
 sky130_fd_sc_hd__dfxtp_1 _17299_ (.CLK(net544),
    .D(_00742_),
    .Q(\fifo_bank_register.bank[5][77] ));
 sky130_fd_sc_hd__dfxtp_1 _17300_ (.CLK(net517),
    .D(_00743_),
    .Q(\fifo_bank_register.bank[5][78] ));
 sky130_fd_sc_hd__dfxtp_1 _17301_ (.CLK(net543),
    .D(_00744_),
    .Q(\fifo_bank_register.bank[5][79] ));
 sky130_fd_sc_hd__dfxtp_1 _17302_ (.CLK(net541),
    .D(_00745_),
    .Q(\fifo_bank_register.bank[5][80] ));
 sky130_fd_sc_hd__dfxtp_1 _17303_ (.CLK(net540),
    .D(_00746_),
    .Q(\fifo_bank_register.bank[5][81] ));
 sky130_fd_sc_hd__dfxtp_1 _17304_ (.CLK(net539),
    .D(_00747_),
    .Q(\fifo_bank_register.bank[5][82] ));
 sky130_fd_sc_hd__dfxtp_1 _17305_ (.CLK(net539),
    .D(_00748_),
    .Q(\fifo_bank_register.bank[5][83] ));
 sky130_fd_sc_hd__dfxtp_1 _17306_ (.CLK(net536),
    .D(_00749_),
    .Q(\fifo_bank_register.bank[5][84] ));
 sky130_fd_sc_hd__dfxtp_1 _17307_ (.CLK(net540),
    .D(_00750_),
    .Q(\fifo_bank_register.bank[5][85] ));
 sky130_fd_sc_hd__dfxtp_1 _17308_ (.CLK(net536),
    .D(_00751_),
    .Q(\fifo_bank_register.bank[5][86] ));
 sky130_fd_sc_hd__dfxtp_1 _17309_ (.CLK(net538),
    .D(_00752_),
    .Q(\fifo_bank_register.bank[5][87] ));
 sky130_fd_sc_hd__dfxtp_1 _17310_ (.CLK(net541),
    .D(_00753_),
    .Q(\fifo_bank_register.bank[5][88] ));
 sky130_fd_sc_hd__dfxtp_1 _17311_ (.CLK(net536),
    .D(_00754_),
    .Q(\fifo_bank_register.bank[5][89] ));
 sky130_fd_sc_hd__dfxtp_1 _17312_ (.CLK(net409),
    .D(_00755_),
    .Q(\fifo_bank_register.bank[5][90] ));
 sky130_fd_sc_hd__dfxtp_1 _17313_ (.CLK(net401),
    .D(_00756_),
    .Q(\fifo_bank_register.bank[5][91] ));
 sky130_fd_sc_hd__dfxtp_1 _17314_ (.CLK(net403),
    .D(_00757_),
    .Q(\fifo_bank_register.bank[5][92] ));
 sky130_fd_sc_hd__dfxtp_1 _17315_ (.CLK(net400),
    .D(_00758_),
    .Q(\fifo_bank_register.bank[5][93] ));
 sky130_fd_sc_hd__dfxtp_1 _17316_ (.CLK(net448),
    .D(_00759_),
    .Q(\fifo_bank_register.bank[5][94] ));
 sky130_fd_sc_hd__dfxtp_1 _17317_ (.CLK(net400),
    .D(_00760_),
    .Q(\fifo_bank_register.bank[5][95] ));
 sky130_fd_sc_hd__dfxtp_1 _17318_ (.CLK(net401),
    .D(_00761_),
    .Q(\fifo_bank_register.bank[5][96] ));
 sky130_fd_sc_hd__dfxtp_1 _17319_ (.CLK(net448),
    .D(_00762_),
    .Q(\fifo_bank_register.bank[5][97] ));
 sky130_fd_sc_hd__dfxtp_1 _17320_ (.CLK(net445),
    .D(_00763_),
    .Q(\fifo_bank_register.bank[5][98] ));
 sky130_fd_sc_hd__dfxtp_1 _17321_ (.CLK(net445),
    .D(_00764_),
    .Q(\fifo_bank_register.bank[5][99] ));
 sky130_fd_sc_hd__dfxtp_1 _17322_ (.CLK(net452),
    .D(_00765_),
    .Q(\fifo_bank_register.bank[5][100] ));
 sky130_fd_sc_hd__dfxtp_1 _17323_ (.CLK(net446),
    .D(_00766_),
    .Q(\fifo_bank_register.bank[5][101] ));
 sky130_fd_sc_hd__dfxtp_1 _17324_ (.CLK(net464),
    .D(_00767_),
    .Q(\fifo_bank_register.bank[5][102] ));
 sky130_fd_sc_hd__dfxtp_1 _17325_ (.CLK(net464),
    .D(_00768_),
    .Q(\fifo_bank_register.bank[5][103] ));
 sky130_fd_sc_hd__dfxtp_1 _17326_ (.CLK(net462),
    .D(_00769_),
    .Q(\fifo_bank_register.bank[5][104] ));
 sky130_fd_sc_hd__dfxtp_1 _17327_ (.CLK(net467),
    .D(_00770_),
    .Q(\fifo_bank_register.bank[5][105] ));
 sky130_fd_sc_hd__dfxtp_1 _17328_ (.CLK(net464),
    .D(_00771_),
    .Q(\fifo_bank_register.bank[5][106] ));
 sky130_fd_sc_hd__dfxtp_1 _17329_ (.CLK(net462),
    .D(_00772_),
    .Q(\fifo_bank_register.bank[5][107] ));
 sky130_fd_sc_hd__dfxtp_1 _17330_ (.CLK(net447),
    .D(_00773_),
    .Q(\fifo_bank_register.bank[5][108] ));
 sky130_fd_sc_hd__dfxtp_1 _17331_ (.CLK(net454),
    .D(_00774_),
    .Q(\fifo_bank_register.bank[5][109] ));
 sky130_fd_sc_hd__dfxtp_1 _17332_ (.CLK(net432),
    .D(_00775_),
    .Q(\fifo_bank_register.bank[5][110] ));
 sky130_fd_sc_hd__dfxtp_1 _17333_ (.CLK(net412),
    .D(_00776_),
    .Q(\fifo_bank_register.bank[5][111] ));
 sky130_fd_sc_hd__dfxtp_1 _17334_ (.CLK(net412),
    .D(_00777_),
    .Q(\fifo_bank_register.bank[5][112] ));
 sky130_fd_sc_hd__dfxtp_1 _17335_ (.CLK(net429),
    .D(_00778_),
    .Q(\fifo_bank_register.bank[5][113] ));
 sky130_fd_sc_hd__dfxtp_1 _17336_ (.CLK(net408),
    .D(_00779_),
    .Q(\fifo_bank_register.bank[5][114] ));
 sky130_fd_sc_hd__dfxtp_1 _17337_ (.CLK(net429),
    .D(_00780_),
    .Q(\fifo_bank_register.bank[5][115] ));
 sky130_fd_sc_hd__dfxtp_1 _17338_ (.CLK(net412),
    .D(_00781_),
    .Q(\fifo_bank_register.bank[5][116] ));
 sky130_fd_sc_hd__dfxtp_1 _17339_ (.CLK(net434),
    .D(_00782_),
    .Q(\fifo_bank_register.bank[5][117] ));
 sky130_fd_sc_hd__dfxtp_1 _17340_ (.CLK(net408),
    .D(_00783_),
    .Q(\fifo_bank_register.bank[5][118] ));
 sky130_fd_sc_hd__dfxtp_1 _17341_ (.CLK(net429),
    .D(_00784_),
    .Q(\fifo_bank_register.bank[5][119] ));
 sky130_fd_sc_hd__dfxtp_1 _17342_ (.CLK(net441),
    .D(_00785_),
    .Q(\fifo_bank_register.bank[5][120] ));
 sky130_fd_sc_hd__dfxtp_1 _17343_ (.CLK(net490),
    .D(_00786_),
    .Q(\fifo_bank_register.bank[5][121] ));
 sky130_fd_sc_hd__dfxtp_1 _17344_ (.CLK(net492),
    .D(_00787_),
    .Q(\fifo_bank_register.bank[5][122] ));
 sky130_fd_sc_hd__dfxtp_1 _17345_ (.CLK(net439),
    .D(_00788_),
    .Q(\fifo_bank_register.bank[5][123] ));
 sky130_fd_sc_hd__dfxtp_1 _17346_ (.CLK(net494),
    .D(_00789_),
    .Q(\fifo_bank_register.bank[5][124] ));
 sky130_fd_sc_hd__dfxtp_1 _17347_ (.CLK(net494),
    .D(_00790_),
    .Q(\fifo_bank_register.bank[5][125] ));
 sky130_fd_sc_hd__dfxtp_1 _17348_ (.CLK(net494),
    .D(_00791_),
    .Q(\fifo_bank_register.bank[5][126] ));
 sky130_fd_sc_hd__dfxtp_1 _17349_ (.CLK(net441),
    .D(_00792_),
    .Q(\fifo_bank_register.bank[5][127] ));
 sky130_fd_sc_hd__dfxtp_1 _17350_ (.CLK(net473),
    .D(_00793_),
    .Q(\fifo_bank_register.bank[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17351_ (.CLK(net490),
    .D(_00794_),
    .Q(\fifo_bank_register.bank[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17352_ (.CLK(net474),
    .D(_00795_),
    .Q(\fifo_bank_register.bank[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17353_ (.CLK(net473),
    .D(_00796_),
    .Q(\fifo_bank_register.bank[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17354_ (.CLK(net474),
    .D(_00797_),
    .Q(\fifo_bank_register.bank[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17355_ (.CLK(net474),
    .D(_00798_),
    .Q(\fifo_bank_register.bank[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17356_ (.CLK(net477),
    .D(_00799_),
    .Q(\fifo_bank_register.bank[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17357_ (.CLK(net477),
    .D(_00800_),
    .Q(\fifo_bank_register.bank[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17358_ (.CLK(net478),
    .D(_00801_),
    .Q(\fifo_bank_register.bank[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17359_ (.CLK(net478),
    .D(_00802_),
    .Q(\fifo_bank_register.bank[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17360_ (.CLK(net496),
    .D(_00803_),
    .Q(\fifo_bank_register.bank[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17361_ (.CLK(net533),
    .D(_00804_),
    .Q(\fifo_bank_register.bank[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17362_ (.CLK(net504),
    .D(_00805_),
    .Q(\fifo_bank_register.bank[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17363_ (.CLK(net505),
    .D(_00806_),
    .Q(\fifo_bank_register.bank[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17364_ (.CLK(net534),
    .D(_00807_),
    .Q(\fifo_bank_register.bank[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17365_ (.CLK(net534),
    .D(_00808_),
    .Q(\fifo_bank_register.bank[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17366_ (.CLK(net496),
    .D(_00809_),
    .Q(\fifo_bank_register.bank[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17367_ (.CLK(net532),
    .D(_00810_),
    .Q(\fifo_bank_register.bank[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17368_ (.CLK(net533),
    .D(_00811_),
    .Q(\fifo_bank_register.bank[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17369_ (.CLK(net505),
    .D(_00812_),
    .Q(\fifo_bank_register.bank[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17370_ (.CLK(net501),
    .D(_00813_),
    .Q(\fifo_bank_register.bank[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17371_ (.CLK(net482),
    .D(_00814_),
    .Q(\fifo_bank_register.bank[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17372_ (.CLK(net500),
    .D(_00815_),
    .Q(\fifo_bank_register.bank[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17373_ (.CLK(net484),
    .D(_00816_),
    .Q(\fifo_bank_register.bank[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17374_ (.CLK(net485),
    .D(_00817_),
    .Q(\fifo_bank_register.bank[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17375_ (.CLK(net509),
    .D(_00818_),
    .Q(\fifo_bank_register.bank[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17376_ (.CLK(net483),
    .D(_00819_),
    .Q(\fifo_bank_register.bank[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17377_ (.CLK(net499),
    .D(_00820_),
    .Q(\fifo_bank_register.bank[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17378_ (.CLK(net485),
    .D(_00821_),
    .Q(\fifo_bank_register.bank[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17379_ (.CLK(net500),
    .D(_00822_),
    .Q(\fifo_bank_register.bank[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17380_ (.CLK(net430),
    .D(_00823_),
    .Q(\fifo_bank_register.bank[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17381_ (.CLK(net437),
    .D(_00824_),
    .Q(\fifo_bank_register.bank[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17382_ (.CLK(net417),
    .D(_00825_),
    .Q(\fifo_bank_register.bank[4][32] ));
 sky130_fd_sc_hd__dfxtp_1 _17383_ (.CLK(net423),
    .D(_00826_),
    .Q(\fifo_bank_register.bank[4][33] ));
 sky130_fd_sc_hd__dfxtp_1 _17384_ (.CLK(net430),
    .D(_00827_),
    .Q(\fifo_bank_register.bank[4][34] ));
 sky130_fd_sc_hd__dfxtp_1 _17385_ (.CLK(net428),
    .D(_00828_),
    .Q(\fifo_bank_register.bank[4][35] ));
 sky130_fd_sc_hd__dfxtp_1 _17386_ (.CLK(net422),
    .D(_00829_),
    .Q(\fifo_bank_register.bank[4][36] ));
 sky130_fd_sc_hd__dfxtp_1 _17387_ (.CLK(net417),
    .D(_00830_),
    .Q(\fifo_bank_register.bank[4][37] ));
 sky130_fd_sc_hd__dfxtp_1 _17388_ (.CLK(net428),
    .D(_00831_),
    .Q(\fifo_bank_register.bank[4][38] ));
 sky130_fd_sc_hd__dfxtp_1 _17389_ (.CLK(net415),
    .D(_00832_),
    .Q(\fifo_bank_register.bank[4][39] ));
 sky130_fd_sc_hd__dfxtp_1 _17390_ (.CLK(net395),
    .D(_00833_),
    .Q(\fifo_bank_register.bank[4][40] ));
 sky130_fd_sc_hd__dfxtp_1 _17391_ (.CLK(net398),
    .D(_00834_),
    .Q(\fifo_bank_register.bank[4][41] ));
 sky130_fd_sc_hd__dfxtp_1 _17392_ (.CLK(net398),
    .D(_00835_),
    .Q(\fifo_bank_register.bank[4][42] ));
 sky130_fd_sc_hd__dfxtp_1 _17393_ (.CLK(net393),
    .D(_00836_),
    .Q(\fifo_bank_register.bank[4][43] ));
 sky130_fd_sc_hd__dfxtp_1 _17394_ (.CLK(net389),
    .D(_00837_),
    .Q(\fifo_bank_register.bank[4][44] ));
 sky130_fd_sc_hd__dfxtp_1 _17395_ (.CLK(net406),
    .D(_00838_),
    .Q(\fifo_bank_register.bank[4][45] ));
 sky130_fd_sc_hd__dfxtp_1 _17396_ (.CLK(net390),
    .D(_00839_),
    .Q(\fifo_bank_register.bank[4][46] ));
 sky130_fd_sc_hd__dfxtp_1 _17397_ (.CLK(net395),
    .D(_00840_),
    .Q(\fifo_bank_register.bank[4][47] ));
 sky130_fd_sc_hd__dfxtp_1 _17398_ (.CLK(net395),
    .D(_00841_),
    .Q(\fifo_bank_register.bank[4][48] ));
 sky130_fd_sc_hd__dfxtp_1 _17399_ (.CLK(net408),
    .D(_00842_),
    .Q(\fifo_bank_register.bank[4][49] ));
 sky130_fd_sc_hd__dfxtp_1 _17400_ (.CLK(net572),
    .D(_00843_),
    .Q(\fifo_bank_register.bank[4][50] ));
 sky130_fd_sc_hd__dfxtp_1 _17401_ (.CLK(net575),
    .D(_00844_),
    .Q(\fifo_bank_register.bank[4][51] ));
 sky130_fd_sc_hd__dfxtp_1 _17402_ (.CLK(net567),
    .D(_00845_),
    .Q(\fifo_bank_register.bank[4][52] ));
 sky130_fd_sc_hd__dfxtp_1 _17403_ (.CLK(net567),
    .D(_00846_),
    .Q(\fifo_bank_register.bank[4][53] ));
 sky130_fd_sc_hd__dfxtp_1 _17404_ (.CLK(net556),
    .D(_00847_),
    .Q(\fifo_bank_register.bank[4][54] ));
 sky130_fd_sc_hd__dfxtp_1 _17405_ (.CLK(net574),
    .D(_00848_),
    .Q(\fifo_bank_register.bank[4][55] ));
 sky130_fd_sc_hd__dfxtp_1 _17406_ (.CLK(net574),
    .D(_00849_),
    .Q(\fifo_bank_register.bank[4][56] ));
 sky130_fd_sc_hd__dfxtp_1 _17407_ (.CLK(net550),
    .D(_00850_),
    .Q(\fifo_bank_register.bank[4][57] ));
 sky130_fd_sc_hd__dfxtp_1 _17408_ (.CLK(net558),
    .D(_00851_),
    .Q(\fifo_bank_register.bank[4][58] ));
 sky130_fd_sc_hd__dfxtp_1 _17409_ (.CLK(net573),
    .D(_00852_),
    .Q(\fifo_bank_register.bank[4][59] ));
 sky130_fd_sc_hd__dfxtp_1 _17410_ (.CLK(net515),
    .D(_00853_),
    .Q(\fifo_bank_register.bank[4][60] ));
 sky130_fd_sc_hd__dfxtp_1 _17411_ (.CLK(net524),
    .D(_00854_),
    .Q(\fifo_bank_register.bank[4][61] ));
 sky130_fd_sc_hd__dfxtp_1 _17412_ (.CLK(net523),
    .D(_00855_),
    .Q(\fifo_bank_register.bank[4][62] ));
 sky130_fd_sc_hd__dfxtp_1 _17413_ (.CLK(net523),
    .D(_00856_),
    .Q(\fifo_bank_register.bank[4][63] ));
 sky130_fd_sc_hd__dfxtp_1 _17414_ (.CLK(net514),
    .D(_00857_),
    .Q(\fifo_bank_register.bank[4][64] ));
 sky130_fd_sc_hd__dfxtp_1 _17415_ (.CLK(net518),
    .D(_00858_),
    .Q(\fifo_bank_register.bank[4][65] ));
 sky130_fd_sc_hd__dfxtp_1 _17416_ (.CLK(net524),
    .D(_00859_),
    .Q(\fifo_bank_register.bank[4][66] ));
 sky130_fd_sc_hd__dfxtp_1 _17417_ (.CLK(net514),
    .D(_00860_),
    .Q(\fifo_bank_register.bank[4][67] ));
 sky130_fd_sc_hd__dfxtp_1 _17418_ (.CLK(net521),
    .D(_00861_),
    .Q(\fifo_bank_register.bank[4][68] ));
 sky130_fd_sc_hd__dfxtp_1 _17419_ (.CLK(net518),
    .D(_00862_),
    .Q(\fifo_bank_register.bank[4][69] ));
 sky130_fd_sc_hd__dfxtp_1 _17420_ (.CLK(net519),
    .D(_00863_),
    .Q(\fifo_bank_register.bank[4][70] ));
 sky130_fd_sc_hd__dfxtp_1 _17421_ (.CLK(net525),
    .D(_00864_),
    .Q(\fifo_bank_register.bank[4][71] ));
 sky130_fd_sc_hd__dfxtp_1 _17422_ (.CLK(net553),
    .D(_00865_),
    .Q(\fifo_bank_register.bank[4][72] ));
 sky130_fd_sc_hd__dfxtp_1 _17423_ (.CLK(net552),
    .D(_00866_),
    .Q(\fifo_bank_register.bank[4][73] ));
 sky130_fd_sc_hd__dfxtp_1 _17424_ (.CLK(net546),
    .D(_00867_),
    .Q(\fifo_bank_register.bank[4][74] ));
 sky130_fd_sc_hd__dfxtp_1 _17425_ (.CLK(net552),
    .D(_00868_),
    .Q(\fifo_bank_register.bank[4][75] ));
 sky130_fd_sc_hd__dfxtp_1 _17426_ (.CLK(net545),
    .D(_00869_),
    .Q(\fifo_bank_register.bank[4][76] ));
 sky130_fd_sc_hd__dfxtp_1 _17427_ (.CLK(net552),
    .D(_00870_),
    .Q(\fifo_bank_register.bank[4][77] ));
 sky130_fd_sc_hd__dfxtp_1 _17428_ (.CLK(net525),
    .D(_00871_),
    .Q(\fifo_bank_register.bank[4][78] ));
 sky130_fd_sc_hd__dfxtp_1 _17429_ (.CLK(net553),
    .D(_00872_),
    .Q(\fifo_bank_register.bank[4][79] ));
 sky130_fd_sc_hd__dfxtp_1 _17430_ (.CLK(net565),
    .D(_00873_),
    .Q(\fifo_bank_register.bank[4][80] ));
 sky130_fd_sc_hd__dfxtp_1 _17431_ (.CLK(net565),
    .D(_00874_),
    .Q(\fifo_bank_register.bank[4][81] ));
 sky130_fd_sc_hd__dfxtp_1 _17432_ (.CLK(net560),
    .D(_00875_),
    .Q(\fifo_bank_register.bank[4][82] ));
 sky130_fd_sc_hd__dfxtp_1 _17433_ (.CLK(net560),
    .D(_00876_),
    .Q(\fifo_bank_register.bank[4][83] ));
 sky130_fd_sc_hd__dfxtp_1 _17434_ (.CLK(net548),
    .D(_00877_),
    .Q(\fifo_bank_register.bank[4][84] ));
 sky130_fd_sc_hd__dfxtp_1 _17435_ (.CLK(net565),
    .D(_00878_),
    .Q(\fifo_bank_register.bank[4][85] ));
 sky130_fd_sc_hd__dfxtp_1 _17436_ (.CLK(net560),
    .D(_00879_),
    .Q(\fifo_bank_register.bank[4][86] ));
 sky130_fd_sc_hd__dfxtp_1 _17437_ (.CLK(net560),
    .D(_00880_),
    .Q(\fifo_bank_register.bank[4][87] ));
 sky130_fd_sc_hd__dfxtp_1 _17438_ (.CLK(net565),
    .D(_00881_),
    .Q(\fifo_bank_register.bank[4][88] ));
 sky130_fd_sc_hd__dfxtp_1 _17439_ (.CLK(net548),
    .D(_00882_),
    .Q(\fifo_bank_register.bank[4][89] ));
 sky130_fd_sc_hd__dfxtp_1 _17440_ (.CLK(net409),
    .D(_00883_),
    .Q(\fifo_bank_register.bank[4][90] ));
 sky130_fd_sc_hd__dfxtp_1 _17441_ (.CLK(net401),
    .D(_00884_),
    .Q(\fifo_bank_register.bank[4][91] ));
 sky130_fd_sc_hd__dfxtp_1 _17442_ (.CLK(net410),
    .D(_00885_),
    .Q(\fifo_bank_register.bank[4][92] ));
 sky130_fd_sc_hd__dfxtp_1 _17443_ (.CLK(net400),
    .D(_00886_),
    .Q(\fifo_bank_register.bank[4][93] ));
 sky130_fd_sc_hd__dfxtp_1 _17444_ (.CLK(net455),
    .D(_00887_),
    .Q(\fifo_bank_register.bank[4][94] ));
 sky130_fd_sc_hd__dfxtp_1 _17445_ (.CLK(net402),
    .D(_00888_),
    .Q(\fifo_bank_register.bank[4][95] ));
 sky130_fd_sc_hd__dfxtp_1 _17446_ (.CLK(net448),
    .D(_00889_),
    .Q(\fifo_bank_register.bank[4][96] ));
 sky130_fd_sc_hd__dfxtp_1 _17447_ (.CLK(net454),
    .D(_00890_),
    .Q(\fifo_bank_register.bank[4][97] ));
 sky130_fd_sc_hd__dfxtp_1 _17448_ (.CLK(net447),
    .D(_00891_),
    .Q(\fifo_bank_register.bank[4][98] ));
 sky130_fd_sc_hd__dfxtp_1 _17449_ (.CLK(net445),
    .D(_00892_),
    .Q(\fifo_bank_register.bank[4][99] ));
 sky130_fd_sc_hd__dfxtp_1 _17450_ (.CLK(net453),
    .D(_00893_),
    .Q(\fifo_bank_register.bank[4][100] ));
 sky130_fd_sc_hd__dfxtp_1 _17451_ (.CLK(net451),
    .D(_00894_),
    .Q(\fifo_bank_register.bank[4][101] ));
 sky130_fd_sc_hd__dfxtp_1 _17452_ (.CLK(net465),
    .D(_00895_),
    .Q(\fifo_bank_register.bank[4][102] ));
 sky130_fd_sc_hd__dfxtp_1 _17453_ (.CLK(net467),
    .D(_00896_),
    .Q(\fifo_bank_register.bank[4][103] ));
 sky130_fd_sc_hd__dfxtp_1 _17454_ (.CLK(net462),
    .D(_00897_),
    .Q(\fifo_bank_register.bank[4][104] ));
 sky130_fd_sc_hd__dfxtp_1 _17455_ (.CLK(net467),
    .D(_00898_),
    .Q(\fifo_bank_register.bank[4][105] ));
 sky130_fd_sc_hd__dfxtp_1 _17456_ (.CLK(net465),
    .D(_00899_),
    .Q(\fifo_bank_register.bank[4][106] ));
 sky130_fd_sc_hd__dfxtp_1 _17457_ (.CLK(net451),
    .D(_00900_),
    .Q(\fifo_bank_register.bank[4][107] ));
 sky130_fd_sc_hd__dfxtp_1 _17458_ (.CLK(net452),
    .D(_00901_),
    .Q(\fifo_bank_register.bank[4][108] ));
 sky130_fd_sc_hd__dfxtp_1 _17459_ (.CLK(net459),
    .D(_00902_),
    .Q(\fifo_bank_register.bank[4][109] ));
 sky130_fd_sc_hd__dfxtp_1 _17460_ (.CLK(net434),
    .D(_00903_),
    .Q(\fifo_bank_register.bank[4][110] ));
 sky130_fd_sc_hd__dfxtp_1 _17461_ (.CLK(net411),
    .D(_00904_),
    .Q(\fifo_bank_register.bank[4][111] ));
 sky130_fd_sc_hd__dfxtp_1 _17462_ (.CLK(net411),
    .D(_00905_),
    .Q(\fifo_bank_register.bank[4][112] ));
 sky130_fd_sc_hd__dfxtp_1 _17463_ (.CLK(net469),
    .D(_00906_),
    .Q(\fifo_bank_register.bank[4][113] ));
 sky130_fd_sc_hd__dfxtp_1 _17464_ (.CLK(net456),
    .D(_00907_),
    .Q(\fifo_bank_register.bank[4][114] ));
 sky130_fd_sc_hd__dfxtp_1 _17465_ (.CLK(net470),
    .D(_00908_),
    .Q(\fifo_bank_register.bank[4][115] ));
 sky130_fd_sc_hd__dfxtp_1 _17466_ (.CLK(net411),
    .D(_00909_),
    .Q(\fifo_bank_register.bank[4][116] ));
 sky130_fd_sc_hd__dfxtp_1 _17467_ (.CLK(net435),
    .D(_00910_),
    .Q(\fifo_bank_register.bank[4][117] ));
 sky130_fd_sc_hd__dfxtp_1 _17468_ (.CLK(net456),
    .D(_00911_),
    .Q(\fifo_bank_register.bank[4][118] ));
 sky130_fd_sc_hd__dfxtp_1 _17469_ (.CLK(net435),
    .D(_00912_),
    .Q(\fifo_bank_register.bank[4][119] ));
 sky130_fd_sc_hd__dfxtp_1 _17470_ (.CLK(net442),
    .D(_00913_),
    .Q(\fifo_bank_register.bank[4][120] ));
 sky130_fd_sc_hd__dfxtp_1 _17471_ (.CLK(net440),
    .D(_00914_),
    .Q(\fifo_bank_register.bank[4][121] ));
 sky130_fd_sc_hd__dfxtp_1 _17472_ (.CLK(net490),
    .D(_00915_),
    .Q(\fifo_bank_register.bank[4][122] ));
 sky130_fd_sc_hd__dfxtp_1 _17473_ (.CLK(net439),
    .D(_00916_),
    .Q(\fifo_bank_register.bank[4][123] ));
 sky130_fd_sc_hd__dfxtp_1 _17474_ (.CLK(net495),
    .D(_00917_),
    .Q(\fifo_bank_register.bank[4][124] ));
 sky130_fd_sc_hd__dfxtp_1 _17475_ (.CLK(net495),
    .D(_00918_),
    .Q(\fifo_bank_register.bank[4][125] ));
 sky130_fd_sc_hd__dfxtp_1 _17476_ (.CLK(net495),
    .D(_00919_),
    .Q(\fifo_bank_register.bank[4][126] ));
 sky130_fd_sc_hd__dfxtp_1 _17477_ (.CLK(net443),
    .D(_00920_),
    .Q(\fifo_bank_register.bank[4][127] ));
 sky130_fd_sc_hd__dfxtp_1 _17478_ (.CLK(net475),
    .D(_00921_),
    .Q(\fifo_bank_register.bank[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17479_ (.CLK(net492),
    .D(_00922_),
    .Q(\fifo_bank_register.bank[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17480_ (.CLK(net476),
    .D(_00923_),
    .Q(\fifo_bank_register.bank[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17481_ (.CLK(net475),
    .D(_00924_),
    .Q(\fifo_bank_register.bank[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17482_ (.CLK(net474),
    .D(_00925_),
    .Q(\fifo_bank_register.bank[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17483_ (.CLK(net476),
    .D(_00926_),
    .Q(\fifo_bank_register.bank[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17484_ (.CLK(net479),
    .D(_00927_),
    .Q(\fifo_bank_register.bank[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17485_ (.CLK(net479),
    .D(_00928_),
    .Q(\fifo_bank_register.bank[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17486_ (.CLK(net492),
    .D(_00929_),
    .Q(\fifo_bank_register.bank[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17487_ (.CLK(net480),
    .D(_00930_),
    .Q(\fifo_bank_register.bank[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17488_ (.CLK(net493),
    .D(_00931_),
    .Q(\fifo_bank_register.bank[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17489_ (.CLK(net503),
    .D(_00932_),
    .Q(\fifo_bank_register.bank[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17490_ (.CLK(net500),
    .D(_00933_),
    .Q(\fifo_bank_register.bank[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17491_ (.CLK(net507),
    .D(_00934_),
    .Q(\fifo_bank_register.bank[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17492_ (.CLK(net503),
    .D(_00935_),
    .Q(\fifo_bank_register.bank[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17493_ (.CLK(net503),
    .D(_00936_),
    .Q(\fifo_bank_register.bank[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17494_ (.CLK(net492),
    .D(_00937_),
    .Q(\fifo_bank_register.bank[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17495_ (.CLK(net497),
    .D(_00938_),
    .Q(\fifo_bank_register.bank[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17496_ (.CLK(net497),
    .D(_00939_),
    .Q(\fifo_bank_register.bank[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17497_ (.CLK(net502),
    .D(_00940_),
    .Q(\fifo_bank_register.bank[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17498_ (.CLK(net501),
    .D(_00941_),
    .Q(\fifo_bank_register.bank[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17499_ (.CLK(net485),
    .D(_00942_),
    .Q(\fifo_bank_register.bank[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17500_ (.CLK(net488),
    .D(_00943_),
    .Q(\fifo_bank_register.bank[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17501_ (.CLK(net487),
    .D(_00944_),
    .Q(\fifo_bank_register.bank[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17502_ (.CLK(net485),
    .D(_00945_),
    .Q(\fifo_bank_register.bank[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17503_ (.CLK(net487),
    .D(_00946_),
    .Q(\fifo_bank_register.bank[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17504_ (.CLK(net487),
    .D(_00947_),
    .Q(\fifo_bank_register.bank[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17505_ (.CLK(net488),
    .D(_00948_),
    .Q(\fifo_bank_register.bank[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17506_ (.CLK(net487),
    .D(_00949_),
    .Q(\fifo_bank_register.bank[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17507_ (.CLK(net499),
    .D(_00950_),
    .Q(\fifo_bank_register.bank[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17508_ (.CLK(net418),
    .D(_00951_),
    .Q(\fifo_bank_register.bank[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17509_ (.CLK(net424),
    .D(_00952_),
    .Q(\fifo_bank_register.bank[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17510_ (.CLK(net419),
    .D(_00953_),
    .Q(\fifo_bank_register.bank[3][32] ));
 sky130_fd_sc_hd__dfxtp_1 _17511_ (.CLK(net424),
    .D(_00954_),
    .Q(\fifo_bank_register.bank[3][33] ));
 sky130_fd_sc_hd__dfxtp_1 _17512_ (.CLK(net418),
    .D(_00955_),
    .Q(\fifo_bank_register.bank[3][34] ));
 sky130_fd_sc_hd__dfxtp_1 _17513_ (.CLK(net416),
    .D(_00956_),
    .Q(\fifo_bank_register.bank[3][35] ));
 sky130_fd_sc_hd__dfxtp_1 _17514_ (.CLK(net422),
    .D(_00957_),
    .Q(\fifo_bank_register.bank[3][36] ));
 sky130_fd_sc_hd__dfxtp_1 _17515_ (.CLK(net414),
    .D(_00958_),
    .Q(\fifo_bank_register.bank[3][37] ));
 sky130_fd_sc_hd__dfxtp_1 _17516_ (.CLK(net416),
    .D(_00959_),
    .Q(\fifo_bank_register.bank[3][38] ));
 sky130_fd_sc_hd__dfxtp_1 _17517_ (.CLK(net414),
    .D(_00960_),
    .Q(\fifo_bank_register.bank[3][39] ));
 sky130_fd_sc_hd__dfxtp_1 _17518_ (.CLK(net392),
    .D(_00961_),
    .Q(\fifo_bank_register.bank[3][40] ));
 sky130_fd_sc_hd__dfxtp_1 _17519_ (.CLK(net398),
    .D(_00962_),
    .Q(\fifo_bank_register.bank[3][41] ));
 sky130_fd_sc_hd__dfxtp_1 _17520_ (.CLK(net389),
    .D(_00963_),
    .Q(\fifo_bank_register.bank[3][42] ));
 sky130_fd_sc_hd__dfxtp_1 _17521_ (.CLK(net392),
    .D(_00964_),
    .Q(\fifo_bank_register.bank[3][43] ));
 sky130_fd_sc_hd__dfxtp_1 _17522_ (.CLK(net391),
    .D(_00965_),
    .Q(\fifo_bank_register.bank[3][44] ));
 sky130_fd_sc_hd__dfxtp_1 _17523_ (.CLK(net394),
    .D(_00966_),
    .Q(\fifo_bank_register.bank[3][45] ));
 sky130_fd_sc_hd__dfxtp_1 _17524_ (.CLK(net391),
    .D(_00967_),
    .Q(\fifo_bank_register.bank[3][46] ));
 sky130_fd_sc_hd__dfxtp_1 _17525_ (.CLK(net394),
    .D(_00968_),
    .Q(\fifo_bank_register.bank[3][47] ));
 sky130_fd_sc_hd__dfxtp_1 _17526_ (.CLK(net392),
    .D(_00969_),
    .Q(\fifo_bank_register.bank[3][48] ));
 sky130_fd_sc_hd__dfxtp_1 _17527_ (.CLK(net405),
    .D(_00970_),
    .Q(\fifo_bank_register.bank[3][49] ));
 sky130_fd_sc_hd__dfxtp_1 _17528_ (.CLK(net556),
    .D(_00971_),
    .Q(\fifo_bank_register.bank[3][50] ));
 sky130_fd_sc_hd__dfxtp_1 _17529_ (.CLK(net570),
    .D(_00972_),
    .Q(\fifo_bank_register.bank[3][51] ));
 sky130_fd_sc_hd__dfxtp_1 _17530_ (.CLK(net562),
    .D(_00973_),
    .Q(\fifo_bank_register.bank[3][52] ));
 sky130_fd_sc_hd__dfxtp_1 _17531_ (.CLK(net562),
    .D(_00974_),
    .Q(\fifo_bank_register.bank[3][53] ));
 sky130_fd_sc_hd__dfxtp_1 _17532_ (.CLK(net556),
    .D(_00975_),
    .Q(\fifo_bank_register.bank[3][54] ));
 sky130_fd_sc_hd__dfxtp_1 _17533_ (.CLK(net570),
    .D(_00976_),
    .Q(\fifo_bank_register.bank[3][55] ));
 sky130_fd_sc_hd__dfxtp_1 _17534_ (.CLK(net570),
    .D(_00977_),
    .Q(\fifo_bank_register.bank[3][56] ));
 sky130_fd_sc_hd__dfxtp_1 _17535_ (.CLK(net550),
    .D(_00978_),
    .Q(\fifo_bank_register.bank[3][57] ));
 sky130_fd_sc_hd__dfxtp_1 _17536_ (.CLK(net556),
    .D(_00979_),
    .Q(\fifo_bank_register.bank[3][58] ));
 sky130_fd_sc_hd__dfxtp_1 _17537_ (.CLK(net570),
    .D(_00980_),
    .Q(\fifo_bank_register.bank[3][59] ));
 sky130_fd_sc_hd__dfxtp_1 _17538_ (.CLK(net513),
    .D(_00981_),
    .Q(\fifo_bank_register.bank[3][60] ));
 sky130_fd_sc_hd__dfxtp_1 _17539_ (.CLK(net526),
    .D(_00982_),
    .Q(\fifo_bank_register.bank[3][61] ));
 sky130_fd_sc_hd__dfxtp_1 _17540_ (.CLK(net521),
    .D(_00983_),
    .Q(\fifo_bank_register.bank[3][62] ));
 sky130_fd_sc_hd__dfxtp_1 _17541_ (.CLK(net522),
    .D(_00984_),
    .Q(\fifo_bank_register.bank[3][63] ));
 sky130_fd_sc_hd__dfxtp_1 _17542_ (.CLK(net512),
    .D(_00985_),
    .Q(\fifo_bank_register.bank[3][64] ));
 sky130_fd_sc_hd__dfxtp_1 _17543_ (.CLK(net521),
    .D(_00986_),
    .Q(\fifo_bank_register.bank[3][65] ));
 sky130_fd_sc_hd__dfxtp_1 _17544_ (.CLK(net522),
    .D(_00987_),
    .Q(\fifo_bank_register.bank[3][66] ));
 sky130_fd_sc_hd__dfxtp_1 _17545_ (.CLK(net515),
    .D(_00988_),
    .Q(\fifo_bank_register.bank[3][67] ));
 sky130_fd_sc_hd__dfxtp_1 _17546_ (.CLK(net522),
    .D(_00989_),
    .Q(\fifo_bank_register.bank[3][68] ));
 sky130_fd_sc_hd__dfxtp_1 _17547_ (.CLK(net513),
    .D(_00990_),
    .Q(\fifo_bank_register.bank[3][69] ));
 sky130_fd_sc_hd__dfxtp_1 _17548_ (.CLK(net517),
    .D(_00991_),
    .Q(\fifo_bank_register.bank[3][70] ));
 sky130_fd_sc_hd__dfxtp_1 _17549_ (.CLK(net517),
    .D(_00992_),
    .Q(\fifo_bank_register.bank[3][71] ));
 sky130_fd_sc_hd__dfxtp_1 _17550_ (.CLK(net544),
    .D(_00993_),
    .Q(\fifo_bank_register.bank[3][72] ));
 sky130_fd_sc_hd__dfxtp_1 _17551_ (.CLK(net543),
    .D(_00994_),
    .Q(\fifo_bank_register.bank[3][73] ));
 sky130_fd_sc_hd__dfxtp_1 _17552_ (.CLK(net547),
    .D(_00995_),
    .Q(\fifo_bank_register.bank[3][74] ));
 sky130_fd_sc_hd__dfxtp_1 _17553_ (.CLK(net543),
    .D(_00996_),
    .Q(\fifo_bank_register.bank[3][75] ));
 sky130_fd_sc_hd__dfxtp_1 _17554_ (.CLK(net543),
    .D(_00997_),
    .Q(\fifo_bank_register.bank[3][76] ));
 sky130_fd_sc_hd__dfxtp_1 _17555_ (.CLK(net544),
    .D(_00998_),
    .Q(\fifo_bank_register.bank[3][77] ));
 sky130_fd_sc_hd__dfxtp_1 _17556_ (.CLK(net517),
    .D(_00999_),
    .Q(\fifo_bank_register.bank[3][78] ));
 sky130_fd_sc_hd__dfxtp_1 _17557_ (.CLK(net547),
    .D(_01000_),
    .Q(\fifo_bank_register.bank[3][79] ));
 sky130_fd_sc_hd__dfxtp_1 _17558_ (.CLK(net540),
    .D(_01001_),
    .Q(\fifo_bank_register.bank[3][80] ));
 sky130_fd_sc_hd__dfxtp_1 _17559_ (.CLK(net540),
    .D(_01002_),
    .Q(\fifo_bank_register.bank[3][81] ));
 sky130_fd_sc_hd__dfxtp_1 _17560_ (.CLK(net538),
    .D(_01003_),
    .Q(\fifo_bank_register.bank[3][82] ));
 sky130_fd_sc_hd__dfxtp_1 _17561_ (.CLK(net538),
    .D(_01004_),
    .Q(\fifo_bank_register.bank[3][83] ));
 sky130_fd_sc_hd__dfxtp_1 _17562_ (.CLK(net537),
    .D(_01005_),
    .Q(\fifo_bank_register.bank[3][84] ));
 sky130_fd_sc_hd__dfxtp_1 _17563_ (.CLK(net540),
    .D(_01006_),
    .Q(\fifo_bank_register.bank[3][85] ));
 sky130_fd_sc_hd__dfxtp_1 _17564_ (.CLK(net538),
    .D(_01007_),
    .Q(\fifo_bank_register.bank[3][86] ));
 sky130_fd_sc_hd__dfxtp_1 _17565_ (.CLK(net538),
    .D(_01008_),
    .Q(\fifo_bank_register.bank[3][87] ));
 sky130_fd_sc_hd__dfxtp_1 _17566_ (.CLK(net540),
    .D(_01009_),
    .Q(\fifo_bank_register.bank[3][88] ));
 sky130_fd_sc_hd__dfxtp_1 _17567_ (.CLK(net536),
    .D(_01010_),
    .Q(\fifo_bank_register.bank[3][89] ));
 sky130_fd_sc_hd__dfxtp_1 _17568_ (.CLK(net402),
    .D(_01011_),
    .Q(\fifo_bank_register.bank[3][90] ));
 sky130_fd_sc_hd__dfxtp_1 _17569_ (.CLK(net401),
    .D(_01012_),
    .Q(\fifo_bank_register.bank[3][91] ));
 sky130_fd_sc_hd__dfxtp_1 _17570_ (.CLK(net403),
    .D(_01013_),
    .Q(\fifo_bank_register.bank[3][92] ));
 sky130_fd_sc_hd__dfxtp_1 _17571_ (.CLK(net400),
    .D(_01014_),
    .Q(\fifo_bank_register.bank[3][93] ));
 sky130_fd_sc_hd__dfxtp_1 _17572_ (.CLK(net448),
    .D(_01015_),
    .Q(\fifo_bank_register.bank[3][94] ));
 sky130_fd_sc_hd__dfxtp_1 _17573_ (.CLK(net400),
    .D(_01016_),
    .Q(\fifo_bank_register.bank[3][95] ));
 sky130_fd_sc_hd__dfxtp_1 _17574_ (.CLK(net445),
    .D(_01017_),
    .Q(\fifo_bank_register.bank[3][96] ));
 sky130_fd_sc_hd__dfxtp_1 _17575_ (.CLK(net448),
    .D(_01018_),
    .Q(\fifo_bank_register.bank[3][97] ));
 sky130_fd_sc_hd__dfxtp_1 _17576_ (.CLK(net445),
    .D(_01019_),
    .Q(\fifo_bank_register.bank[3][98] ));
 sky130_fd_sc_hd__dfxtp_1 _17577_ (.CLK(net445),
    .D(_01020_),
    .Q(\fifo_bank_register.bank[3][99] ));
 sky130_fd_sc_hd__dfxtp_1 _17578_ (.CLK(net447),
    .D(_01021_),
    .Q(\fifo_bank_register.bank[3][100] ));
 sky130_fd_sc_hd__dfxtp_1 _17579_ (.CLK(net450),
    .D(_01022_),
    .Q(\fifo_bank_register.bank[3][101] ));
 sky130_fd_sc_hd__dfxtp_1 _17580_ (.CLK(net464),
    .D(_01023_),
    .Q(\fifo_bank_register.bank[3][102] ));
 sky130_fd_sc_hd__dfxtp_1 _17581_ (.CLK(net464),
    .D(_01024_),
    .Q(\fifo_bank_register.bank[3][103] ));
 sky130_fd_sc_hd__dfxtp_1 _17582_ (.CLK(net462),
    .D(_01025_),
    .Q(\fifo_bank_register.bank[3][104] ));
 sky130_fd_sc_hd__dfxtp_1 _17583_ (.CLK(net464),
    .D(_01026_),
    .Q(\fifo_bank_register.bank[3][105] ));
 sky130_fd_sc_hd__dfxtp_1 _17584_ (.CLK(net462),
    .D(_01027_),
    .Q(\fifo_bank_register.bank[3][106] ));
 sky130_fd_sc_hd__dfxtp_1 _17585_ (.CLK(net462),
    .D(_01028_),
    .Q(\fifo_bank_register.bank[3][107] ));
 sky130_fd_sc_hd__dfxtp_1 _17586_ (.CLK(net451),
    .D(_01029_),
    .Q(\fifo_bank_register.bank[3][108] ));
 sky130_fd_sc_hd__dfxtp_1 _17587_ (.CLK(net458),
    .D(_01030_),
    .Q(\fifo_bank_register.bank[3][109] ));
 sky130_fd_sc_hd__dfxtp_1 _17588_ (.CLK(net432),
    .D(_01031_),
    .Q(\fifo_bank_register.bank[3][110] ));
 sky130_fd_sc_hd__dfxtp_1 _17589_ (.CLK(net409),
    .D(_01032_),
    .Q(\fifo_bank_register.bank[3][111] ));
 sky130_fd_sc_hd__dfxtp_1 _17590_ (.CLK(net412),
    .D(_01033_),
    .Q(\fifo_bank_register.bank[3][112] ));
 sky130_fd_sc_hd__dfxtp_1 _17591_ (.CLK(net429),
    .D(_01034_),
    .Q(\fifo_bank_register.bank[3][113] ));
 sky130_fd_sc_hd__dfxtp_1 _17592_ (.CLK(net408),
    .D(_01035_),
    .Q(\fifo_bank_register.bank[3][114] ));
 sky130_fd_sc_hd__dfxtp_1 _17593_ (.CLK(net432),
    .D(_01036_),
    .Q(\fifo_bank_register.bank[3][115] ));
 sky130_fd_sc_hd__dfxtp_1 _17594_ (.CLK(net409),
    .D(_01037_),
    .Q(\fifo_bank_register.bank[3][116] ));
 sky130_fd_sc_hd__dfxtp_1 _17595_ (.CLK(net432),
    .D(_01038_),
    .Q(\fifo_bank_register.bank[3][117] ));
 sky130_fd_sc_hd__dfxtp_1 _17596_ (.CLK(net408),
    .D(_01039_),
    .Q(\fifo_bank_register.bank[3][118] ));
 sky130_fd_sc_hd__dfxtp_1 _17597_ (.CLK(net429),
    .D(_01040_),
    .Q(\fifo_bank_register.bank[3][119] ));
 sky130_fd_sc_hd__dfxtp_1 _17598_ (.CLK(net441),
    .D(_01041_),
    .Q(\fifo_bank_register.bank[3][120] ));
 sky130_fd_sc_hd__dfxtp_1 _17599_ (.CLK(net439),
    .D(_01042_),
    .Q(\fifo_bank_register.bank[3][121] ));
 sky130_fd_sc_hd__dfxtp_1 _17600_ (.CLK(net492),
    .D(_01043_),
    .Q(\fifo_bank_register.bank[3][122] ));
 sky130_fd_sc_hd__dfxtp_1 _17601_ (.CLK(net438),
    .D(_01044_),
    .Q(\fifo_bank_register.bank[3][123] ));
 sky130_fd_sc_hd__dfxtp_1 _17602_ (.CLK(net494),
    .D(_01045_),
    .Q(\fifo_bank_register.bank[3][124] ));
 sky130_fd_sc_hd__dfxtp_1 _17603_ (.CLK(net490),
    .D(_01046_),
    .Q(\fifo_bank_register.bank[3][125] ));
 sky130_fd_sc_hd__dfxtp_1 _17604_ (.CLK(net494),
    .D(_01047_),
    .Q(\fifo_bank_register.bank[3][126] ));
 sky130_fd_sc_hd__dfxtp_1 _17605_ (.CLK(net440),
    .D(_01048_),
    .Q(\fifo_bank_register.bank[3][127] ));
 sky130_fd_sc_hd__dfxtp_1 _17606_ (.CLK(net475),
    .D(_01049_),
    .Q(\fifo_bank_register.bank[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17607_ (.CLK(net492),
    .D(_01050_),
    .Q(\fifo_bank_register.bank[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17608_ (.CLK(net475),
    .D(_01051_),
    .Q(\fifo_bank_register.bank[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17609_ (.CLK(net475),
    .D(_01052_),
    .Q(\fifo_bank_register.bank[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17610_ (.CLK(net475),
    .D(_01053_),
    .Q(\fifo_bank_register.bank[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17611_ (.CLK(net476),
    .D(_01054_),
    .Q(\fifo_bank_register.bank[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17612_ (.CLK(net479),
    .D(_01055_),
    .Q(\fifo_bank_register.bank[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17613_ (.CLK(net477),
    .D(_01056_),
    .Q(\fifo_bank_register.bank[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17614_ (.CLK(net480),
    .D(_01057_),
    .Q(\fifo_bank_register.bank[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17615_ (.CLK(net479),
    .D(_01058_),
    .Q(\fifo_bank_register.bank[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17616_ (.CLK(net496),
    .D(_01059_),
    .Q(\fifo_bank_register.bank[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17617_ (.CLK(net503),
    .D(_01060_),
    .Q(\fifo_bank_register.bank[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17618_ (.CLK(net500),
    .D(_01061_),
    .Q(\fifo_bank_register.bank[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17619_ (.CLK(net505),
    .D(_01062_),
    .Q(\fifo_bank_register.bank[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17620_ (.CLK(net506),
    .D(_01063_),
    .Q(\fifo_bank_register.bank[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17621_ (.CLK(net534),
    .D(_01064_),
    .Q(\fifo_bank_register.bank[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17622_ (.CLK(net496),
    .D(_01065_),
    .Q(\fifo_bank_register.bank[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17623_ (.CLK(net497),
    .D(_01066_),
    .Q(\fifo_bank_register.bank[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17624_ (.CLK(net503),
    .D(_01067_),
    .Q(\fifo_bank_register.bank[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17625_ (.CLK(net501),
    .D(_01068_),
    .Q(\fifo_bank_register.bank[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17626_ (.CLK(net512),
    .D(_01069_),
    .Q(\fifo_bank_register.bank[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17627_ (.CLK(net483),
    .D(_01070_),
    .Q(\fifo_bank_register.bank[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17628_ (.CLK(net501),
    .D(_01071_),
    .Q(\fifo_bank_register.bank[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17629_ (.CLK(net487),
    .D(_01072_),
    .Q(\fifo_bank_register.bank[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17630_ (.CLK(net485),
    .D(_01073_),
    .Q(\fifo_bank_register.bank[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17631_ (.CLK(net508),
    .D(_01074_),
    .Q(\fifo_bank_register.bank[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17632_ (.CLK(net508),
    .D(_01075_),
    .Q(\fifo_bank_register.bank[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17633_ (.CLK(net486),
    .D(_01076_),
    .Q(\fifo_bank_register.bank[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17634_ (.CLK(net486),
    .D(_01077_),
    .Q(\fifo_bank_register.bank[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17635_ (.CLK(net499),
    .D(_01078_),
    .Q(\fifo_bank_register.bank[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17636_ (.CLK(net418),
    .D(_01079_),
    .Q(\fifo_bank_register.bank[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17637_ (.CLK(net423),
    .D(_01080_),
    .Q(\fifo_bank_register.bank[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17638_ (.CLK(net419),
    .D(_01081_),
    .Q(\fifo_bank_register.bank[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 _17639_ (.CLK(net424),
    .D(_01082_),
    .Q(\fifo_bank_register.bank[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 _17640_ (.CLK(net418),
    .D(_01083_),
    .Q(\fifo_bank_register.bank[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 _17641_ (.CLK(net416),
    .D(_01084_),
    .Q(\fifo_bank_register.bank[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 _17642_ (.CLK(net422),
    .D(_01085_),
    .Q(\fifo_bank_register.bank[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 _17643_ (.CLK(net414),
    .D(_01086_),
    .Q(\fifo_bank_register.bank[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 _17644_ (.CLK(net416),
    .D(_01087_),
    .Q(\fifo_bank_register.bank[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 _17645_ (.CLK(net414),
    .D(_01088_),
    .Q(\fifo_bank_register.bank[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 _17646_ (.CLK(net397),
    .D(_01089_),
    .Q(\fifo_bank_register.bank[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 _17647_ (.CLK(net398),
    .D(_01090_),
    .Q(\fifo_bank_register.bank[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 _17648_ (.CLK(net389),
    .D(_01091_),
    .Q(\fifo_bank_register.bank[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 _17649_ (.CLK(net392),
    .D(_01092_),
    .Q(\fifo_bank_register.bank[2][43] ));
 sky130_fd_sc_hd__dfxtp_1 _17650_ (.CLK(net391),
    .D(_01093_),
    .Q(\fifo_bank_register.bank[2][44] ));
 sky130_fd_sc_hd__dfxtp_1 _17651_ (.CLK(net405),
    .D(_01094_),
    .Q(\fifo_bank_register.bank[2][45] ));
 sky130_fd_sc_hd__dfxtp_1 _17652_ (.CLK(net391),
    .D(_01095_),
    .Q(\fifo_bank_register.bank[2][46] ));
 sky130_fd_sc_hd__dfxtp_1 _17653_ (.CLK(net396),
    .D(_01096_),
    .Q(\fifo_bank_register.bank[2][47] ));
 sky130_fd_sc_hd__dfxtp_1 _17654_ (.CLK(net397),
    .D(_01097_),
    .Q(\fifo_bank_register.bank[2][48] ));
 sky130_fd_sc_hd__dfxtp_1 _17655_ (.CLK(net407),
    .D(_01098_),
    .Q(\fifo_bank_register.bank[2][49] ));
 sky130_fd_sc_hd__dfxtp_1 _17656_ (.CLK(net556),
    .D(_01099_),
    .Q(\fifo_bank_register.bank[2][50] ));
 sky130_fd_sc_hd__dfxtp_1 _17657_ (.CLK(net573),
    .D(_01100_),
    .Q(\fifo_bank_register.bank[2][51] ));
 sky130_fd_sc_hd__dfxtp_1 _17658_ (.CLK(net563),
    .D(_01101_),
    .Q(\fifo_bank_register.bank[2][52] ));
 sky130_fd_sc_hd__dfxtp_1 _17659_ (.CLK(net562),
    .D(_01102_),
    .Q(\fifo_bank_register.bank[2][53] ));
 sky130_fd_sc_hd__dfxtp_1 _17660_ (.CLK(net556),
    .D(_01103_),
    .Q(\fifo_bank_register.bank[2][54] ));
 sky130_fd_sc_hd__dfxtp_1 _17661_ (.CLK(net571),
    .D(_01104_),
    .Q(\fifo_bank_register.bank[2][55] ));
 sky130_fd_sc_hd__dfxtp_1 _17662_ (.CLK(net571),
    .D(_01105_),
    .Q(\fifo_bank_register.bank[2][56] ));
 sky130_fd_sc_hd__dfxtp_1 _17663_ (.CLK(net550),
    .D(_01106_),
    .Q(\fifo_bank_register.bank[2][57] ));
 sky130_fd_sc_hd__dfxtp_1 _17664_ (.CLK(net557),
    .D(_01107_),
    .Q(\fifo_bank_register.bank[2][58] ));
 sky130_fd_sc_hd__dfxtp_1 _17665_ (.CLK(net572),
    .D(_01108_),
    .Q(\fifo_bank_register.bank[2][59] ));
 sky130_fd_sc_hd__dfxtp_1 _17666_ (.CLK(net513),
    .D(_01109_),
    .Q(\fifo_bank_register.bank[2][60] ));
 sky130_fd_sc_hd__dfxtp_1 _17667_ (.CLK(net526),
    .D(_01110_),
    .Q(\fifo_bank_register.bank[2][61] ));
 sky130_fd_sc_hd__dfxtp_1 _17668_ (.CLK(net523),
    .D(_01111_),
    .Q(\fifo_bank_register.bank[2][62] ));
 sky130_fd_sc_hd__dfxtp_1 _17669_ (.CLK(net524),
    .D(_01112_),
    .Q(\fifo_bank_register.bank[2][63] ));
 sky130_fd_sc_hd__dfxtp_1 _17670_ (.CLK(net512),
    .D(_01113_),
    .Q(\fifo_bank_register.bank[2][64] ));
 sky130_fd_sc_hd__dfxtp_1 _17671_ (.CLK(net526),
    .D(_01114_),
    .Q(\fifo_bank_register.bank[2][65] ));
 sky130_fd_sc_hd__dfxtp_1 _17672_ (.CLK(net521),
    .D(_01115_),
    .Q(\fifo_bank_register.bank[2][66] ));
 sky130_fd_sc_hd__dfxtp_1 _17673_ (.CLK(net515),
    .D(_01116_),
    .Q(\fifo_bank_register.bank[2][67] ));
 sky130_fd_sc_hd__dfxtp_1 _17674_ (.CLK(net521),
    .D(_01117_),
    .Q(\fifo_bank_register.bank[2][68] ));
 sky130_fd_sc_hd__dfxtp_1 _17675_ (.CLK(net516),
    .D(_01118_),
    .Q(\fifo_bank_register.bank[2][69] ));
 sky130_fd_sc_hd__dfxtp_1 _17676_ (.CLK(net519),
    .D(_01119_),
    .Q(\fifo_bank_register.bank[2][70] ));
 sky130_fd_sc_hd__dfxtp_1 _17677_ (.CLK(net517),
    .D(_01120_),
    .Q(\fifo_bank_register.bank[2][71] ));
 sky130_fd_sc_hd__dfxtp_1 _17678_ (.CLK(net544),
    .D(_01121_),
    .Q(\fifo_bank_register.bank[2][72] ));
 sky130_fd_sc_hd__dfxtp_1 _17679_ (.CLK(net543),
    .D(_01122_),
    .Q(\fifo_bank_register.bank[2][73] ));
 sky130_fd_sc_hd__dfxtp_1 _17680_ (.CLK(net549),
    .D(_01123_),
    .Q(\fifo_bank_register.bank[2][74] ));
 sky130_fd_sc_hd__dfxtp_1 _17681_ (.CLK(net544),
    .D(_01124_),
    .Q(\fifo_bank_register.bank[2][75] ));
 sky130_fd_sc_hd__dfxtp_1 _17682_ (.CLK(net543),
    .D(_01125_),
    .Q(\fifo_bank_register.bank[2][76] ));
 sky130_fd_sc_hd__dfxtp_1 _17683_ (.CLK(net546),
    .D(_01126_),
    .Q(\fifo_bank_register.bank[2][77] ));
 sky130_fd_sc_hd__dfxtp_1 _17684_ (.CLK(net517),
    .D(_01127_),
    .Q(\fifo_bank_register.bank[2][78] ));
 sky130_fd_sc_hd__dfxtp_1 _17685_ (.CLK(net547),
    .D(_01128_),
    .Q(\fifo_bank_register.bank[2][79] ));
 sky130_fd_sc_hd__dfxtp_1 _17686_ (.CLK(net541),
    .D(_01129_),
    .Q(\fifo_bank_register.bank[2][80] ));
 sky130_fd_sc_hd__dfxtp_1 _17687_ (.CLK(net540),
    .D(_01130_),
    .Q(\fifo_bank_register.bank[2][81] ));
 sky130_fd_sc_hd__dfxtp_1 _17688_ (.CLK(net539),
    .D(_01131_),
    .Q(\fifo_bank_register.bank[2][82] ));
 sky130_fd_sc_hd__dfxtp_1 _17689_ (.CLK(net539),
    .D(_01132_),
    .Q(\fifo_bank_register.bank[2][83] ));
 sky130_fd_sc_hd__dfxtp_1 _17690_ (.CLK(net536),
    .D(_01133_),
    .Q(\fifo_bank_register.bank[2][84] ));
 sky130_fd_sc_hd__dfxtp_1 _17691_ (.CLK(net540),
    .D(_01134_),
    .Q(\fifo_bank_register.bank[2][85] ));
 sky130_fd_sc_hd__dfxtp_1 _17692_ (.CLK(net538),
    .D(_01135_),
    .Q(\fifo_bank_register.bank[2][86] ));
 sky130_fd_sc_hd__dfxtp_1 _17693_ (.CLK(net538),
    .D(_01136_),
    .Q(\fifo_bank_register.bank[2][87] ));
 sky130_fd_sc_hd__dfxtp_1 _17694_ (.CLK(net541),
    .D(_01137_),
    .Q(\fifo_bank_register.bank[2][88] ));
 sky130_fd_sc_hd__dfxtp_1 _17695_ (.CLK(net536),
    .D(_01138_),
    .Q(\fifo_bank_register.bank[2][89] ));
 sky130_fd_sc_hd__dfxtp_1 _17696_ (.CLK(net409),
    .D(_01139_),
    .Q(\fifo_bank_register.bank[2][90] ));
 sky130_fd_sc_hd__dfxtp_1 _17697_ (.CLK(net401),
    .D(_01140_),
    .Q(\fifo_bank_register.bank[2][91] ));
 sky130_fd_sc_hd__dfxtp_1 _17698_ (.CLK(net410),
    .D(_01141_),
    .Q(\fifo_bank_register.bank[2][92] ));
 sky130_fd_sc_hd__dfxtp_1 _17699_ (.CLK(net400),
    .D(_01142_),
    .Q(\fifo_bank_register.bank[2][93] ));
 sky130_fd_sc_hd__dfxtp_1 _17700_ (.CLK(net447),
    .D(_01143_),
    .Q(\fifo_bank_register.bank[2][94] ));
 sky130_fd_sc_hd__dfxtp_1 _17701_ (.CLK(net400),
    .D(_01144_),
    .Q(\fifo_bank_register.bank[2][95] ));
 sky130_fd_sc_hd__dfxtp_1 _17702_ (.CLK(net445),
    .D(_01145_),
    .Q(\fifo_bank_register.bank[2][96] ));
 sky130_fd_sc_hd__dfxtp_1 _17703_ (.CLK(net448),
    .D(_01146_),
    .Q(\fifo_bank_register.bank[2][97] ));
 sky130_fd_sc_hd__dfxtp_1 _17704_ (.CLK(net446),
    .D(_01147_),
    .Q(\fifo_bank_register.bank[2][98] ));
 sky130_fd_sc_hd__dfxtp_1 _17705_ (.CLK(net446),
    .D(_01148_),
    .Q(\fifo_bank_register.bank[2][99] ));
 sky130_fd_sc_hd__dfxtp_1 _17706_ (.CLK(net452),
    .D(_01149_),
    .Q(\fifo_bank_register.bank[2][100] ));
 sky130_fd_sc_hd__dfxtp_1 _17707_ (.CLK(net450),
    .D(_01150_),
    .Q(\fifo_bank_register.bank[2][101] ));
 sky130_fd_sc_hd__dfxtp_1 _17708_ (.CLK(net464),
    .D(_01151_),
    .Q(\fifo_bank_register.bank[2][102] ));
 sky130_fd_sc_hd__dfxtp_1 _17709_ (.CLK(net453),
    .D(_01152_),
    .Q(\fifo_bank_register.bank[2][103] ));
 sky130_fd_sc_hd__dfxtp_1 _17710_ (.CLK(net462),
    .D(_01153_),
    .Q(\fifo_bank_register.bank[2][104] ));
 sky130_fd_sc_hd__dfxtp_1 _17711_ (.CLK(net467),
    .D(_01154_),
    .Q(\fifo_bank_register.bank[2][105] ));
 sky130_fd_sc_hd__dfxtp_1 _17712_ (.CLK(net464),
    .D(_01155_),
    .Q(\fifo_bank_register.bank[2][106] ));
 sky130_fd_sc_hd__dfxtp_1 _17713_ (.CLK(net462),
    .D(_01156_),
    .Q(\fifo_bank_register.bank[2][107] ));
 sky130_fd_sc_hd__dfxtp_1 _17714_ (.CLK(net450),
    .D(_01157_),
    .Q(\fifo_bank_register.bank[2][108] ));
 sky130_fd_sc_hd__dfxtp_1 _17715_ (.CLK(net458),
    .D(_01158_),
    .Q(\fifo_bank_register.bank[2][109] ));
 sky130_fd_sc_hd__dfxtp_1 _17716_ (.CLK(net434),
    .D(_01159_),
    .Q(\fifo_bank_register.bank[2][110] ));
 sky130_fd_sc_hd__dfxtp_1 _17717_ (.CLK(net412),
    .D(_01160_),
    .Q(\fifo_bank_register.bank[2][111] ));
 sky130_fd_sc_hd__dfxtp_1 _17718_ (.CLK(net432),
    .D(_01161_),
    .Q(\fifo_bank_register.bank[2][112] ));
 sky130_fd_sc_hd__dfxtp_1 _17719_ (.CLK(net432),
    .D(_01162_),
    .Q(\fifo_bank_register.bank[2][113] ));
 sky130_fd_sc_hd__dfxtp_1 _17720_ (.CLK(net408),
    .D(_01163_),
    .Q(\fifo_bank_register.bank[2][114] ));
 sky130_fd_sc_hd__dfxtp_1 _17721_ (.CLK(net430),
    .D(_01164_),
    .Q(\fifo_bank_register.bank[2][115] ));
 sky130_fd_sc_hd__dfxtp_1 _17722_ (.CLK(net412),
    .D(_01165_),
    .Q(\fifo_bank_register.bank[2][116] ));
 sky130_fd_sc_hd__dfxtp_1 _17723_ (.CLK(net434),
    .D(_01166_),
    .Q(\fifo_bank_register.bank[2][117] ));
 sky130_fd_sc_hd__dfxtp_1 _17724_ (.CLK(net407),
    .D(_01167_),
    .Q(\fifo_bank_register.bank[2][118] ));
 sky130_fd_sc_hd__dfxtp_1 _17725_ (.CLK(net430),
    .D(_01168_),
    .Q(\fifo_bank_register.bank[2][119] ));
 sky130_fd_sc_hd__dfxtp_1 _17726_ (.CLK(net441),
    .D(_01169_),
    .Q(\fifo_bank_register.bank[2][120] ));
 sky130_fd_sc_hd__dfxtp_1 _17727_ (.CLK(net491),
    .D(_01170_),
    .Q(\fifo_bank_register.bank[2][121] ));
 sky130_fd_sc_hd__dfxtp_1 _17728_ (.CLK(net493),
    .D(_01171_),
    .Q(\fifo_bank_register.bank[2][122] ));
 sky130_fd_sc_hd__dfxtp_1 _17729_ (.CLK(net439),
    .D(_01172_),
    .Q(\fifo_bank_register.bank[2][123] ));
 sky130_fd_sc_hd__dfxtp_1 _17730_ (.CLK(net494),
    .D(_01173_),
    .Q(\fifo_bank_register.bank[2][124] ));
 sky130_fd_sc_hd__dfxtp_1 _17731_ (.CLK(net494),
    .D(_01174_),
    .Q(\fifo_bank_register.bank[2][125] ));
 sky130_fd_sc_hd__dfxtp_1 _17732_ (.CLK(net494),
    .D(_01175_),
    .Q(\fifo_bank_register.bank[2][126] ));
 sky130_fd_sc_hd__dfxtp_1 _17733_ (.CLK(net441),
    .D(_01176_),
    .Q(\fifo_bank_register.bank[2][127] ));
 sky130_fd_sc_hd__dfxtp_1 _17734_ (.CLK(net473),
    .D(_01177_),
    .Q(\fifo_bank_register.bank[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17735_ (.CLK(net439),
    .D(_01178_),
    .Q(\fifo_bank_register.bank[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17736_ (.CLK(net420),
    .D(_01179_),
    .Q(\fifo_bank_register.bank[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17737_ (.CLK(net473),
    .D(_01180_),
    .Q(\fifo_bank_register.bank[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17738_ (.CLK(net474),
    .D(_01181_),
    .Q(\fifo_bank_register.bank[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17739_ (.CLK(net473),
    .D(_01182_),
    .Q(\fifo_bank_register.bank[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17740_ (.CLK(net477),
    .D(_01183_),
    .Q(\fifo_bank_register.bank[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17741_ (.CLK(net477),
    .D(_01184_),
    .Q(\fifo_bank_register.bank[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17742_ (.CLK(net477),
    .D(_01185_),
    .Q(\fifo_bank_register.bank[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17743_ (.CLK(net478),
    .D(_01186_),
    .Q(\fifo_bank_register.bank[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17744_ (.CLK(net503),
    .D(_01187_),
    .Q(\fifo_bank_register.bank[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17745_ (.CLK(net533),
    .D(_01188_),
    .Q(\fifo_bank_register.bank[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17746_ (.CLK(net504),
    .D(_01189_),
    .Q(\fifo_bank_register.bank[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17747_ (.CLK(net516),
    .D(_01190_),
    .Q(\fifo_bank_register.bank[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17748_ (.CLK(net534),
    .D(_01191_),
    .Q(\fifo_bank_register.bank[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17749_ (.CLK(net517),
    .D(_01192_),
    .Q(\fifo_bank_register.bank[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17750_ (.CLK(net497),
    .D(_01193_),
    .Q(\fifo_bank_register.bank[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17751_ (.CLK(net532),
    .D(_01194_),
    .Q(\fifo_bank_register.bank[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17752_ (.CLK(net533),
    .D(_01195_),
    .Q(\fifo_bank_register.bank[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17753_ (.CLK(net516),
    .D(_01196_),
    .Q(\fifo_bank_register.bank[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17754_ (.CLK(net501),
    .D(_01197_),
    .Q(\fifo_bank_register.bank[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17755_ (.CLK(net482),
    .D(_01198_),
    .Q(\fifo_bank_register.bank[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17756_ (.CLK(net501),
    .D(_01199_),
    .Q(\fifo_bank_register.bank[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17757_ (.CLK(net483),
    .D(_01200_),
    .Q(\fifo_bank_register.bank[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17758_ (.CLK(net482),
    .D(_01201_),
    .Q(\fifo_bank_register.bank[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17759_ (.CLK(net488),
    .D(_01202_),
    .Q(\fifo_bank_register.bank[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17760_ (.CLK(net483),
    .D(_01203_),
    .Q(\fifo_bank_register.bank[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17761_ (.CLK(net486),
    .D(_01204_),
    .Q(\fifo_bank_register.bank[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17762_ (.CLK(net486),
    .D(_01205_),
    .Q(\fifo_bank_register.bank[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17763_ (.CLK(net499),
    .D(_01206_),
    .Q(\fifo_bank_register.bank[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17764_ (.CLK(net437),
    .D(_01207_),
    .Q(\fifo_bank_register.bank[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17765_ (.CLK(net437),
    .D(_01208_),
    .Q(\fifo_bank_register.bank[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17766_ (.CLK(net417),
    .D(_01209_),
    .Q(\fifo_bank_register.bank[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 _17767_ (.CLK(net423),
    .D(_01210_),
    .Q(\fifo_bank_register.bank[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 _17768_ (.CLK(net430),
    .D(_01211_),
    .Q(\fifo_bank_register.bank[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 _17769_ (.CLK(net428),
    .D(_01212_),
    .Q(\fifo_bank_register.bank[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 _17770_ (.CLK(net422),
    .D(_01213_),
    .Q(\fifo_bank_register.bank[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 _17771_ (.CLK(net417),
    .D(_01214_),
    .Q(\fifo_bank_register.bank[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 _17772_ (.CLK(net416),
    .D(_01215_),
    .Q(\fifo_bank_register.bank[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 _17773_ (.CLK(net415),
    .D(_01216_),
    .Q(\fifo_bank_register.bank[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 _17774_ (.CLK(net395),
    .D(_01217_),
    .Q(\fifo_bank_register.bank[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 _17775_ (.CLK(net398),
    .D(_01218_),
    .Q(\fifo_bank_register.bank[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 _17776_ (.CLK(net394),
    .D(_01219_),
    .Q(\fifo_bank_register.bank[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 _17777_ (.CLK(net393),
    .D(_01220_),
    .Q(\fifo_bank_register.bank[1][43] ));
 sky130_fd_sc_hd__dfxtp_1 _17778_ (.CLK(net389),
    .D(_01221_),
    .Q(\fifo_bank_register.bank[1][44] ));
 sky130_fd_sc_hd__dfxtp_1 _17779_ (.CLK(net405),
    .D(_01222_),
    .Q(\fifo_bank_register.bank[1][45] ));
 sky130_fd_sc_hd__dfxtp_1 _17780_ (.CLK(net394),
    .D(_01223_),
    .Q(\fifo_bank_register.bank[1][46] ));
 sky130_fd_sc_hd__dfxtp_1 _17781_ (.CLK(net393),
    .D(_01224_),
    .Q(\fifo_bank_register.bank[1][47] ));
 sky130_fd_sc_hd__dfxtp_1 _17782_ (.CLK(net393),
    .D(_01225_),
    .Q(\fifo_bank_register.bank[1][48] ));
 sky130_fd_sc_hd__dfxtp_1 _17783_ (.CLK(net407),
    .D(_01226_),
    .Q(\fifo_bank_register.bank[1][49] ));
 sky130_fd_sc_hd__dfxtp_1 _17784_ (.CLK(net557),
    .D(_01227_),
    .Q(\fifo_bank_register.bank[1][50] ));
 sky130_fd_sc_hd__dfxtp_1 _17785_ (.CLK(net573),
    .D(_01228_),
    .Q(\fifo_bank_register.bank[1][51] ));
 sky130_fd_sc_hd__dfxtp_1 _17786_ (.CLK(net563),
    .D(_01229_),
    .Q(\fifo_bank_register.bank[1][52] ));
 sky130_fd_sc_hd__dfxtp_1 _17787_ (.CLK(net562),
    .D(_01230_),
    .Q(\fifo_bank_register.bank[1][53] ));
 sky130_fd_sc_hd__dfxtp_1 _17788_ (.CLK(net570),
    .D(_01231_),
    .Q(\fifo_bank_register.bank[1][54] ));
 sky130_fd_sc_hd__dfxtp_1 _17789_ (.CLK(net571),
    .D(_01232_),
    .Q(\fifo_bank_register.bank[1][55] ));
 sky130_fd_sc_hd__dfxtp_1 _17790_ (.CLK(net571),
    .D(_01233_),
    .Q(\fifo_bank_register.bank[1][56] ));
 sky130_fd_sc_hd__dfxtp_1 _17791_ (.CLK(net550),
    .D(_01234_),
    .Q(\fifo_bank_register.bank[1][57] ));
 sky130_fd_sc_hd__dfxtp_1 _17792_ (.CLK(net558),
    .D(_01235_),
    .Q(\fifo_bank_register.bank[1][58] ));
 sky130_fd_sc_hd__dfxtp_1 _17793_ (.CLK(net572),
    .D(_01236_),
    .Q(\fifo_bank_register.bank[1][59] ));
 sky130_fd_sc_hd__dfxtp_1 _17794_ (.CLK(net514),
    .D(_01237_),
    .Q(\fifo_bank_register.bank[1][60] ));
 sky130_fd_sc_hd__dfxtp_1 _17795_ (.CLK(net527),
    .D(_01238_),
    .Q(\fifo_bank_register.bank[1][61] ));
 sky130_fd_sc_hd__dfxtp_1 _17796_ (.CLK(net511),
    .D(_01239_),
    .Q(\fifo_bank_register.bank[1][62] ));
 sky130_fd_sc_hd__dfxtp_1 _17797_ (.CLK(net524),
    .D(_01240_),
    .Q(\fifo_bank_register.bank[1][63] ));
 sky130_fd_sc_hd__dfxtp_1 _17798_ (.CLK(net509),
    .D(_01241_),
    .Q(\fifo_bank_register.bank[1][64] ));
 sky130_fd_sc_hd__dfxtp_1 _17799_ (.CLK(net518),
    .D(_01242_),
    .Q(\fifo_bank_register.bank[1][65] ));
 sky130_fd_sc_hd__dfxtp_1 _17800_ (.CLK(net527),
    .D(_01243_),
    .Q(\fifo_bank_register.bank[1][66] ));
 sky130_fd_sc_hd__dfxtp_1 _17801_ (.CLK(net511),
    .D(_01244_),
    .Q(\fifo_bank_register.bank[1][67] ));
 sky130_fd_sc_hd__dfxtp_1 _17802_ (.CLK(net511),
    .D(_01245_),
    .Q(\fifo_bank_register.bank[1][68] ));
 sky130_fd_sc_hd__dfxtp_1 _17803_ (.CLK(net518),
    .D(_01246_),
    .Q(\fifo_bank_register.bank[1][69] ));
 sky130_fd_sc_hd__dfxtp_1 _17804_ (.CLK(net519),
    .D(_01247_),
    .Q(\fifo_bank_register.bank[1][70] ));
 sky130_fd_sc_hd__dfxtp_1 _17805_ (.CLK(net525),
    .D(_01248_),
    .Q(\fifo_bank_register.bank[1][71] ));
 sky130_fd_sc_hd__dfxtp_1 _17806_ (.CLK(net552),
    .D(_01249_),
    .Q(\fifo_bank_register.bank[1][72] ));
 sky130_fd_sc_hd__dfxtp_1 _17807_ (.CLK(net552),
    .D(_01250_),
    .Q(\fifo_bank_register.bank[1][73] ));
 sky130_fd_sc_hd__dfxtp_1 _17808_ (.CLK(net546),
    .D(_01251_),
    .Q(\fifo_bank_register.bank[1][74] ));
 sky130_fd_sc_hd__dfxtp_1 _17809_ (.CLK(net552),
    .D(_01252_),
    .Q(\fifo_bank_register.bank[1][75] ));
 sky130_fd_sc_hd__dfxtp_1 _17810_ (.CLK(net545),
    .D(_01253_),
    .Q(\fifo_bank_register.bank[1][76] ));
 sky130_fd_sc_hd__dfxtp_1 _17811_ (.CLK(net553),
    .D(_01254_),
    .Q(\fifo_bank_register.bank[1][77] ));
 sky130_fd_sc_hd__dfxtp_1 _17812_ (.CLK(net525),
    .D(_01255_),
    .Q(\fifo_bank_register.bank[1][78] ));
 sky130_fd_sc_hd__dfxtp_1 _17813_ (.CLK(net546),
    .D(_01256_),
    .Q(\fifo_bank_register.bank[1][79] ));
 sky130_fd_sc_hd__dfxtp_1 _17814_ (.CLK(net566),
    .D(_01257_),
    .Q(\fifo_bank_register.bank[1][80] ));
 sky130_fd_sc_hd__dfxtp_1 _17815_ (.CLK(net561),
    .D(_01258_),
    .Q(\fifo_bank_register.bank[1][81] ));
 sky130_fd_sc_hd__dfxtp_1 _17816_ (.CLK(net560),
    .D(_01259_),
    .Q(\fifo_bank_register.bank[1][82] ));
 sky130_fd_sc_hd__dfxtp_1 _17817_ (.CLK(net561),
    .D(_01260_),
    .Q(\fifo_bank_register.bank[1][83] ));
 sky130_fd_sc_hd__dfxtp_1 _17818_ (.CLK(net547),
    .D(_01261_),
    .Q(\fifo_bank_register.bank[1][84] ));
 sky130_fd_sc_hd__dfxtp_1 _17819_ (.CLK(net566),
    .D(_01262_),
    .Q(\fifo_bank_register.bank[1][85] ));
 sky130_fd_sc_hd__dfxtp_1 _17820_ (.CLK(net548),
    .D(_01263_),
    .Q(\fifo_bank_register.bank[1][86] ));
 sky130_fd_sc_hd__dfxtp_1 _17821_ (.CLK(net561),
    .D(_01264_),
    .Q(\fifo_bank_register.bank[1][87] ));
 sky130_fd_sc_hd__dfxtp_1 _17822_ (.CLK(net566),
    .D(_01265_),
    .Q(\fifo_bank_register.bank[1][88] ));
 sky130_fd_sc_hd__dfxtp_1 _17823_ (.CLK(net547),
    .D(_01266_),
    .Q(\fifo_bank_register.bank[1][89] ));
 sky130_fd_sc_hd__dfxtp_1 _17824_ (.CLK(net409),
    .D(_01267_),
    .Q(\fifo_bank_register.bank[1][90] ));
 sky130_fd_sc_hd__dfxtp_1 _17825_ (.CLK(net401),
    .D(_01268_),
    .Q(\fifo_bank_register.bank[1][91] ));
 sky130_fd_sc_hd__dfxtp_1 _17826_ (.CLK(net410),
    .D(_01269_),
    .Q(\fifo_bank_register.bank[1][92] ));
 sky130_fd_sc_hd__dfxtp_1 _17827_ (.CLK(net404),
    .D(_01270_),
    .Q(\fifo_bank_register.bank[1][93] ));
 sky130_fd_sc_hd__dfxtp_1 _17828_ (.CLK(net454),
    .D(_01271_),
    .Q(\fifo_bank_register.bank[1][94] ));
 sky130_fd_sc_hd__dfxtp_1 _17829_ (.CLK(net402),
    .D(_01272_),
    .Q(\fifo_bank_register.bank[1][95] ));
 sky130_fd_sc_hd__dfxtp_1 _17830_ (.CLK(net445),
    .D(_01273_),
    .Q(\fifo_bank_register.bank[1][96] ));
 sky130_fd_sc_hd__dfxtp_1 _17831_ (.CLK(net454),
    .D(_01274_),
    .Q(\fifo_bank_register.bank[1][97] ));
 sky130_fd_sc_hd__dfxtp_1 _17832_ (.CLK(net448),
    .D(_01275_),
    .Q(\fifo_bank_register.bank[1][98] ));
 sky130_fd_sc_hd__dfxtp_1 _17833_ (.CLK(net448),
    .D(_01276_),
    .Q(\fifo_bank_register.bank[1][99] ));
 sky130_fd_sc_hd__dfxtp_1 _17834_ (.CLK(net452),
    .D(_01277_),
    .Q(\fifo_bank_register.bank[1][100] ));
 sky130_fd_sc_hd__dfxtp_1 _17835_ (.CLK(net450),
    .D(_01278_),
    .Q(\fifo_bank_register.bank[1][101] ));
 sky130_fd_sc_hd__dfxtp_1 _17836_ (.CLK(net465),
    .D(_01279_),
    .Q(\fifo_bank_register.bank[1][102] ));
 sky130_fd_sc_hd__dfxtp_1 _17837_ (.CLK(net458),
    .D(_01280_),
    .Q(\fifo_bank_register.bank[1][103] ));
 sky130_fd_sc_hd__dfxtp_1 _17838_ (.CLK(net463),
    .D(_01281_),
    .Q(\fifo_bank_register.bank[1][104] ));
 sky130_fd_sc_hd__dfxtp_1 _17839_ (.CLK(net468),
    .D(_01282_),
    .Q(\fifo_bank_register.bank[1][105] ));
 sky130_fd_sc_hd__dfxtp_1 _17840_ (.CLK(net465),
    .D(_01283_),
    .Q(\fifo_bank_register.bank[1][106] ));
 sky130_fd_sc_hd__dfxtp_1 _17841_ (.CLK(net451),
    .D(_01284_),
    .Q(\fifo_bank_register.bank[1][107] ));
 sky130_fd_sc_hd__dfxtp_1 _17842_ (.CLK(net453),
    .D(_01285_),
    .Q(\fifo_bank_register.bank[1][108] ));
 sky130_fd_sc_hd__dfxtp_1 _17843_ (.CLK(net458),
    .D(_01286_),
    .Q(\fifo_bank_register.bank[1][109] ));
 sky130_fd_sc_hd__dfxtp_1 _17844_ (.CLK(net432),
    .D(_01287_),
    .Q(\fifo_bank_register.bank[1][110] ));
 sky130_fd_sc_hd__dfxtp_1 _17845_ (.CLK(net411),
    .D(_01288_),
    .Q(\fifo_bank_register.bank[1][111] ));
 sky130_fd_sc_hd__dfxtp_1 _17846_ (.CLK(net433),
    .D(_01289_),
    .Q(\fifo_bank_register.bank[1][112] ));
 sky130_fd_sc_hd__dfxtp_1 _17847_ (.CLK(net469),
    .D(_01290_),
    .Q(\fifo_bank_register.bank[1][113] ));
 sky130_fd_sc_hd__dfxtp_1 _17848_ (.CLK(net457),
    .D(_01291_),
    .Q(\fifo_bank_register.bank[1][114] ));
 sky130_fd_sc_hd__dfxtp_1 _17849_ (.CLK(net469),
    .D(_01292_),
    .Q(\fifo_bank_register.bank[1][115] ));
 sky130_fd_sc_hd__dfxtp_1 _17850_ (.CLK(net456),
    .D(_01293_),
    .Q(\fifo_bank_register.bank[1][116] ));
 sky130_fd_sc_hd__dfxtp_1 _17851_ (.CLK(net433),
    .D(_01294_),
    .Q(\fifo_bank_register.bank[1][117] ));
 sky130_fd_sc_hd__dfxtp_1 _17852_ (.CLK(net470),
    .D(_01295_),
    .Q(\fifo_bank_register.bank[1][118] ));
 sky130_fd_sc_hd__dfxtp_1 _17853_ (.CLK(net469),
    .D(_01296_),
    .Q(\fifo_bank_register.bank[1][119] ));
 sky130_fd_sc_hd__dfxtp_1 _17854_ (.CLK(net471),
    .D(_01297_),
    .Q(\fifo_bank_register.bank[1][120] ));
 sky130_fd_sc_hd__dfxtp_1 _17855_ (.CLK(net491),
    .D(_01298_),
    .Q(\fifo_bank_register.bank[1][121] ));
 sky130_fd_sc_hd__dfxtp_1 _17856_ (.CLK(net493),
    .D(_01299_),
    .Q(\fifo_bank_register.bank[1][122] ));
 sky130_fd_sc_hd__dfxtp_1 _17857_ (.CLK(net439),
    .D(_01300_),
    .Q(\fifo_bank_register.bank[1][123] ));
 sky130_fd_sc_hd__dfxtp_1 _17858_ (.CLK(net531),
    .D(_01301_),
    .Q(\fifo_bank_register.bank[1][124] ));
 sky130_fd_sc_hd__dfxtp_1 _17859_ (.CLK(net496),
    .D(_01302_),
    .Q(\fifo_bank_register.bank[1][125] ));
 sky130_fd_sc_hd__dfxtp_1 _17860_ (.CLK(net531),
    .D(_01303_),
    .Q(\fifo_bank_register.bank[1][126] ));
 sky130_fd_sc_hd__dfxtp_1 _17861_ (.CLK(net471),
    .D(_01304_),
    .Q(\fifo_bank_register.bank[1][127] ));
 sky130_fd_sc_hd__dfxtp_1 _17862_ (.CLK(net421),
    .D(_01305_),
    .Q(\fifo_bank_register.bank[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _17863_ (.CLK(net439),
    .D(_01306_),
    .Q(\fifo_bank_register.bank[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _17864_ (.CLK(net420),
    .D(_01307_),
    .Q(\fifo_bank_register.bank[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _17865_ (.CLK(net420),
    .D(_01308_),
    .Q(\fifo_bank_register.bank[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _17866_ (.CLK(net420),
    .D(_01309_),
    .Q(\fifo_bank_register.bank[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _17867_ (.CLK(net421),
    .D(_01310_),
    .Q(\fifo_bank_register.bank[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _17868_ (.CLK(net425),
    .D(_01311_),
    .Q(\fifo_bank_register.bank[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _17869_ (.CLK(net425),
    .D(_01312_),
    .Q(\fifo_bank_register.bank[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _17870_ (.CLK(net426),
    .D(_01313_),
    .Q(\fifo_bank_register.bank[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _17871_ (.CLK(net426),
    .D(_01314_),
    .Q(\fifo_bank_register.bank[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _17872_ (.CLK(net500),
    .D(_01315_),
    .Q(\fifo_bank_register.bank[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _17873_ (.CLK(net533),
    .D(_01316_),
    .Q(\fifo_bank_register.bank[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _17874_ (.CLK(net500),
    .D(_01317_),
    .Q(\fifo_bank_register.bank[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _17875_ (.CLK(net506),
    .D(_01318_),
    .Q(\fifo_bank_register.bank[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _17876_ (.CLK(net535),
    .D(_01319_),
    .Q(\fifo_bank_register.bank[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _17877_ (.CLK(net535),
    .D(_01320_),
    .Q(\fifo_bank_register.bank[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _17878_ (.CLK(net497),
    .D(_01321_),
    .Q(\fifo_bank_register.bank[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _17879_ (.CLK(net532),
    .D(_01322_),
    .Q(\fifo_bank_register.bank[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _17880_ (.CLK(net535),
    .D(_01323_),
    .Q(\fifo_bank_register.bank[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _17881_ (.CLK(net502),
    .D(_01324_),
    .Q(\fifo_bank_register.bank[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _17882_ (.CLK(net513),
    .D(_01325_),
    .Q(\fifo_bank_register.bank[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _17883_ (.CLK(net482),
    .D(_01326_),
    .Q(\fifo_bank_register.bank[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _17884_ (.CLK(net502),
    .D(_01327_),
    .Q(\fifo_bank_register.bank[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _17885_ (.CLK(net483),
    .D(_01328_),
    .Q(\fifo_bank_register.bank[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _17886_ (.CLK(net482),
    .D(_01329_),
    .Q(\fifo_bank_register.bank[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _17887_ (.CLK(net508),
    .D(_01330_),
    .Q(\fifo_bank_register.bank[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _17888_ (.CLK(net510),
    .D(_01331_),
    .Q(\fifo_bank_register.bank[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _17889_ (.CLK(net480),
    .D(_01332_),
    .Q(\fifo_bank_register.bank[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _17890_ (.CLK(net485),
    .D(_01333_),
    .Q(\fifo_bank_register.bank[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _17891_ (.CLK(net492),
    .D(_01334_),
    .Q(\fifo_bank_register.bank[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _17892_ (.CLK(net438),
    .D(_01335_),
    .Q(\fifo_bank_register.bank[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _17893_ (.CLK(net438),
    .D(_01336_),
    .Q(\fifo_bank_register.bank[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _17894_ (.CLK(net418),
    .D(_01337_),
    .Q(\fifo_bank_register.bank[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 _17895_ (.CLK(net425),
    .D(_01338_),
    .Q(\fifo_bank_register.bank[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 _17896_ (.CLK(net431),
    .D(_01339_),
    .Q(\fifo_bank_register.bank[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 _17897_ (.CLK(net429),
    .D(_01340_),
    .Q(\fifo_bank_register.bank[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 _17898_ (.CLK(net425),
    .D(_01341_),
    .Q(\fifo_bank_register.bank[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 _17899_ (.CLK(net417),
    .D(_01342_),
    .Q(\fifo_bank_register.bank[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 _17900_ (.CLK(net428),
    .D(_01343_),
    .Q(\fifo_bank_register.bank[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 _17901_ (.CLK(net415),
    .D(_01344_),
    .Q(\fifo_bank_register.bank[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 _17902_ (.CLK(net395),
    .D(_01345_),
    .Q(\fifo_bank_register.bank[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 _17903_ (.CLK(net398),
    .D(_01346_),
    .Q(\fifo_bank_register.bank[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 _17904_ (.CLK(net399),
    .D(_01347_),
    .Q(\fifo_bank_register.bank[0][42] ));
 sky130_fd_sc_hd__dfxtp_1 _17905_ (.CLK(net393),
    .D(_01348_),
    .Q(\fifo_bank_register.bank[0][43] ));
 sky130_fd_sc_hd__dfxtp_1 _17906_ (.CLK(net389),
    .D(_01349_),
    .Q(\fifo_bank_register.bank[0][44] ));
 sky130_fd_sc_hd__dfxtp_1 _17907_ (.CLK(net406),
    .D(_01350_),
    .Q(\fifo_bank_register.bank[0][45] ));
 sky130_fd_sc_hd__dfxtp_1 _17908_ (.CLK(net390),
    .D(_01351_),
    .Q(\fifo_bank_register.bank[0][46] ));
 sky130_fd_sc_hd__dfxtp_1 _17909_ (.CLK(net396),
    .D(_01352_),
    .Q(\fifo_bank_register.bank[0][47] ));
 sky130_fd_sc_hd__dfxtp_1 _17910_ (.CLK(net396),
    .D(_01353_),
    .Q(\fifo_bank_register.bank[0][48] ));
 sky130_fd_sc_hd__dfxtp_1 _17911_ (.CLK(net408),
    .D(_01354_),
    .Q(\fifo_bank_register.bank[0][49] ));
 sky130_fd_sc_hd__dfxtp_1 _17912_ (.CLK(net557),
    .D(_01355_),
    .Q(\fifo_bank_register.bank[0][50] ));
 sky130_fd_sc_hd__dfxtp_1 _17913_ (.CLK(net575),
    .D(_01356_),
    .Q(\fifo_bank_register.bank[0][51] ));
 sky130_fd_sc_hd__dfxtp_1 _17914_ (.CLK(net567),
    .D(_01357_),
    .Q(\fifo_bank_register.bank[0][52] ));
 sky130_fd_sc_hd__dfxtp_1 _17915_ (.CLK(net567),
    .D(_01358_),
    .Q(\fifo_bank_register.bank[0][53] ));
 sky130_fd_sc_hd__dfxtp_1 _17916_ (.CLK(net555),
    .D(_01359_),
    .Q(\fifo_bank_register.bank[0][54] ));
 sky130_fd_sc_hd__dfxtp_1 _17917_ (.CLK(net575),
    .D(_01360_),
    .Q(\fifo_bank_register.bank[0][55] ));
 sky130_fd_sc_hd__dfxtp_1 _17918_ (.CLK(net574),
    .D(_01361_),
    .Q(\fifo_bank_register.bank[0][56] ));
 sky130_fd_sc_hd__dfxtp_1 _17919_ (.CLK(net549),
    .D(_01362_),
    .Q(\fifo_bank_register.bank[0][57] ));
 sky130_fd_sc_hd__dfxtp_1 _17920_ (.CLK(net557),
    .D(_01363_),
    .Q(\fifo_bank_register.bank[0][58] ));
 sky130_fd_sc_hd__dfxtp_1 _17921_ (.CLK(net573),
    .D(_01364_),
    .Q(\fifo_bank_register.bank[0][59] ));
 sky130_fd_sc_hd__dfxtp_1 _17922_ (.CLK(net513),
    .D(_01365_),
    .Q(\fifo_bank_register.bank[0][60] ));
 sky130_fd_sc_hd__dfxtp_1 _17923_ (.CLK(net527),
    .D(_01366_),
    .Q(\fifo_bank_register.bank[0][61] ));
 sky130_fd_sc_hd__dfxtp_1 _17924_ (.CLK(net523),
    .D(_01367_),
    .Q(\fifo_bank_register.bank[0][62] ));
 sky130_fd_sc_hd__dfxtp_1 _17925_ (.CLK(net524),
    .D(_01368_),
    .Q(\fifo_bank_register.bank[0][63] ));
 sky130_fd_sc_hd__dfxtp_1 _17926_ (.CLK(net512),
    .D(_01369_),
    .Q(\fifo_bank_register.bank[0][64] ));
 sky130_fd_sc_hd__dfxtp_1 _17927_ (.CLK(net526),
    .D(_01370_),
    .Q(\fifo_bank_register.bank[0][65] ));
 sky130_fd_sc_hd__dfxtp_1 _17928_ (.CLK(net527),
    .D(_01371_),
    .Q(\fifo_bank_register.bank[0][66] ));
 sky130_fd_sc_hd__dfxtp_1 _17929_ (.CLK(net514),
    .D(_01372_),
    .Q(\fifo_bank_register.bank[0][67] ));
 sky130_fd_sc_hd__dfxtp_1 _17930_ (.CLK(net511),
    .D(_01373_),
    .Q(\fifo_bank_register.bank[0][68] ));
 sky130_fd_sc_hd__dfxtp_1 _17931_ (.CLK(net516),
    .D(_01374_),
    .Q(\fifo_bank_register.bank[0][69] ));
 sky130_fd_sc_hd__dfxtp_1 _17932_ (.CLK(net519),
    .D(_01375_),
    .Q(\fifo_bank_register.bank[0][70] ));
 sky130_fd_sc_hd__dfxtp_1 _17933_ (.CLK(net528),
    .D(_01376_),
    .Q(\fifo_bank_register.bank[0][71] ));
 sky130_fd_sc_hd__dfxtp_1 _17934_ (.CLK(net554),
    .D(_01377_),
    .Q(\fifo_bank_register.bank[0][72] ));
 sky130_fd_sc_hd__dfxtp_1 _17935_ (.CLK(net554),
    .D(_01378_),
    .Q(\fifo_bank_register.bank[0][73] ));
 sky130_fd_sc_hd__dfxtp_1 _17936_ (.CLK(net549),
    .D(_01379_),
    .Q(\fifo_bank_register.bank[0][74] ));
 sky130_fd_sc_hd__dfxtp_1 _17937_ (.CLK(net552),
    .D(_01380_),
    .Q(\fifo_bank_register.bank[0][75] ));
 sky130_fd_sc_hd__dfxtp_1 _17938_ (.CLK(net545),
    .D(_01381_),
    .Q(\fifo_bank_register.bank[0][76] ));
 sky130_fd_sc_hd__dfxtp_1 _17939_ (.CLK(net555),
    .D(_01382_),
    .Q(\fifo_bank_register.bank[0][77] ));
 sky130_fd_sc_hd__dfxtp_1 _17940_ (.CLK(net525),
    .D(_01383_),
    .Q(\fifo_bank_register.bank[0][78] ));
 sky130_fd_sc_hd__dfxtp_1 _17941_ (.CLK(net549),
    .D(_01384_),
    .Q(\fifo_bank_register.bank[0][79] ));
 sky130_fd_sc_hd__dfxtp_1 _17942_ (.CLK(net566),
    .D(_01385_),
    .Q(\fifo_bank_register.bank[0][80] ));
 sky130_fd_sc_hd__dfxtp_1 _17943_ (.CLK(net565),
    .D(_01386_),
    .Q(\fifo_bank_register.bank[0][81] ));
 sky130_fd_sc_hd__dfxtp_1 _17944_ (.CLK(net562),
    .D(_01387_),
    .Q(\fifo_bank_register.bank[0][82] ));
 sky130_fd_sc_hd__dfxtp_1 _17945_ (.CLK(net563),
    .D(_01388_),
    .Q(\fifo_bank_register.bank[0][83] ));
 sky130_fd_sc_hd__dfxtp_1 _17946_ (.CLK(net536),
    .D(_01389_),
    .Q(\fifo_bank_register.bank[0][84] ));
 sky130_fd_sc_hd__dfxtp_1 _17947_ (.CLK(net568),
    .D(_01390_),
    .Q(\fifo_bank_register.bank[0][85] ));
 sky130_fd_sc_hd__dfxtp_1 _17948_ (.CLK(net538),
    .D(_01391_),
    .Q(\fifo_bank_register.bank[0][86] ));
 sky130_fd_sc_hd__dfxtp_1 _17949_ (.CLK(net564),
    .D(_01392_),
    .Q(\fifo_bank_register.bank[0][87] ));
 sky130_fd_sc_hd__dfxtp_1 _17950_ (.CLK(net541),
    .D(_01393_),
    .Q(\fifo_bank_register.bank[0][88] ));
 sky130_fd_sc_hd__dfxtp_1 _17951_ (.CLK(net547),
    .D(_01394_),
    .Q(\fifo_bank_register.bank[0][89] ));
 sky130_fd_sc_hd__dfxtp_1 _17952_ (.CLK(net406),
    .D(_01395_),
    .Q(\fifo_bank_register.bank[0][90] ));
 sky130_fd_sc_hd__dfxtp_1 _17953_ (.CLK(net403),
    .D(_01396_),
    .Q(\fifo_bank_register.bank[0][91] ));
 sky130_fd_sc_hd__dfxtp_1 _17954_ (.CLK(net410),
    .D(_01397_),
    .Q(\fifo_bank_register.bank[0][92] ));
 sky130_fd_sc_hd__dfxtp_1 _17955_ (.CLK(net399),
    .D(_01398_),
    .Q(\fifo_bank_register.bank[0][93] ));
 sky130_fd_sc_hd__dfxtp_1 _17956_ (.CLK(net455),
    .D(_01399_),
    .Q(\fifo_bank_register.bank[0][94] ));
 sky130_fd_sc_hd__dfxtp_1 _17957_ (.CLK(net402),
    .D(_01400_),
    .Q(\fifo_bank_register.bank[0][95] ));
 sky130_fd_sc_hd__dfxtp_1 _17958_ (.CLK(net403),
    .D(_01401_),
    .Q(\fifo_bank_register.bank[0][96] ));
 sky130_fd_sc_hd__dfxtp_1 _17959_ (.CLK(net455),
    .D(_01402_),
    .Q(\fifo_bank_register.bank[0][97] ));
 sky130_fd_sc_hd__dfxtp_1 _17960_ (.CLK(net447),
    .D(_01403_),
    .Q(\fifo_bank_register.bank[0][98] ));
 sky130_fd_sc_hd__dfxtp_1 _17961_ (.CLK(net447),
    .D(_01404_),
    .Q(\fifo_bank_register.bank[0][99] ));
 sky130_fd_sc_hd__dfxtp_1 _17962_ (.CLK(net452),
    .D(_01405_),
    .Q(\fifo_bank_register.bank[0][100] ));
 sky130_fd_sc_hd__dfxtp_1 _17963_ (.CLK(net450),
    .D(_01406_),
    .Q(\fifo_bank_register.bank[0][101] ));
 sky130_fd_sc_hd__dfxtp_1 _17964_ (.CLK(net466),
    .D(_01407_),
    .Q(\fifo_bank_register.bank[0][102] ));
 sky130_fd_sc_hd__dfxtp_1 _17965_ (.CLK(net467),
    .D(_01408_),
    .Q(\fifo_bank_register.bank[0][103] ));
 sky130_fd_sc_hd__dfxtp_1 _17966_ (.CLK(net463),
    .D(_01409_),
    .Q(\fifo_bank_register.bank[0][104] ));
 sky130_fd_sc_hd__dfxtp_1 _17967_ (.CLK(net467),
    .D(_01410_),
    .Q(\fifo_bank_register.bank[0][105] ));
 sky130_fd_sc_hd__dfxtp_1 _17968_ (.CLK(net465),
    .D(_01411_),
    .Q(\fifo_bank_register.bank[0][106] ));
 sky130_fd_sc_hd__dfxtp_1 _17969_ (.CLK(net451),
    .D(_01412_),
    .Q(\fifo_bank_register.bank[0][107] ));
 sky130_fd_sc_hd__dfxtp_1 _17970_ (.CLK(net452),
    .D(_01413_),
    .Q(\fifo_bank_register.bank[0][108] ));
 sky130_fd_sc_hd__dfxtp_1 _17971_ (.CLK(net458),
    .D(_01414_),
    .Q(\fifo_bank_register.bank[0][109] ));
 sky130_fd_sc_hd__dfxtp_1 _17972_ (.CLK(net434),
    .D(_01415_),
    .Q(\fifo_bank_register.bank[0][110] ));
 sky130_fd_sc_hd__dfxtp_1 _17973_ (.CLK(net411),
    .D(_01416_),
    .Q(\fifo_bank_register.bank[0][111] ));
 sky130_fd_sc_hd__dfxtp_1 _17974_ (.CLK(net433),
    .D(_01417_),
    .Q(\fifo_bank_register.bank[0][112] ));
 sky130_fd_sc_hd__dfxtp_1 _17975_ (.CLK(net469),
    .D(_01418_),
    .Q(\fifo_bank_register.bank[0][113] ));
 sky130_fd_sc_hd__dfxtp_1 _17976_ (.CLK(net457),
    .D(_01419_),
    .Q(\fifo_bank_register.bank[0][114] ));
 sky130_fd_sc_hd__dfxtp_1 _17977_ (.CLK(net470),
    .D(_01420_),
    .Q(\fifo_bank_register.bank[0][115] ));
 sky130_fd_sc_hd__dfxtp_1 _17978_ (.CLK(net456),
    .D(_01421_),
    .Q(\fifo_bank_register.bank[0][116] ));
 sky130_fd_sc_hd__dfxtp_1 _17979_ (.CLK(net435),
    .D(_01422_),
    .Q(\fifo_bank_register.bank[0][117] ));
 sky130_fd_sc_hd__dfxtp_1 _17980_ (.CLK(net457),
    .D(_01423_),
    .Q(\fifo_bank_register.bank[0][118] ));
 sky130_fd_sc_hd__dfxtp_1 _17981_ (.CLK(net435),
    .D(_01424_),
    .Q(\fifo_bank_register.bank[0][119] ));
 sky130_fd_sc_hd__dfxtp_1 _17982_ (.CLK(net472),
    .D(_01425_),
    .Q(\fifo_bank_register.bank[0][120] ));
 sky130_fd_sc_hd__dfxtp_1 _17983_ (.CLK(net491),
    .D(_01426_),
    .Q(\fifo_bank_register.bank[0][121] ));
 sky130_fd_sc_hd__dfxtp_1 _17984_ (.CLK(net491),
    .D(_01427_),
    .Q(\fifo_bank_register.bank[0][122] ));
 sky130_fd_sc_hd__dfxtp_1 _17985_ (.CLK(net437),
    .D(_01428_),
    .Q(\fifo_bank_register.bank[0][123] ));
 sky130_fd_sc_hd__dfxtp_1 _17986_ (.CLK(net531),
    .D(_01429_),
    .Q(\fifo_bank_register.bank[0][124] ));
 sky130_fd_sc_hd__dfxtp_1 _17987_ (.CLK(net531),
    .D(_01430_),
    .Q(\fifo_bank_register.bank[0][125] ));
 sky130_fd_sc_hd__dfxtp_1 _17988_ (.CLK(net531),
    .D(_01431_),
    .Q(\fifo_bank_register.bank[0][126] ));
 sky130_fd_sc_hd__dfxtp_1 _17989_ (.CLK(net443),
    .D(_01432_),
    .Q(\fifo_bank_register.bank[0][127] ));
 sky130_fd_sc_hd__dfrtp_4 _17990_ (.CLK(net442),
    .D(_01433_),
    .RESET_B(net596),
    .Q(\fifo_bank_register.read_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _17991_ (.CLK(net438),
    .D(_01434_),
    .RESET_B(net597),
    .Q(\fifo_bank_register.read_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 _17992_ (.CLK(net437),
    .D(_01435_),
    .RESET_B(net597),
    .Q(\fifo_bank_register.read_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_2 _17993_ (.CLK(net442),
    .D(_01436_),
    .RESET_B(net597),
    .Q(\fifo_bank_register.read_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_1 _17994_ (.CLK(net442),
    .D(_01437_),
    .RESET_B(net597),
    .Q(\fifo_bank_register.write_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 _17995_ (.CLK(net442),
    .D(_01438_),
    .RESET_B(net602),
    .Q(\fifo_bank_register.write_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _17996_ (.CLK(net442),
    .D(_01439_),
    .RESET_B(net596),
    .Q(\fifo_bank_register.write_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _17997_ (.CLK(net434),
    .D(_01440_),
    .RESET_B(net596),
    .Q(\fifo_bank_register.write_ptr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _17998_ (.CLK(net421),
    .D(_01441_),
    .Q(\fifo_bank_register.data_out[0] ));
 sky130_fd_sc_hd__dfxtp_4 _17999_ (.CLK(net440),
    .D(_01442_),
    .Q(\fifo_bank_register.data_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _18000_ (.CLK(net420),
    .D(_01443_),
    .Q(\fifo_bank_register.data_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _18001_ (.CLK(net420),
    .D(_01444_),
    .Q(\fifo_bank_register.data_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _18002_ (.CLK(net422),
    .D(_01445_),
    .Q(\fifo_bank_register.data_out[4] ));
 sky130_fd_sc_hd__dfxtp_4 _18003_ (.CLK(net420),
    .D(_01446_),
    .Q(\fifo_bank_register.data_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _18004_ (.CLK(net425),
    .D(_01447_),
    .Q(\fifo_bank_register.data_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _18005_ (.CLK(net425),
    .D(_01448_),
    .Q(\fifo_bank_register.data_out[7] ));
 sky130_fd_sc_hd__dfxtp_2 _18006_ (.CLK(net426),
    .D(_01449_),
    .Q(\fifo_bank_register.data_out[8] ));
 sky130_fd_sc_hd__dfxtp_1 _18007_ (.CLK(net426),
    .D(_01450_),
    .Q(\fifo_bank_register.data_out[9] ));
 sky130_fd_sc_hd__dfxtp_1 _18008_ (.CLK(net493),
    .D(_01451_),
    .Q(\fifo_bank_register.data_out[10] ));
 sky130_fd_sc_hd__dfxtp_1 _18009_ (.CLK(net535),
    .D(_01452_),
    .Q(\fifo_bank_register.data_out[11] ));
 sky130_fd_sc_hd__dfxtp_1 _18010_ (.CLK(net500),
    .D(_01453_),
    .Q(\fifo_bank_register.data_out[12] ));
 sky130_fd_sc_hd__dfxtp_2 _18011_ (.CLK(net506),
    .D(_01454_),
    .Q(\fifo_bank_register.data_out[13] ));
 sky130_fd_sc_hd__dfxtp_1 _18012_ (.CLK(net534),
    .D(_01455_),
    .Q(\fifo_bank_register.data_out[14] ));
 sky130_fd_sc_hd__dfxtp_1 _18013_ (.CLK(net535),
    .D(_01456_),
    .Q(\fifo_bank_register.data_out[15] ));
 sky130_fd_sc_hd__dfxtp_4 _18014_ (.CLK(net471),
    .D(_01457_),
    .Q(\fifo_bank_register.data_out[16] ));
 sky130_fd_sc_hd__dfxtp_2 _18015_ (.CLK(net531),
    .D(_01458_),
    .Q(\fifo_bank_register.data_out[17] ));
 sky130_fd_sc_hd__dfxtp_2 _18016_ (.CLK(net533),
    .D(_01459_),
    .Q(\fifo_bank_register.data_out[18] ));
 sky130_fd_sc_hd__dfxtp_1 _18017_ (.CLK(net502),
    .D(_01460_),
    .Q(\fifo_bank_register.data_out[19] ));
 sky130_fd_sc_hd__dfxtp_4 _18018_ (.CLK(net516),
    .D(_01461_),
    .Q(\fifo_bank_register.data_out[20] ));
 sky130_fd_sc_hd__dfxtp_1 _18019_ (.CLK(net482),
    .D(_01462_),
    .Q(\fifo_bank_register.data_out[21] ));
 sky130_fd_sc_hd__dfxtp_2 _18020_ (.CLK(net513),
    .D(_01463_),
    .Q(\fifo_bank_register.data_out[22] ));
 sky130_fd_sc_hd__dfxtp_1 _18021_ (.CLK(net483),
    .D(_01464_),
    .Q(\fifo_bank_register.data_out[23] ));
 sky130_fd_sc_hd__dfxtp_1 _18022_ (.CLK(net482),
    .D(_01465_),
    .Q(\fifo_bank_register.data_out[24] ));
 sky130_fd_sc_hd__dfxtp_1 _18023_ (.CLK(net513),
    .D(_01466_),
    .Q(\fifo_bank_register.data_out[25] ));
 sky130_fd_sc_hd__dfxtp_1 _18024_ (.CLK(net510),
    .D(_01467_),
    .Q(\fifo_bank_register.data_out[26] ));
 sky130_fd_sc_hd__dfxtp_2 _18025_ (.CLK(net426),
    .D(_01468_),
    .Q(\fifo_bank_register.data_out[27] ));
 sky130_fd_sc_hd__dfxtp_1 _18026_ (.CLK(net485),
    .D(_01469_),
    .Q(\fifo_bank_register.data_out[28] ));
 sky130_fd_sc_hd__dfxtp_1 _18027_ (.CLK(net480),
    .D(_01470_),
    .Q(\fifo_bank_register.data_out[29] ));
 sky130_fd_sc_hd__dfxtp_4 _18028_ (.CLK(net438),
    .D(_01471_),
    .Q(\fifo_bank_register.data_out[30] ));
 sky130_fd_sc_hd__dfxtp_1 _18029_ (.CLK(net438),
    .D(_01472_),
    .Q(\fifo_bank_register.data_out[31] ));
 sky130_fd_sc_hd__dfxtp_1 _18030_ (.CLK(net416),
    .D(_01473_),
    .Q(\fifo_bank_register.data_out[32] ));
 sky130_fd_sc_hd__dfxtp_1 _18031_ (.CLK(net426),
    .D(_01474_),
    .Q(\fifo_bank_register.data_out[33] ));
 sky130_fd_sc_hd__dfxtp_1 _18032_ (.CLK(net431),
    .D(_01475_),
    .Q(\fifo_bank_register.data_out[34] ));
 sky130_fd_sc_hd__dfxtp_4 _18033_ (.CLK(net429),
    .D(_01476_),
    .Q(\fifo_bank_register.data_out[35] ));
 sky130_fd_sc_hd__dfxtp_1 _18034_ (.CLK(net425),
    .D(_01477_),
    .Q(\fifo_bank_register.data_out[36] ));
 sky130_fd_sc_hd__dfxtp_4 _18035_ (.CLK(net415),
    .D(_01478_),
    .Q(\fifo_bank_register.data_out[37] ));
 sky130_fd_sc_hd__dfxtp_4 _18036_ (.CLK(net407),
    .D(_01479_),
    .Q(\fifo_bank_register.data_out[38] ));
 sky130_fd_sc_hd__dfxtp_1 _18037_ (.CLK(net415),
    .D(_01480_),
    .Q(\fifo_bank_register.data_out[39] ));
 sky130_fd_sc_hd__dfxtp_1 _18038_ (.CLK(net415),
    .D(_01481_),
    .Q(\fifo_bank_register.data_out[40] ));
 sky130_fd_sc_hd__dfxtp_2 _18039_ (.CLK(net399),
    .D(_01482_),
    .Q(\fifo_bank_register.data_out[41] ));
 sky130_fd_sc_hd__dfxtp_2 _18040_ (.CLK(net399),
    .D(_01483_),
    .Q(\fifo_bank_register.data_out[42] ));
 sky130_fd_sc_hd__dfxtp_2 _18041_ (.CLK(net407),
    .D(_01484_),
    .Q(\fifo_bank_register.data_out[43] ));
 sky130_fd_sc_hd__dfxtp_1 _18042_ (.CLK(net389),
    .D(_01485_),
    .Q(\fifo_bank_register.data_out[44] ));
 sky130_fd_sc_hd__dfxtp_1 _18043_ (.CLK(net406),
    .D(_01486_),
    .Q(\fifo_bank_register.data_out[45] ));
 sky130_fd_sc_hd__dfxtp_1 _18044_ (.CLK(net390),
    .D(_01487_),
    .Q(\fifo_bank_register.data_out[46] ));
 sky130_fd_sc_hd__dfxtp_1 _18045_ (.CLK(net395),
    .D(_01488_),
    .Q(\fifo_bank_register.data_out[47] ));
 sky130_fd_sc_hd__dfxtp_1 _18046_ (.CLK(net415),
    .D(_01489_),
    .Q(\fifo_bank_register.data_out[48] ));
 sky130_fd_sc_hd__dfxtp_4 _18047_ (.CLK(net429),
    .D(_01490_),
    .Q(\fifo_bank_register.data_out[49] ));
 sky130_fd_sc_hd__dfxtp_1 _18048_ (.CLK(net557),
    .D(_01491_),
    .Q(\fifo_bank_register.data_out[50] ));
 sky130_fd_sc_hd__dfxtp_1 _18049_ (.CLK(net574),
    .D(_01492_),
    .Q(\fifo_bank_register.data_out[51] ));
 sky130_fd_sc_hd__dfxtp_2 _18050_ (.CLK(net567),
    .D(_01493_),
    .Q(\fifo_bank_register.data_out[52] ));
 sky130_fd_sc_hd__dfxtp_2 _18051_ (.CLK(net568),
    .D(_01494_),
    .Q(\fifo_bank_register.data_out[53] ));
 sky130_fd_sc_hd__dfxtp_2 _18052_ (.CLK(net555),
    .D(_01495_),
    .Q(\fifo_bank_register.data_out[54] ));
 sky130_fd_sc_hd__dfxtp_1 _18053_ (.CLK(net574),
    .D(_01496_),
    .Q(\fifo_bank_register.data_out[55] ));
 sky130_fd_sc_hd__dfxtp_4 _18054_ (.CLK(net574),
    .D(_01497_),
    .Q(\fifo_bank_register.data_out[56] ));
 sky130_fd_sc_hd__dfxtp_1 _18055_ (.CLK(net549),
    .D(_01498_),
    .Q(\fifo_bank_register.data_out[57] ));
 sky130_fd_sc_hd__dfxtp_1 _18056_ (.CLK(net557),
    .D(_01499_),
    .Q(\fifo_bank_register.data_out[58] ));
 sky130_fd_sc_hd__dfxtp_2 _18057_ (.CLK(net574),
    .D(_01500_),
    .Q(\fifo_bank_register.data_out[59] ));
 sky130_fd_sc_hd__dfxtp_1 _18058_ (.CLK(net513),
    .D(_01501_),
    .Q(\fifo_bank_register.data_out[60] ));
 sky130_fd_sc_hd__dfxtp_1 _18059_ (.CLK(net528),
    .D(_01502_),
    .Q(\fifo_bank_register.data_out[61] ));
 sky130_fd_sc_hd__dfxtp_1 _18060_ (.CLK(net523),
    .D(_01503_),
    .Q(\fifo_bank_register.data_out[62] ));
 sky130_fd_sc_hd__dfxtp_1 _18061_ (.CLK(net575),
    .D(_01504_),
    .Q(\fifo_bank_register.data_out[63] ));
 sky130_fd_sc_hd__dfxtp_2 _18062_ (.CLK(net512),
    .D(_01505_),
    .Q(\fifo_bank_register.data_out[64] ));
 sky130_fd_sc_hd__dfxtp_2 _18063_ (.CLK(net567),
    .D(_01506_),
    .Q(\fifo_bank_register.data_out[65] ));
 sky130_fd_sc_hd__dfxtp_1 _18064_ (.CLK(net573),
    .D(_01507_),
    .Q(\fifo_bank_register.data_out[66] ));
 sky130_fd_sc_hd__dfxtp_1 _18065_ (.CLK(net508),
    .D(_01508_),
    .Q(\fifo_bank_register.data_out[67] ));
 sky130_fd_sc_hd__dfxtp_1 _18066_ (.CLK(net509),
    .D(_01509_),
    .Q(\fifo_bank_register.data_out[68] ));
 sky130_fd_sc_hd__dfxtp_2 _18067_ (.CLK(net516),
    .D(_01510_),
    .Q(\fifo_bank_register.data_out[69] ));
 sky130_fd_sc_hd__dfxtp_1 _18068_ (.CLK(net516),
    .D(_01511_),
    .Q(\fifo_bank_register.data_out[70] ));
 sky130_fd_sc_hd__dfxtp_1 _18069_ (.CLK(net527),
    .D(_01512_),
    .Q(\fifo_bank_register.data_out[71] ));
 sky130_fd_sc_hd__dfxtp_1 _18070_ (.CLK(net557),
    .D(_01513_),
    .Q(\fifo_bank_register.data_out[72] ));
 sky130_fd_sc_hd__dfxtp_1 _18071_ (.CLK(net554),
    .D(_01514_),
    .Q(\fifo_bank_register.data_out[73] ));
 sky130_fd_sc_hd__dfxtp_2 _18072_ (.CLK(net549),
    .D(_01515_),
    .Q(\fifo_bank_register.data_out[74] ));
 sky130_fd_sc_hd__dfxtp_1 _18073_ (.CLK(net555),
    .D(_01516_),
    .Q(\fifo_bank_register.data_out[75] ));
 sky130_fd_sc_hd__dfxtp_2 _18074_ (.CLK(net516),
    .D(_01517_),
    .Q(\fifo_bank_register.data_out[76] ));
 sky130_fd_sc_hd__dfxtp_1 _18075_ (.CLK(net555),
    .D(_01518_),
    .Q(\fifo_bank_register.data_out[77] ));
 sky130_fd_sc_hd__dfxtp_1 _18076_ (.CLK(net519),
    .D(_01519_),
    .Q(\fifo_bank_register.data_out[78] ));
 sky130_fd_sc_hd__dfxtp_1 _18077_ (.CLK(net568),
    .D(_01520_),
    .Q(\fifo_bank_register.data_out[79] ));
 sky130_fd_sc_hd__dfxtp_2 _18078_ (.CLK(net566),
    .D(_01521_),
    .Q(\fifo_bank_register.data_out[80] ));
 sky130_fd_sc_hd__dfxtp_1 _18079_ (.CLK(net566),
    .D(_01522_),
    .Q(\fifo_bank_register.data_out[81] ));
 sky130_fd_sc_hd__dfxtp_1 _18080_ (.CLK(net568),
    .D(_01523_),
    .Q(\fifo_bank_register.data_out[82] ));
 sky130_fd_sc_hd__dfxtp_1 _18081_ (.CLK(net568),
    .D(_01524_),
    .Q(\fifo_bank_register.data_out[83] ));
 sky130_fd_sc_hd__dfxtp_2 _18082_ (.CLK(net537),
    .D(_01525_),
    .Q(\fifo_bank_register.data_out[84] ));
 sky130_fd_sc_hd__dfxtp_1 _18083_ (.CLK(net568),
    .D(_01526_),
    .Q(\fifo_bank_register.data_out[85] ));
 sky130_fd_sc_hd__dfxtp_2 _18084_ (.CLK(net560),
    .D(_01527_),
    .Q(\fifo_bank_register.data_out[86] ));
 sky130_fd_sc_hd__dfxtp_2 _18085_ (.CLK(net542),
    .D(_01528_),
    .Q(\fifo_bank_register.data_out[87] ));
 sky130_fd_sc_hd__dfxtp_2 _18086_ (.CLK(net541),
    .D(_01529_),
    .Q(\fifo_bank_register.data_out[88] ));
 sky130_fd_sc_hd__dfxtp_1 _18087_ (.CLK(net472),
    .D(_01530_),
    .Q(\fifo_bank_register.data_out[89] ));
 sky130_fd_sc_hd__dfxtp_1 _18088_ (.CLK(net405),
    .D(_01531_),
    .Q(\fifo_bank_register.data_out[90] ));
 sky130_fd_sc_hd__dfxtp_1 _18089_ (.CLK(net472),
    .D(_01532_),
    .Q(\fifo_bank_register.data_out[91] ));
 sky130_fd_sc_hd__dfxtp_2 _18090_ (.CLK(net456),
    .D(_01533_),
    .Q(\fifo_bank_register.data_out[92] ));
 sky130_fd_sc_hd__dfxtp_1 _18091_ (.CLK(net434),
    .D(_01534_),
    .Q(\fifo_bank_register.data_out[93] ));
 sky130_fd_sc_hd__dfxtp_1 _18092_ (.CLK(net460),
    .D(_01535_),
    .Q(\fifo_bank_register.data_out[94] ));
 sky130_fd_sc_hd__dfxtp_1 _18093_ (.CLK(net399),
    .D(_01536_),
    .Q(\fifo_bank_register.data_out[95] ));
 sky130_fd_sc_hd__dfxtp_1 _18094_ (.CLK(net398),
    .D(_01537_),
    .Q(\fifo_bank_register.data_out[96] ));
 sky130_fd_sc_hd__dfxtp_1 _18095_ (.CLK(net457),
    .D(_01538_),
    .Q(\fifo_bank_register.data_out[97] ));
 sky130_fd_sc_hd__dfxtp_1 _18096_ (.CLK(net458),
    .D(_01539_),
    .Q(\fifo_bank_register.data_out[98] ));
 sky130_fd_sc_hd__dfxtp_1 _18097_ (.CLK(net463),
    .D(_01540_),
    .Q(\fifo_bank_register.data_out[99] ));
 sky130_fd_sc_hd__dfxtp_1 _18098_ (.CLK(net458),
    .D(_01541_),
    .Q(\fifo_bank_register.data_out[100] ));
 sky130_fd_sc_hd__dfxtp_1 _18099_ (.CLK(net450),
    .D(_01542_),
    .Q(\fifo_bank_register.data_out[101] ));
 sky130_fd_sc_hd__dfxtp_1 _18100_ (.CLK(net466),
    .D(_01543_),
    .Q(\fifo_bank_register.data_out[102] ));
 sky130_fd_sc_hd__dfxtp_1 _18101_ (.CLK(net459),
    .D(_01544_),
    .Q(\fifo_bank_register.data_out[103] ));
 sky130_fd_sc_hd__dfxtp_2 _18102_ (.CLK(net466),
    .D(_01545_),
    .Q(\fifo_bank_register.data_out[104] ));
 sky130_fd_sc_hd__dfxtp_1 _18103_ (.CLK(net468),
    .D(_01546_),
    .Q(\fifo_bank_register.data_out[105] ));
 sky130_fd_sc_hd__dfxtp_1 _18104_ (.CLK(net466),
    .D(_01547_),
    .Q(\fifo_bank_register.data_out[106] ));
 sky130_fd_sc_hd__dfxtp_1 _18105_ (.CLK(net451),
    .D(_01548_),
    .Q(\fifo_bank_register.data_out[107] ));
 sky130_fd_sc_hd__dfxtp_1 _18106_ (.CLK(net450),
    .D(_01549_),
    .Q(\fifo_bank_register.data_out[108] ));
 sky130_fd_sc_hd__dfxtp_2 _18107_ (.CLK(net459),
    .D(_01550_),
    .Q(\fifo_bank_register.data_out[109] ));
 sky130_fd_sc_hd__dfxtp_2 _18108_ (.CLK(net470),
    .D(_01551_),
    .Q(\fifo_bank_register.data_out[110] ));
 sky130_fd_sc_hd__dfxtp_2 _18109_ (.CLK(net454),
    .D(_01552_),
    .Q(\fifo_bank_register.data_out[111] ));
 sky130_fd_sc_hd__dfxtp_1 _18110_ (.CLK(net470),
    .D(_01553_),
    .Q(\fifo_bank_register.data_out[112] ));
 sky130_fd_sc_hd__dfxtp_1 _18111_ (.CLK(net470),
    .D(_01554_),
    .Q(\fifo_bank_register.data_out[113] ));
 sky130_fd_sc_hd__dfxtp_2 _18112_ (.CLK(net454),
    .D(_01555_),
    .Q(\fifo_bank_register.data_out[114] ));
 sky130_fd_sc_hd__dfxtp_4 _18113_ (.CLK(net471),
    .D(_01556_),
    .Q(\fifo_bank_register.data_out[115] ));
 sky130_fd_sc_hd__dfxtp_1 _18114_ (.CLK(net457),
    .D(_01557_),
    .Q(\fifo_bank_register.data_out[116] ));
 sky130_fd_sc_hd__dfxtp_1 _18115_ (.CLK(net442),
    .D(_01558_),
    .Q(\fifo_bank_register.data_out[117] ));
 sky130_fd_sc_hd__dfxtp_2 _18116_ (.CLK(net457),
    .D(_01559_),
    .Q(\fifo_bank_register.data_out[118] ));
 sky130_fd_sc_hd__dfxtp_1 _18117_ (.CLK(net431),
    .D(_01560_),
    .Q(\fifo_bank_register.data_out[119] ));
 sky130_fd_sc_hd__dfxtp_2 _18118_ (.CLK(net471),
    .D(_01561_),
    .Q(\fifo_bank_register.data_out[120] ));
 sky130_fd_sc_hd__dfxtp_1 _18119_ (.CLK(net490),
    .D(_01562_),
    .Q(\fifo_bank_register.data_out[121] ));
 sky130_fd_sc_hd__dfxtp_1 _18120_ (.CLK(net428),
    .D(_01563_),
    .Q(\fifo_bank_register.data_out[122] ));
 sky130_fd_sc_hd__dfxtp_1 _18121_ (.CLK(net428),
    .D(_01564_),
    .Q(\fifo_bank_register.data_out[123] ));
 sky130_fd_sc_hd__dfxtp_1 _18122_ (.CLK(net531),
    .D(_01565_),
    .Q(\fifo_bank_register.data_out[124] ));
 sky130_fd_sc_hd__dfxtp_1 _18123_ (.CLK(net531),
    .D(_01566_),
    .Q(\fifo_bank_register.data_out[125] ));
 sky130_fd_sc_hd__dfxtp_1 _18124_ (.CLK(net531),
    .D(_01567_),
    .Q(\fifo_bank_register.data_out[126] ));
 sky130_fd_sc_hd__dfxtp_1 _18125_ (.CLK(net442),
    .D(_01568_),
    .Q(\fifo_bank_register.data_out[127] ));
 sky130_fd_sc_hd__dfrtp_4 _18126_ (.CLK(clknet_leaf_20_clk),
    .D(_01569_),
    .RESET_B(net640),
    .Q(\sub1.data_o[80] ));
 sky130_fd_sc_hd__dfrtp_4 _18127_ (.CLK(clknet_leaf_20_clk),
    .D(_01570_),
    .RESET_B(net640),
    .Q(\sub1.data_o[81] ));
 sky130_fd_sc_hd__dfrtp_4 _18128_ (.CLK(clknet_leaf_21_clk),
    .D(_01571_),
    .RESET_B(net639),
    .Q(\sub1.data_o[82] ));
 sky130_fd_sc_hd__dfrtp_4 _18129_ (.CLK(clknet_leaf_24_clk),
    .D(_01572_),
    .RESET_B(net643),
    .Q(\sub1.data_o[83] ));
 sky130_fd_sc_hd__dfrtp_4 _18130_ (.CLK(clknet_leaf_28_clk),
    .D(_01573_),
    .RESET_B(net641),
    .Q(\sub1.data_o[84] ));
 sky130_fd_sc_hd__dfrtp_4 _18131_ (.CLK(clknet_leaf_22_clk),
    .D(_01574_),
    .RESET_B(net643),
    .Q(\sub1.data_o[85] ));
 sky130_fd_sc_hd__dfrtp_4 _18132_ (.CLK(clknet_leaf_24_clk),
    .D(_01575_),
    .RESET_B(net643),
    .Q(\sub1.data_o[86] ));
 sky130_fd_sc_hd__dfrtp_4 _18133_ (.CLK(clknet_leaf_28_clk),
    .D(_01576_),
    .RESET_B(net643),
    .Q(\sub1.data_o[87] ));
 sky130_fd_sc_hd__dfrtp_2 _18134_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.intermediate_to_invert_var[0] ),
    .RESET_B(net656),
    .Q(\sbox1.inversion_to_invert_var[0] ));
 sky130_fd_sc_hd__dfrtp_4 _18135_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.intermediate_to_invert_var[1] ),
    .RESET_B(net656),
    .Q(\sbox1.inversion_to_invert_var[1] ));
 sky130_fd_sc_hd__dfrtp_1 _18136_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.intermediate_to_invert_var[2] ),
    .RESET_B(net656),
    .Q(\sbox1.inversion_to_invert_var[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18137_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.intermediate_to_invert_var[3] ),
    .RESET_B(net656),
    .Q(\sbox1.inversion_to_invert_var[3] ));
 sky130_fd_sc_hd__dfrtp_2 _18138_ (.CLK(clknet_leaf_42_clk),
    .D(\sbox1.next_alph[0] ),
    .RESET_B(net656),
    .Q(\sbox1.alph[0] ));
 sky130_fd_sc_hd__dfrtp_1 _18139_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.next_alph[1] ),
    .RESET_B(net656),
    .Q(\sbox1.alph[1] ));
 sky130_fd_sc_hd__dfrtp_1 _18140_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.next_alph[2] ),
    .RESET_B(net657),
    .Q(\sbox1.alph[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18141_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.next_alph[3] ),
    .RESET_B(net657),
    .Q(\sbox1.alph[3] ));
 sky130_fd_sc_hd__dfrtp_1 _18142_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.ah[0] ),
    .RESET_B(net656),
    .Q(\sbox1.ah_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _18143_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.ah[1] ),
    .RESET_B(net657),
    .Q(\sbox1.ah_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 _18144_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.ah[2] ),
    .RESET_B(net656),
    .Q(\sbox1.ah_reg[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18145_ (.CLK(clknet_leaf_53_clk),
    .D(\sbox1.ah[3] ),
    .RESET_B(net656),
    .Q(\sbox1.ah_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _18146_ (.CLK(clknet_leaf_64_clk),
    .D(_01577_),
    .RESET_B(net603),
    .Q(\ks1.col[0] ));
 sky130_fd_sc_hd__dfrtp_2 _18147_ (.CLK(clknet_leaf_78_clk),
    .D(_01578_),
    .RESET_B(net579),
    .Q(\ks1.col[1] ));
 sky130_fd_sc_hd__dfrtp_4 _18148_ (.CLK(clknet_leaf_82_clk),
    .D(_01579_),
    .RESET_B(net587),
    .Q(\ks1.col[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18149_ (.CLK(clknet_leaf_82_clk),
    .D(_01580_),
    .RESET_B(net585),
    .Q(\ks1.col[3] ));
 sky130_fd_sc_hd__dfrtp_2 _18150_ (.CLK(clknet_leaf_81_clk),
    .D(_01581_),
    .RESET_B(net586),
    .Q(\ks1.col[4] ));
 sky130_fd_sc_hd__dfrtp_4 _18151_ (.CLK(clknet_leaf_81_clk),
    .D(_01582_),
    .RESET_B(net578),
    .Q(\ks1.col[5] ));
 sky130_fd_sc_hd__dfrtp_2 _18152_ (.CLK(clknet_leaf_81_clk),
    .D(_01583_),
    .RESET_B(net586),
    .Q(\ks1.col[6] ));
 sky130_fd_sc_hd__dfrtp_4 _18153_ (.CLK(clknet_leaf_81_clk),
    .D(_01584_),
    .RESET_B(net578),
    .Q(\ks1.col[7] ));
 sky130_fd_sc_hd__dfrtp_1 _18154_ (.CLK(clknet_leaf_49_clk),
    .D(_01585_),
    .RESET_B(net615),
    .Q(\ks1.col[24] ));
 sky130_fd_sc_hd__dfrtp_4 _18155_ (.CLK(clknet_leaf_48_clk),
    .D(_01586_),
    .RESET_B(net610),
    .Q(\ks1.col[25] ));
 sky130_fd_sc_hd__dfrtp_2 _18156_ (.CLK(clknet_leaf_67_clk),
    .D(_01587_),
    .RESET_B(net610),
    .Q(\ks1.col[26] ));
 sky130_fd_sc_hd__dfrtp_2 _18157_ (.CLK(clknet_leaf_67_clk),
    .D(_01588_),
    .RESET_B(net606),
    .Q(\ks1.col[27] ));
 sky130_fd_sc_hd__dfrtp_4 _18158_ (.CLK(clknet_leaf_49_clk),
    .D(_01589_),
    .RESET_B(net616),
    .Q(\ks1.col[28] ));
 sky130_fd_sc_hd__dfrtp_2 _18159_ (.CLK(clknet_leaf_48_clk),
    .D(_01590_),
    .RESET_B(net610),
    .Q(\ks1.col[29] ));
 sky130_fd_sc_hd__dfrtp_2 _18160_ (.CLK(clknet_leaf_48_clk),
    .D(_01591_),
    .RESET_B(net612),
    .Q(\ks1.col[30] ));
 sky130_fd_sc_hd__dfrtp_2 _18161_ (.CLK(clknet_leaf_49_clk),
    .D(_01592_),
    .RESET_B(net611),
    .Q(\ks1.col[31] ));
 sky130_fd_sc_hd__dfrtp_1 _18162_ (.CLK(clknet_leaf_81_clk),
    .D(_01593_),
    .RESET_B(net578),
    .Q(\ks1.col[16] ));
 sky130_fd_sc_hd__dfrtp_4 _18163_ (.CLK(clknet_leaf_76_clk),
    .D(_01594_),
    .RESET_B(net589),
    .Q(\ks1.col[17] ));
 sky130_fd_sc_hd__dfrtp_4 _18164_ (.CLK(clknet_leaf_82_clk),
    .D(_01595_),
    .RESET_B(net587),
    .Q(\ks1.col[18] ));
 sky130_fd_sc_hd__dfrtp_2 _18165_ (.CLK(clknet_leaf_75_clk),
    .D(_01596_),
    .RESET_B(net587),
    .Q(\ks1.col[19] ));
 sky130_fd_sc_hd__dfrtp_4 _18166_ (.CLK(clknet_leaf_81_clk),
    .D(_01597_),
    .RESET_B(net586),
    .Q(\ks1.col[20] ));
 sky130_fd_sc_hd__dfrtp_1 _18167_ (.CLK(clknet_leaf_81_clk),
    .D(_01598_),
    .RESET_B(net588),
    .Q(\ks1.col[21] ));
 sky130_fd_sc_hd__dfrtp_1 _18168_ (.CLK(clknet_leaf_4_clk),
    .D(_01599_),
    .RESET_B(net591),
    .Q(\ks1.col[22] ));
 sky130_fd_sc_hd__dfrtp_1 _18169_ (.CLK(clknet_leaf_77_clk),
    .D(_01600_),
    .RESET_B(net589),
    .Q(\ks1.col[23] ));
 sky130_fd_sc_hd__dfrtp_1 _18170_ (.CLK(clknet_leaf_11_clk),
    .D(_01601_),
    .RESET_B(net631),
    .Q(\mix1.data_reg[64] ));
 sky130_fd_sc_hd__dfrtp_1 _18171_ (.CLK(clknet_leaf_17_clk),
    .D(_01602_),
    .RESET_B(net633),
    .Q(\mix1.data_reg[65] ));
 sky130_fd_sc_hd__dfrtp_1 _18172_ (.CLK(clknet_leaf_20_clk),
    .D(_01603_),
    .RESET_B(net640),
    .Q(\mix1.data_reg[66] ));
 sky130_fd_sc_hd__dfrtp_1 _18173_ (.CLK(clknet_leaf_20_clk),
    .D(_01604_),
    .RESET_B(net640),
    .Q(\mix1.data_reg[67] ));
 sky130_fd_sc_hd__dfrtp_1 _18174_ (.CLK(clknet_leaf_20_clk),
    .D(_01605_),
    .RESET_B(net640),
    .Q(\mix1.data_reg[68] ));
 sky130_fd_sc_hd__dfrtp_1 _18175_ (.CLK(clknet_leaf_12_clk),
    .D(_01606_),
    .RESET_B(net627),
    .Q(\mix1.data_reg[69] ));
 sky130_fd_sc_hd__dfrtp_1 _18176_ (.CLK(clknet_leaf_13_clk),
    .D(_01607_),
    .RESET_B(net627),
    .Q(\mix1.data_reg[70] ));
 sky130_fd_sc_hd__dfrtp_1 _18177_ (.CLK(clknet_leaf_13_clk),
    .D(_01608_),
    .RESET_B(net627),
    .Q(\mix1.data_reg[71] ));
 sky130_fd_sc_hd__dfrtp_1 _18178_ (.CLK(clknet_leaf_12_clk),
    .D(_01609_),
    .RESET_B(net621),
    .Q(\mix1.data_reg[72] ));
 sky130_fd_sc_hd__dfrtp_1 _18179_ (.CLK(clknet_leaf_12_clk),
    .D(_01610_),
    .RESET_B(net621),
    .Q(\mix1.data_reg[73] ));
 sky130_fd_sc_hd__dfrtp_1 _18180_ (.CLK(clknet_leaf_0_clk),
    .D(_01611_),
    .RESET_B(net619),
    .Q(\mix1.data_reg[74] ));
 sky130_fd_sc_hd__dfrtp_1 _18181_ (.CLK(clknet_leaf_1_clk),
    .D(_01612_),
    .RESET_B(net619),
    .Q(\mix1.data_reg[75] ));
 sky130_fd_sc_hd__dfrtp_1 _18182_ (.CLK(clknet_leaf_0_clk),
    .D(_01613_),
    .RESET_B(net619),
    .Q(\mix1.data_reg[76] ));
 sky130_fd_sc_hd__dfrtp_1 _18183_ (.CLK(clknet_leaf_1_clk),
    .D(_01614_),
    .RESET_B(net619),
    .Q(\mix1.data_reg[77] ));
 sky130_fd_sc_hd__dfrtp_1 _18184_ (.CLK(clknet_leaf_1_clk),
    .D(_01615_),
    .RESET_B(net619),
    .Q(\mix1.data_reg[78] ));
 sky130_fd_sc_hd__dfrtp_1 _18185_ (.CLK(clknet_leaf_14_clk),
    .D(_01616_),
    .RESET_B(net629),
    .Q(\mix1.data_reg[79] ));
 sky130_fd_sc_hd__dfrtp_1 _18186_ (.CLK(clknet_leaf_18_clk),
    .D(_01617_),
    .RESET_B(net638),
    .Q(\mix1.data_reg[80] ));
 sky130_fd_sc_hd__dfrtp_1 _18187_ (.CLK(clknet_leaf_18_clk),
    .D(_01618_),
    .RESET_B(net638),
    .Q(\mix1.data_reg[81] ));
 sky130_fd_sc_hd__dfrtp_1 _18188_ (.CLK(clknet_leaf_18_clk),
    .D(_01619_),
    .RESET_B(net638),
    .Q(\mix1.data_reg[82] ));
 sky130_fd_sc_hd__dfrtp_1 _18189_ (.CLK(clknet_leaf_24_clk),
    .D(_01620_),
    .RESET_B(net647),
    .Q(\mix1.data_reg[83] ));
 sky130_fd_sc_hd__dfrtp_1 _18190_ (.CLK(clknet_leaf_24_clk),
    .D(_01621_),
    .RESET_B(net644),
    .Q(\mix1.data_reg[84] ));
 sky130_fd_sc_hd__dfrtp_1 _18191_ (.CLK(clknet_leaf_24_clk),
    .D(_01622_),
    .RESET_B(net644),
    .Q(\mix1.data_reg[85] ));
 sky130_fd_sc_hd__dfrtp_1 _18192_ (.CLK(clknet_leaf_24_clk),
    .D(_01623_),
    .RESET_B(net647),
    .Q(\mix1.data_reg[86] ));
 sky130_fd_sc_hd__dfrtp_1 _18193_ (.CLK(clknet_leaf_24_clk),
    .D(_01624_),
    .RESET_B(net647),
    .Q(\mix1.data_reg[87] ));
 sky130_fd_sc_hd__dfrtp_1 _18194_ (.CLK(clknet_leaf_24_clk),
    .D(_01625_),
    .RESET_B(net647),
    .Q(\mix1.data_reg[88] ));
 sky130_fd_sc_hd__dfrtp_1 _18195_ (.CLK(clknet_leaf_25_clk),
    .D(_01626_),
    .RESET_B(net647),
    .Q(\mix1.data_reg[89] ));
 sky130_fd_sc_hd__dfrtp_1 _18196_ (.CLK(clknet_leaf_25_clk),
    .D(_01627_),
    .RESET_B(net648),
    .Q(\mix1.data_reg[90] ));
 sky130_fd_sc_hd__dfrtp_1 _18197_ (.CLK(clknet_leaf_25_clk),
    .D(_01628_),
    .RESET_B(net648),
    .Q(\mix1.data_reg[91] ));
 sky130_fd_sc_hd__dfrtp_1 _18198_ (.CLK(clknet_leaf_25_clk),
    .D(_01629_),
    .RESET_B(net648),
    .Q(\mix1.data_reg[92] ));
 sky130_fd_sc_hd__dfrtp_1 _18199_ (.CLK(clknet_leaf_10_clk),
    .D(_01630_),
    .RESET_B(net623),
    .Q(\mix1.data_reg[93] ));
 sky130_fd_sc_hd__dfrtp_1 _18200_ (.CLK(clknet_leaf_11_clk),
    .D(_01631_),
    .RESET_B(net622),
    .Q(\mix1.data_reg[94] ));
 sky130_fd_sc_hd__dfrtp_1 _18201_ (.CLK(clknet_leaf_12_clk),
    .D(_01632_),
    .RESET_B(net622),
    .Q(\mix1.data_reg[95] ));
 sky130_fd_sc_hd__dfrtp_1 _18202_ (.CLK(clknet_leaf_16_clk),
    .D(_01633_),
    .RESET_B(net637),
    .Q(\mix1.data_reg[32] ));
 sky130_fd_sc_hd__dfrtp_1 _18203_ (.CLK(clknet_leaf_15_clk),
    .D(_01634_),
    .RESET_B(net637),
    .Q(\mix1.data_reg[33] ));
 sky130_fd_sc_hd__dfrtp_1 _18204_ (.CLK(clknet_leaf_18_clk),
    .D(_01635_),
    .RESET_B(net636),
    .Q(\mix1.data_reg[34] ));
 sky130_fd_sc_hd__dfrtp_1 _18205_ (.CLK(clknet_leaf_18_clk),
    .D(_01636_),
    .RESET_B(net636),
    .Q(\mix1.data_reg[35] ));
 sky130_fd_sc_hd__dfrtp_1 _18206_ (.CLK(clknet_leaf_18_clk),
    .D(_01637_),
    .RESET_B(net636),
    .Q(\mix1.data_reg[36] ));
 sky130_fd_sc_hd__dfrtp_1 _18207_ (.CLK(clknet_leaf_15_clk),
    .D(_01638_),
    .RESET_B(net636),
    .Q(\mix1.data_reg[37] ));
 sky130_fd_sc_hd__dfrtp_1 _18208_ (.CLK(clknet_leaf_15_clk),
    .D(_01639_),
    .RESET_B(net629),
    .Q(\mix1.data_reg[38] ));
 sky130_fd_sc_hd__dfrtp_1 _18209_ (.CLK(clknet_leaf_15_clk),
    .D(_01640_),
    .RESET_B(net629),
    .Q(\mix1.data_reg[39] ));
 sky130_fd_sc_hd__dfrtp_1 _18210_ (.CLK(clknet_leaf_14_clk),
    .D(_01641_),
    .RESET_B(net629),
    .Q(\mix1.data_reg[40] ));
 sky130_fd_sc_hd__dfrtp_1 _18211_ (.CLK(clknet_leaf_12_clk),
    .D(_01642_),
    .RESET_B(net621),
    .Q(\mix1.data_reg[41] ));
 sky130_fd_sc_hd__dfrtp_1 _18212_ (.CLK(clknet_leaf_84_clk),
    .D(_01643_),
    .RESET_B(net581),
    .Q(\mix1.data_reg[42] ));
 sky130_fd_sc_hd__dfrtp_1 _18213_ (.CLK(clknet_leaf_84_clk),
    .D(_01644_),
    .RESET_B(net581),
    .Q(\mix1.data_reg[43] ));
 sky130_fd_sc_hd__dfrtp_1 _18214_ (.CLK(clknet_leaf_84_clk),
    .D(_01645_),
    .RESET_B(net581),
    .Q(\mix1.data_reg[44] ));
 sky130_fd_sc_hd__dfrtp_1 _18215_ (.CLK(clknet_leaf_84_clk),
    .D(_01646_),
    .RESET_B(net581),
    .Q(\mix1.data_reg[45] ));
 sky130_fd_sc_hd__dfrtp_1 _18216_ (.CLK(clknet_leaf_84_clk),
    .D(_01647_),
    .RESET_B(net581),
    .Q(\mix1.data_reg[46] ));
 sky130_fd_sc_hd__dfrtp_1 _18217_ (.CLK(clknet_leaf_0_clk),
    .D(_01648_),
    .RESET_B(net619),
    .Q(\mix1.data_reg[47] ));
 sky130_fd_sc_hd__dfrtp_1 _18218_ (.CLK(clknet_leaf_15_clk),
    .D(_01649_),
    .RESET_B(net629),
    .Q(\mix1.data_reg[48] ));
 sky130_fd_sc_hd__dfrtp_1 _18219_ (.CLK(clknet_leaf_19_clk),
    .D(_01650_),
    .RESET_B(net640),
    .Q(\mix1.data_reg[49] ));
 sky130_fd_sc_hd__dfrtp_1 _18220_ (.CLK(clknet_leaf_19_clk),
    .D(_01651_),
    .RESET_B(net640),
    .Q(\mix1.data_reg[50] ));
 sky130_fd_sc_hd__dfrtp_1 _18221_ (.CLK(clknet_leaf_36_clk),
    .D(_01652_),
    .RESET_B(net665),
    .Q(\mix1.data_reg[51] ));
 sky130_fd_sc_hd__dfrtp_1 _18222_ (.CLK(clknet_leaf_37_clk),
    .D(_01653_),
    .RESET_B(net666),
    .Q(\mix1.data_reg[52] ));
 sky130_fd_sc_hd__dfrtp_1 _18223_ (.CLK(clknet_leaf_37_clk),
    .D(_01654_),
    .RESET_B(net666),
    .Q(\mix1.data_reg[53] ));
 sky130_fd_sc_hd__dfrtp_1 _18224_ (.CLK(clknet_leaf_36_clk),
    .D(_01655_),
    .RESET_B(net665),
    .Q(\mix1.data_reg[54] ));
 sky130_fd_sc_hd__dfrtp_1 _18225_ (.CLK(clknet_leaf_36_clk),
    .D(_01656_),
    .RESET_B(net665),
    .Q(\mix1.data_reg[55] ));
 sky130_fd_sc_hd__dfrtp_1 _18226_ (.CLK(clknet_leaf_37_clk),
    .D(_01657_),
    .RESET_B(net666),
    .Q(\mix1.data_reg[56] ));
 sky130_fd_sc_hd__dfrtp_1 _18227_ (.CLK(clknet_leaf_36_clk),
    .D(_01658_),
    .RESET_B(net665),
    .Q(\mix1.data_reg[57] ));
 sky130_fd_sc_hd__dfrtp_1 _18228_ (.CLK(clknet_leaf_37_clk),
    .D(_01659_),
    .RESET_B(net666),
    .Q(\mix1.data_reg[58] ));
 sky130_fd_sc_hd__dfrtp_1 _18229_ (.CLK(clknet_leaf_38_clk),
    .D(_01660_),
    .RESET_B(net668),
    .Q(\mix1.data_reg[59] ));
 sky130_fd_sc_hd__dfrtp_1 _18230_ (.CLK(clknet_leaf_38_clk),
    .D(_01661_),
    .RESET_B(net668),
    .Q(\mix1.data_reg[60] ));
 sky130_fd_sc_hd__dfrtp_1 _18231_ (.CLK(clknet_leaf_36_clk),
    .D(_01662_),
    .RESET_B(net664),
    .Q(\mix1.data_reg[61] ));
 sky130_fd_sc_hd__dfrtp_2 _18232_ (.CLK(clknet_leaf_9_clk),
    .D(_01663_),
    .RESET_B(net631),
    .Q(\mix1.data_reg[62] ));
 sky130_fd_sc_hd__dfrtp_2 _18233_ (.CLK(clknet_leaf_11_clk),
    .D(_01664_),
    .RESET_B(net622),
    .Q(\mix1.data_reg[63] ));
 sky130_fd_sc_hd__dfrtp_2 _18234_ (.CLK(clknet_leaf_27_clk),
    .D(_01665_),
    .RESET_B(net641),
    .Q(\sub1.data_o[0] ));
 sky130_fd_sc_hd__dfrtp_2 _18235_ (.CLK(clknet_leaf_29_clk),
    .D(_01666_),
    .RESET_B(net635),
    .Q(\sub1.data_o[1] ));
 sky130_fd_sc_hd__dfrtp_2 _18236_ (.CLK(clknet_leaf_32_clk),
    .D(_01667_),
    .RESET_B(net653),
    .Q(\sub1.data_o[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18237_ (.CLK(clknet_leaf_26_clk),
    .D(_01668_),
    .RESET_B(net642),
    .Q(\sub1.data_o[3] ));
 sky130_fd_sc_hd__dfrtp_4 _18238_ (.CLK(clknet_leaf_32_clk),
    .D(_01669_),
    .RESET_B(net661),
    .Q(\sub1.data_o[4] ));
 sky130_fd_sc_hd__dfrtp_2 _18239_ (.CLK(clknet_leaf_32_clk),
    .D(_01670_),
    .RESET_B(net661),
    .Q(\sub1.data_o[5] ));
 sky130_fd_sc_hd__dfrtp_2 _18240_ (.CLK(clknet_leaf_39_clk),
    .D(_01671_),
    .RESET_B(net663),
    .Q(\sub1.data_o[6] ));
 sky130_fd_sc_hd__dfrtp_4 _18241_ (.CLK(clknet_leaf_35_clk),
    .D(_01672_),
    .RESET_B(net662),
    .Q(\sub1.data_o[7] ));
 sky130_fd_sc_hd__dfrtp_4 _18242_ (.CLK(clknet_leaf_10_clk),
    .D(_01673_),
    .RESET_B(net623),
    .Q(\sub1.data_o[8] ));
 sky130_fd_sc_hd__dfrtp_4 _18243_ (.CLK(clknet_leaf_2_clk),
    .D(_01674_),
    .RESET_B(net623),
    .Q(\sub1.data_o[9] ));
 sky130_fd_sc_hd__dfrtp_4 _18244_ (.CLK(clknet_leaf_10_clk),
    .D(_01675_),
    .RESET_B(net625),
    .Q(\sub1.data_o[10] ));
 sky130_fd_sc_hd__dfrtp_4 _18245_ (.CLK(clknet_leaf_2_clk),
    .D(_01676_),
    .RESET_B(net625),
    .Q(\sub1.data_o[11] ));
 sky130_fd_sc_hd__dfrtp_4 _18246_ (.CLK(clknet_leaf_10_clk),
    .D(_01677_),
    .RESET_B(net625),
    .Q(\sub1.data_o[12] ));
 sky130_fd_sc_hd__dfrtp_4 _18247_ (.CLK(clknet_leaf_2_clk),
    .D(_01678_),
    .RESET_B(net625),
    .Q(\sub1.data_o[13] ));
 sky130_fd_sc_hd__dfrtp_4 _18248_ (.CLK(clknet_leaf_10_clk),
    .D(_01679_),
    .RESET_B(net623),
    .Q(\sub1.data_o[14] ));
 sky130_fd_sc_hd__dfrtp_4 _18249_ (.CLK(clknet_leaf_1_clk),
    .D(_01680_),
    .RESET_B(net623),
    .Q(\sub1.data_o[15] ));
 sky130_fd_sc_hd__dfrtp_4 _18250_ (.CLK(clknet_leaf_21_clk),
    .D(_01681_),
    .RESET_B(net643),
    .Q(\sub1.data_o[16] ));
 sky130_fd_sc_hd__dfrtp_4 _18251_ (.CLK(clknet_leaf_23_clk),
    .D(_01682_),
    .RESET_B(net643),
    .Q(\sub1.data_o[17] ));
 sky130_fd_sc_hd__dfrtp_4 _18252_ (.CLK(clknet_leaf_21_clk),
    .D(_01683_),
    .RESET_B(net641),
    .Q(\sub1.data_o[18] ));
 sky130_fd_sc_hd__dfrtp_4 _18253_ (.CLK(clknet_leaf_22_clk),
    .D(_01684_),
    .RESET_B(net643),
    .Q(\sub1.data_o[19] ));
 sky130_fd_sc_hd__dfrtp_4 _18254_ (.CLK(clknet_leaf_21_clk),
    .D(_01685_),
    .RESET_B(net641),
    .Q(\sub1.data_o[20] ));
 sky130_fd_sc_hd__dfrtp_4 _18255_ (.CLK(clknet_leaf_22_clk),
    .D(_01686_),
    .RESET_B(net646),
    .Q(\sub1.data_o[21] ));
 sky130_fd_sc_hd__dfrtp_4 _18256_ (.CLK(clknet_leaf_22_clk),
    .D(_01687_),
    .RESET_B(net646),
    .Q(\sub1.data_o[22] ));
 sky130_fd_sc_hd__dfrtp_4 _18257_ (.CLK(clknet_leaf_21_clk),
    .D(_01688_),
    .RESET_B(net646),
    .Q(\sub1.data_o[23] ));
 sky130_fd_sc_hd__dfrtp_4 _18258_ (.CLK(clknet_leaf_47_clk),
    .D(_01689_),
    .RESET_B(net652),
    .Q(\sub1.data_o[24] ));
 sky130_fd_sc_hd__dfrtp_4 _18259_ (.CLK(clknet_leaf_43_clk),
    .D(_01690_),
    .RESET_B(net655),
    .Q(\sub1.data_o[25] ));
 sky130_fd_sc_hd__dfrtp_2 _18260_ (.CLK(clknet_leaf_51_clk),
    .D(_01691_),
    .RESET_B(net655),
    .Q(\sub1.data_o[26] ));
 sky130_fd_sc_hd__dfrtp_4 _18261_ (.CLK(clknet_leaf_42_clk),
    .D(_01692_),
    .RESET_B(net655),
    .Q(\sub1.data_o[27] ));
 sky130_fd_sc_hd__dfrtp_2 _18262_ (.CLK(clknet_leaf_43_clk),
    .D(_01693_),
    .RESET_B(net658),
    .Q(\sub1.data_o[28] ));
 sky130_fd_sc_hd__dfrtp_2 _18263_ (.CLK(clknet_leaf_52_clk),
    .D(_01694_),
    .RESET_B(net655),
    .Q(\sub1.data_o[29] ));
 sky130_fd_sc_hd__dfrtp_4 _18264_ (.CLK(clknet_leaf_52_clk),
    .D(_01695_),
    .RESET_B(net655),
    .Q(\sub1.data_o[30] ));
 sky130_fd_sc_hd__dfrtp_2 _18265_ (.CLK(clknet_leaf_43_clk),
    .D(_01696_),
    .RESET_B(net655),
    .Q(\sub1.data_o[31] ));
 sky130_fd_sc_hd__dfrtp_4 _18266_ (.CLK(clknet_leaf_34_clk),
    .D(_01697_),
    .RESET_B(net661),
    .Q(\sub1.data_o[32] ));
 sky130_fd_sc_hd__dfrtp_4 _18267_ (.CLK(clknet_leaf_32_clk),
    .D(_01698_),
    .RESET_B(net661),
    .Q(\sub1.data_o[33] ));
 sky130_fd_sc_hd__dfrtp_4 _18268_ (.CLK(clknet_leaf_33_clk),
    .D(_01699_),
    .RESET_B(net663),
    .Q(\sub1.data_o[34] ));
 sky130_fd_sc_hd__dfrtp_4 _18269_ (.CLK(clknet_leaf_34_clk),
    .D(_01700_),
    .RESET_B(net662),
    .Q(\sub1.data_o[35] ));
 sky130_fd_sc_hd__dfrtp_4 _18270_ (.CLK(clknet_leaf_33_clk),
    .D(_01701_),
    .RESET_B(net653),
    .Q(\sub1.data_o[36] ));
 sky130_fd_sc_hd__dfrtp_4 _18271_ (.CLK(clknet_leaf_32_clk),
    .D(_01702_),
    .RESET_B(net661),
    .Q(\sub1.data_o[37] ));
 sky130_fd_sc_hd__dfrtp_2 _18272_ (.CLK(clknet_leaf_34_clk),
    .D(_01703_),
    .RESET_B(net662),
    .Q(\sub1.data_o[38] ));
 sky130_fd_sc_hd__dfrtp_4 _18273_ (.CLK(clknet_leaf_34_clk),
    .D(_01704_),
    .RESET_B(net662),
    .Q(\sub1.data_o[39] ));
 sky130_fd_sc_hd__dfrtp_4 _18274_ (.CLK(clknet_leaf_3_clk),
    .D(_01705_),
    .RESET_B(net583),
    .Q(\sub1.data_o[40] ));
 sky130_fd_sc_hd__dfrtp_4 _18275_ (.CLK(clknet_leaf_3_clk),
    .D(_01706_),
    .RESET_B(net583),
    .Q(\sub1.data_o[41] ));
 sky130_fd_sc_hd__dfrtp_4 _18276_ (.CLK(clknet_leaf_2_clk),
    .D(_01707_),
    .RESET_B(net583),
    .Q(\sub1.data_o[42] ));
 sky130_fd_sc_hd__dfrtp_4 _18277_ (.CLK(clknet_leaf_3_clk),
    .D(_01708_),
    .RESET_B(net583),
    .Q(\sub1.data_o[43] ));
 sky130_fd_sc_hd__dfrtp_4 _18278_ (.CLK(clknet_leaf_5_clk),
    .D(_01709_),
    .RESET_B(net592),
    .Q(\sub1.data_o[44] ));
 sky130_fd_sc_hd__dfrtp_4 _18279_ (.CLK(clknet_leaf_5_clk),
    .D(_01710_),
    .RESET_B(net592),
    .Q(\sub1.data_o[45] ));
 sky130_fd_sc_hd__dfrtp_4 _18280_ (.CLK(clknet_leaf_1_clk),
    .D(_01711_),
    .RESET_B(net583),
    .Q(\sub1.data_o[46] ));
 sky130_fd_sc_hd__dfrtp_4 _18281_ (.CLK(clknet_leaf_3_clk),
    .D(_01712_),
    .RESET_B(net624),
    .Q(\sub1.data_o[47] ));
 sky130_fd_sc_hd__dfrtp_4 _18282_ (.CLK(clknet_leaf_22_clk),
    .D(_01713_),
    .RESET_B(net643),
    .Q(\sub1.data_o[48] ));
 sky130_fd_sc_hd__dfrtp_4 _18283_ (.CLK(clknet_leaf_22_clk),
    .D(_01714_),
    .RESET_B(net643),
    .Q(\sub1.data_o[49] ));
 sky130_fd_sc_hd__dfrtp_4 _18284_ (.CLK(clknet_leaf_21_clk),
    .D(_01715_),
    .RESET_B(net641),
    .Q(\sub1.data_o[50] ));
 sky130_fd_sc_hd__dfrtp_4 _18285_ (.CLK(clknet_leaf_26_clk),
    .D(_01716_),
    .RESET_B(net649),
    .Q(\sub1.data_o[51] ));
 sky130_fd_sc_hd__dfrtp_4 _18286_ (.CLK(clknet_leaf_26_clk),
    .D(_01717_),
    .RESET_B(net642),
    .Q(\sub1.data_o[52] ));
 sky130_fd_sc_hd__dfrtp_4 _18287_ (.CLK(clknet_leaf_26_clk),
    .D(_01718_),
    .RESET_B(net649),
    .Q(\sub1.data_o[53] ));
 sky130_fd_sc_hd__dfrtp_4 _18288_ (.CLK(clknet_leaf_26_clk),
    .D(_01719_),
    .RESET_B(net649),
    .Q(\sub1.data_o[54] ));
 sky130_fd_sc_hd__dfrtp_4 _18289_ (.CLK(clknet_leaf_26_clk),
    .D(_01720_),
    .RESET_B(net649),
    .Q(\sub1.data_o[55] ));
 sky130_fd_sc_hd__dfrtp_1 _18290_ (.CLK(clknet_leaf_46_clk),
    .D(_01721_),
    .RESET_B(net652),
    .Q(\sub1.data_o[56] ));
 sky130_fd_sc_hd__dfrtp_1 _18291_ (.CLK(clknet_leaf_71_clk),
    .D(_01722_),
    .RESET_B(net652),
    .Q(\sub1.data_o[57] ));
 sky130_fd_sc_hd__dfrtp_1 _18292_ (.CLK(clknet_leaf_46_clk),
    .D(_01723_),
    .RESET_B(net651),
    .Q(\sub1.data_o[58] ));
 sky130_fd_sc_hd__dfrtp_2 _18293_ (.CLK(clknet_leaf_47_clk),
    .D(_01724_),
    .RESET_B(net652),
    .Q(\sub1.data_o[59] ));
 sky130_fd_sc_hd__dfrtp_1 _18294_ (.CLK(clknet_leaf_45_clk),
    .D(_01725_),
    .RESET_B(net652),
    .Q(\sub1.data_o[60] ));
 sky130_fd_sc_hd__dfrtp_2 _18295_ (.CLK(clknet_leaf_47_clk),
    .D(_01726_),
    .RESET_B(net651),
    .Q(\sub1.data_o[61] ));
 sky130_fd_sc_hd__dfrtp_2 _18296_ (.CLK(clknet_leaf_51_clk),
    .D(_01727_),
    .RESET_B(net651),
    .Q(\sub1.data_o[62] ));
 sky130_fd_sc_hd__dfrtp_1 _18297_ (.CLK(clknet_leaf_46_clk),
    .D(_01728_),
    .RESET_B(net652),
    .Q(\sub1.data_o[63] ));
 sky130_fd_sc_hd__dfrtp_4 _18298_ (.CLK(clknet_leaf_27_clk),
    .D(_01729_),
    .RESET_B(net642),
    .Q(\sub1.data_o[64] ));
 sky130_fd_sc_hd__dfrtp_4 _18299_ (.CLK(clknet_leaf_29_clk),
    .D(_01730_),
    .RESET_B(net642),
    .Q(\sub1.data_o[65] ));
 sky130_fd_sc_hd__dfrtp_4 _18300_ (.CLK(clknet_leaf_30_clk),
    .D(_01731_),
    .RESET_B(net642),
    .Q(\sub1.data_o[66] ));
 sky130_fd_sc_hd__dfrtp_4 _18301_ (.CLK(clknet_leaf_27_clk),
    .D(_01732_),
    .RESET_B(net642),
    .Q(\sub1.data_o[67] ));
 sky130_fd_sc_hd__dfrtp_4 _18302_ (.CLK(clknet_leaf_32_clk),
    .D(_01733_),
    .RESET_B(net661),
    .Q(\sub1.data_o[68] ));
 sky130_fd_sc_hd__dfrtp_4 _18303_ (.CLK(clknet_leaf_34_clk),
    .D(_01734_),
    .RESET_B(net661),
    .Q(\sub1.data_o[69] ));
 sky130_fd_sc_hd__dfrtp_4 _18304_ (.CLK(clknet_leaf_34_clk),
    .D(_01735_),
    .RESET_B(net661),
    .Q(\sub1.data_o[70] ));
 sky130_fd_sc_hd__dfrtp_4 _18305_ (.CLK(clknet_leaf_34_clk),
    .D(_01736_),
    .RESET_B(net662),
    .Q(\sub1.data_o[71] ));
 sky130_fd_sc_hd__dfrtp_4 _18306_ (.CLK(clknet_leaf_1_clk),
    .D(_01737_),
    .RESET_B(net624),
    .Q(\sub1.data_o[72] ));
 sky130_fd_sc_hd__dfrtp_4 _18307_ (.CLK(clknet_leaf_1_clk),
    .D(_01738_),
    .RESET_B(net624),
    .Q(\sub1.data_o[73] ));
 sky130_fd_sc_hd__dfrtp_2 _18308_ (.CLK(clknet_leaf_2_clk),
    .D(_01739_),
    .RESET_B(net624),
    .Q(\sub1.data_o[74] ));
 sky130_fd_sc_hd__dfrtp_2 _18309_ (.CLK(clknet_leaf_2_clk),
    .D(_01740_),
    .RESET_B(net624),
    .Q(\sub1.data_o[75] ));
 sky130_fd_sc_hd__dfrtp_2 _18310_ (.CLK(clknet_leaf_2_clk),
    .D(_01741_),
    .RESET_B(net624),
    .Q(\sub1.data_o[76] ));
 sky130_fd_sc_hd__dfrtp_2 _18311_ (.CLK(clknet_leaf_5_clk),
    .D(_01742_),
    .RESET_B(net624),
    .Q(\sub1.data_o[77] ));
 sky130_fd_sc_hd__dfrtp_4 _18312_ (.CLK(clknet_leaf_1_clk),
    .D(_01743_),
    .RESET_B(net624),
    .Q(\sub1.data_o[78] ));
 sky130_fd_sc_hd__dfrtp_4 _18313_ (.CLK(clknet_leaf_1_clk),
    .D(_01744_),
    .RESET_B(net624),
    .Q(\sub1.data_o[79] ));
 sky130_fd_sc_hd__dfrtp_4 _18314_ (.CLK(clknet_leaf_21_clk),
    .D(\sub1.next_ready_o ),
    .RESET_B(net643),
    .Q(\sub1.ready_o ));
 sky130_fd_sc_hd__dfrtp_4 _18315_ (.CLK(clknet_leaf_9_clk),
    .D(_01745_),
    .RESET_B(net633),
    .Q(\mix1.data_o[0] ));
 sky130_fd_sc_hd__dfrtp_4 _18316_ (.CLK(clknet_leaf_17_clk),
    .D(_01746_),
    .RESET_B(net633),
    .Q(\mix1.data_o[1] ));
 sky130_fd_sc_hd__dfrtp_4 _18317_ (.CLK(clknet_leaf_9_clk),
    .D(_01747_),
    .RESET_B(net633),
    .Q(\mix1.data_o[2] ));
 sky130_fd_sc_hd__dfrtp_4 _18318_ (.CLK(clknet_leaf_8_clk),
    .D(_01748_),
    .RESET_B(net632),
    .Q(\mix1.data_o[3] ));
 sky130_fd_sc_hd__dfrtp_4 _18319_ (.CLK(clknet_leaf_8_clk),
    .D(_01749_),
    .RESET_B(net633),
    .Q(\mix1.data_o[4] ));
 sky130_fd_sc_hd__dfrtp_4 _18320_ (.CLK(clknet_leaf_9_clk),
    .D(_01750_),
    .RESET_B(net633),
    .Q(\mix1.data_o[5] ));
 sky130_fd_sc_hd__dfrtp_4 _18321_ (.CLK(clknet_leaf_8_clk),
    .D(_01751_),
    .RESET_B(net634),
    .Q(\mix1.data_o[6] ));
 sky130_fd_sc_hd__dfrtp_4 _18322_ (.CLK(clknet_leaf_9_clk),
    .D(_01752_),
    .RESET_B(net631),
    .Q(\mix1.data_o[7] ));
 sky130_fd_sc_hd__dfrtp_4 _18323_ (.CLK(clknet_leaf_9_clk),
    .D(_01753_),
    .RESET_B(net631),
    .Q(\mix1.data_o[8] ));
 sky130_fd_sc_hd__dfrtp_4 _18324_ (.CLK(clknet_leaf_9_clk),
    .D(_01754_),
    .RESET_B(net631),
    .Q(\mix1.data_o[9] ));
 sky130_fd_sc_hd__dfrtp_4 _18325_ (.CLK(clknet_leaf_11_clk),
    .D(_01755_),
    .RESET_B(net628),
    .Q(\mix1.data_o[10] ));
 sky130_fd_sc_hd__dfrtp_4 _18326_ (.CLK(clknet_leaf_11_clk),
    .D(_01756_),
    .RESET_B(net631),
    .Q(\mix1.data_o[11] ));
 sky130_fd_sc_hd__dfrtp_4 _18327_ (.CLK(clknet_leaf_11_clk),
    .D(_01757_),
    .RESET_B(net631),
    .Q(\mix1.data_o[12] ));
 sky130_fd_sc_hd__dfrtp_4 _18328_ (.CLK(clknet_leaf_9_clk),
    .D(_01758_),
    .RESET_B(net631),
    .Q(\mix1.data_o[13] ));
 sky130_fd_sc_hd__dfrtp_4 _18329_ (.CLK(clknet_leaf_11_clk),
    .D(_01759_),
    .RESET_B(net628),
    .Q(\mix1.data_o[14] ));
 sky130_fd_sc_hd__dfrtp_4 _18330_ (.CLK(clknet_leaf_11_clk),
    .D(_01760_),
    .RESET_B(net628),
    .Q(\mix1.data_o[15] ));
 sky130_fd_sc_hd__dfrtp_4 _18331_ (.CLK(clknet_leaf_16_clk),
    .D(_01761_),
    .RESET_B(net630),
    .Q(\mix1.data_o[16] ));
 sky130_fd_sc_hd__dfrtp_4 _18332_ (.CLK(clknet_leaf_16_clk),
    .D(_01762_),
    .RESET_B(net637),
    .Q(\mix1.data_o[17] ));
 sky130_fd_sc_hd__dfrtp_4 _18333_ (.CLK(clknet_leaf_16_clk),
    .D(_01763_),
    .RESET_B(net630),
    .Q(\mix1.data_o[18] ));
 sky130_fd_sc_hd__dfrtp_4 _18334_ (.CLK(clknet_leaf_35_clk),
    .D(_01764_),
    .RESET_B(net664),
    .Q(\mix1.data_o[19] ));
 sky130_fd_sc_hd__dfrtp_4 _18335_ (.CLK(clknet_leaf_37_clk),
    .D(_01765_),
    .RESET_B(net664),
    .Q(\mix1.data_o[20] ));
 sky130_fd_sc_hd__dfrtp_4 _18336_ (.CLK(clknet_leaf_37_clk),
    .D(_01766_),
    .RESET_B(net664),
    .Q(\mix1.data_o[21] ));
 sky130_fd_sc_hd__dfrtp_4 _18337_ (.CLK(clknet_leaf_35_clk),
    .D(_01767_),
    .RESET_B(net664),
    .Q(\mix1.data_o[22] ));
 sky130_fd_sc_hd__dfrtp_4 _18338_ (.CLK(clknet_leaf_35_clk),
    .D(_01768_),
    .RESET_B(net664),
    .Q(\mix1.data_o[23] ));
 sky130_fd_sc_hd__dfrtp_4 _18339_ (.CLK(clknet_leaf_35_clk),
    .D(_01769_),
    .RESET_B(net664),
    .Q(\mix1.data_o[24] ));
 sky130_fd_sc_hd__dfrtp_4 _18340_ (.CLK(clknet_leaf_35_clk),
    .D(_01770_),
    .RESET_B(net664),
    .Q(\mix1.data_o[25] ));
 sky130_fd_sc_hd__dfrtp_4 _18341_ (.CLK(clknet_leaf_37_clk),
    .D(_01771_),
    .RESET_B(net668),
    .Q(\mix1.data_o[26] ));
 sky130_fd_sc_hd__dfrtp_4 _18342_ (.CLK(clknet_leaf_38_clk),
    .D(_01772_),
    .RESET_B(net668),
    .Q(\mix1.data_o[27] ));
 sky130_fd_sc_hd__dfrtp_4 _18343_ (.CLK(clknet_leaf_38_clk),
    .D(_01773_),
    .RESET_B(net668),
    .Q(\mix1.data_o[28] ));
 sky130_fd_sc_hd__dfrtp_4 _18344_ (.CLK(clknet_leaf_11_clk),
    .D(_01774_),
    .RESET_B(net623),
    .Q(\mix1.data_o[29] ));
 sky130_fd_sc_hd__dfrtp_4 _18345_ (.CLK(clknet_leaf_11_clk),
    .D(_01775_),
    .RESET_B(net631),
    .Q(\mix1.data_o[30] ));
 sky130_fd_sc_hd__dfrtp_4 _18346_ (.CLK(clknet_leaf_11_clk),
    .D(_01776_),
    .RESET_B(net623),
    .Q(\mix1.data_o[31] ));
 sky130_fd_sc_hd__dfrtp_4 _18347_ (.CLK(clknet_leaf_18_clk),
    .D(_01777_),
    .RESET_B(net637),
    .Q(\mix1.data_o[32] ));
 sky130_fd_sc_hd__dfrtp_4 _18348_ (.CLK(clknet_leaf_16_clk),
    .D(_01778_),
    .RESET_B(net637),
    .Q(\mix1.data_o[33] ));
 sky130_fd_sc_hd__dfrtp_4 _18349_ (.CLK(clknet_leaf_15_clk),
    .D(_01779_),
    .RESET_B(net636),
    .Q(\mix1.data_o[34] ));
 sky130_fd_sc_hd__dfrtp_4 _18350_ (.CLK(clknet_leaf_18_clk),
    .D(_01780_),
    .RESET_B(net637),
    .Q(\mix1.data_o[35] ));
 sky130_fd_sc_hd__dfrtp_4 _18351_ (.CLK(clknet_leaf_15_clk),
    .D(_01781_),
    .RESET_B(net636),
    .Q(\mix1.data_o[36] ));
 sky130_fd_sc_hd__dfrtp_4 _18352_ (.CLK(clknet_leaf_15_clk),
    .D(_01782_),
    .RESET_B(net636),
    .Q(\mix1.data_o[37] ));
 sky130_fd_sc_hd__dfrtp_4 _18353_ (.CLK(clknet_leaf_15_clk),
    .D(_01783_),
    .RESET_B(net629),
    .Q(\mix1.data_o[38] ));
 sky130_fd_sc_hd__dfrtp_4 _18354_ (.CLK(clknet_leaf_15_clk),
    .D(_01784_),
    .RESET_B(net629),
    .Q(\mix1.data_o[39] ));
 sky130_fd_sc_hd__dfrtp_4 _18355_ (.CLK(clknet_leaf_14_clk),
    .D(_01785_),
    .RESET_B(net627),
    .Q(\mix1.data_o[40] ));
 sky130_fd_sc_hd__dfrtp_4 _18356_ (.CLK(clknet_leaf_12_clk),
    .D(_01786_),
    .RESET_B(net621),
    .Q(\mix1.data_o[41] ));
 sky130_fd_sc_hd__dfrtp_4 _18357_ (.CLK(clknet_leaf_84_clk),
    .D(_01787_),
    .RESET_B(net581),
    .Q(\mix1.data_o[42] ));
 sky130_fd_sc_hd__dfrtp_4 _18358_ (.CLK(clknet_leaf_83_clk),
    .D(_01788_),
    .RESET_B(net581),
    .Q(\mix1.data_o[43] ));
 sky130_fd_sc_hd__dfrtp_4 _18359_ (.CLK(clknet_leaf_84_clk),
    .D(_01789_),
    .RESET_B(net581),
    .Q(\mix1.data_o[44] ));
 sky130_fd_sc_hd__dfrtp_4 _18360_ (.CLK(clknet_leaf_1_clk),
    .D(_01790_),
    .RESET_B(net581),
    .Q(\mix1.data_o[45] ));
 sky130_fd_sc_hd__dfrtp_4 _18361_ (.CLK(clknet_leaf_84_clk),
    .D(_01791_),
    .RESET_B(net582),
    .Q(\mix1.data_o[46] ));
 sky130_fd_sc_hd__dfrtp_4 _18362_ (.CLK(clknet_leaf_0_clk),
    .D(_01792_),
    .RESET_B(net619),
    .Q(\mix1.data_o[47] ));
 sky130_fd_sc_hd__dfrtp_4 _18363_ (.CLK(clknet_leaf_15_clk),
    .D(_01793_),
    .RESET_B(net630),
    .Q(\mix1.data_o[48] ));
 sky130_fd_sc_hd__dfrtp_2 _18364_ (.CLK(clknet_leaf_35_clk),
    .D(_01794_),
    .RESET_B(net667),
    .Q(\mix1.data_o[49] ));
 sky130_fd_sc_hd__dfrtp_4 _18365_ (.CLK(clknet_leaf_35_clk),
    .D(_01795_),
    .RESET_B(net664),
    .Q(\mix1.data_o[50] ));
 sky130_fd_sc_hd__dfrtp_4 _18366_ (.CLK(clknet_leaf_36_clk),
    .D(_01796_),
    .RESET_B(net665),
    .Q(\mix1.data_o[51] ));
 sky130_fd_sc_hd__dfrtp_2 _18367_ (.CLK(clknet_leaf_37_clk),
    .D(_01797_),
    .RESET_B(net667),
    .Q(\mix1.data_o[52] ));
 sky130_fd_sc_hd__dfrtp_2 _18368_ (.CLK(clknet_leaf_37_clk),
    .D(_01798_),
    .RESET_B(net666),
    .Q(\mix1.data_o[53] ));
 sky130_fd_sc_hd__dfrtp_4 _18369_ (.CLK(clknet_leaf_37_clk),
    .D(_01799_),
    .RESET_B(net666),
    .Q(\mix1.data_o[54] ));
 sky130_fd_sc_hd__dfrtp_1 _18370_ (.CLK(clknet_leaf_36_clk),
    .D(_01800_),
    .RESET_B(net665),
    .Q(\mix1.data_o[55] ));
 sky130_fd_sc_hd__dfrtp_4 _18371_ (.CLK(clknet_leaf_37_clk),
    .D(_01801_),
    .RESET_B(net667),
    .Q(\mix1.data_o[56] ));
 sky130_fd_sc_hd__dfrtp_4 _18372_ (.CLK(clknet_leaf_37_clk),
    .D(_01802_),
    .RESET_B(net667),
    .Q(\mix1.data_o[57] ));
 sky130_fd_sc_hd__dfrtp_4 _18373_ (.CLK(clknet_leaf_37_clk),
    .D(_01803_),
    .RESET_B(net668),
    .Q(\mix1.data_o[58] ));
 sky130_fd_sc_hd__dfrtp_4 _18374_ (.CLK(clknet_leaf_38_clk),
    .D(_01804_),
    .RESET_B(net668),
    .Q(\mix1.data_o[59] ));
 sky130_fd_sc_hd__dfrtp_4 _18375_ (.CLK(clknet_leaf_38_clk),
    .D(_01805_),
    .RESET_B(net669),
    .Q(\mix1.data_o[60] ));
 sky130_fd_sc_hd__dfrtp_4 _18376_ (.CLK(clknet_leaf_35_clk),
    .D(_01806_),
    .RESET_B(net664),
    .Q(\mix1.data_o[61] ));
 sky130_fd_sc_hd__dfrtp_1 _18377_ (.CLK(clknet_3_6__leaf_clk),
    .D(_01807_),
    .RESET_B(net653),
    .Q(\mix1.data_o[62] ));
 sky130_fd_sc_hd__dfrtp_1 _18378_ (.CLK(clknet_leaf_46_clk),
    .D(_01808_),
    .RESET_B(net652),
    .Q(\mix1.data_o[63] ));
 sky130_fd_sc_hd__dfrtp_2 _18379_ (.CLK(clknet_3_3__leaf_clk),
    .D(_01809_),
    .RESET_B(net635),
    .Q(\mix1.data_o[64] ));
 sky130_fd_sc_hd__dfrtp_4 _18380_ (.CLK(clknet_leaf_30_clk),
    .D(_01810_),
    .RESET_B(net635),
    .Q(\mix1.data_o[65] ));
 sky130_fd_sc_hd__dfrtp_4 _18381_ (.CLK(clknet_leaf_36_clk),
    .D(_01811_),
    .RESET_B(net665),
    .Q(\mix1.data_o[66] ));
 sky130_fd_sc_hd__dfrtp_4 _18382_ (.CLK(clknet_leaf_26_clk),
    .D(_01812_),
    .RESET_B(net648),
    .Q(\mix1.data_o[67] ));
 sky130_fd_sc_hd__dfrtp_4 _18383_ (.CLK(clknet_leaf_25_clk),
    .D(_01813_),
    .RESET_B(net648),
    .Q(\mix1.data_o[68] ));
 sky130_fd_sc_hd__dfrtp_4 _18384_ (.CLK(clknet_leaf_12_clk),
    .D(_01814_),
    .RESET_B(net621),
    .Q(\mix1.data_o[69] ));
 sky130_fd_sc_hd__dfrtp_4 _18385_ (.CLK(clknet_leaf_12_clk),
    .D(_01815_),
    .RESET_B(net621),
    .Q(\mix1.data_o[70] ));
 sky130_fd_sc_hd__dfrtp_4 _18386_ (.CLK(clknet_leaf_0_clk),
    .D(_01816_),
    .RESET_B(net621),
    .Q(\mix1.data_o[71] ));
 sky130_fd_sc_hd__dfrtp_4 _18387_ (.CLK(clknet_leaf_12_clk),
    .D(_01817_),
    .RESET_B(net621),
    .Q(\mix1.data_o[72] ));
 sky130_fd_sc_hd__dfrtp_4 _18388_ (.CLK(clknet_leaf_12_clk),
    .D(_01818_),
    .RESET_B(net622),
    .Q(\mix1.data_o[73] ));
 sky130_fd_sc_hd__dfrtp_2 _18389_ (.CLK(clknet_leaf_0_clk),
    .D(_01819_),
    .RESET_B(net619),
    .Q(\mix1.data_o[74] ));
 sky130_fd_sc_hd__dfrtp_4 _18390_ (.CLK(clknet_leaf_84_clk),
    .D(_01820_),
    .RESET_B(net619),
    .Q(\mix1.data_o[75] ));
 sky130_fd_sc_hd__dfrtp_2 _18391_ (.CLK(clknet_leaf_0_clk),
    .D(_01821_),
    .RESET_B(net620),
    .Q(\mix1.data_o[76] ));
 sky130_fd_sc_hd__dfrtp_4 _18392_ (.CLK(clknet_leaf_1_clk),
    .D(_01822_),
    .RESET_B(net620),
    .Q(\mix1.data_o[77] ));
 sky130_fd_sc_hd__dfrtp_4 _18393_ (.CLK(clknet_leaf_1_clk),
    .D(_01823_),
    .RESET_B(net620),
    .Q(\mix1.data_o[78] ));
 sky130_fd_sc_hd__dfrtp_4 _18394_ (.CLK(clknet_leaf_14_clk),
    .D(_01824_),
    .RESET_B(net629),
    .Q(\mix1.data_o[79] ));
 sky130_fd_sc_hd__dfrtp_4 _18395_ (.CLK(clknet_leaf_18_clk),
    .D(_01825_),
    .RESET_B(net638),
    .Q(\mix1.data_o[80] ));
 sky130_fd_sc_hd__dfrtp_4 _18396_ (.CLK(clknet_leaf_19_clk),
    .D(_01826_),
    .RESET_B(net640),
    .Q(\mix1.data_o[81] ));
 sky130_fd_sc_hd__dfrtp_4 _18397_ (.CLK(clknet_leaf_18_clk),
    .D(_01827_),
    .RESET_B(net638),
    .Q(\mix1.data_o[82] ));
 sky130_fd_sc_hd__dfrtp_2 _18398_ (.CLK(clknet_leaf_24_clk),
    .D(_01828_),
    .RESET_B(net647),
    .Q(\mix1.data_o[83] ));
 sky130_fd_sc_hd__dfrtp_2 _18399_ (.CLK(clknet_leaf_24_clk),
    .D(_01829_),
    .RESET_B(net646),
    .Q(\mix1.data_o[84] ));
 sky130_fd_sc_hd__dfrtp_2 _18400_ (.CLK(clknet_leaf_24_clk),
    .D(_01830_),
    .RESET_B(net647),
    .Q(\mix1.data_o[85] ));
 sky130_fd_sc_hd__dfrtp_2 _18401_ (.CLK(clknet_leaf_24_clk),
    .D(_01831_),
    .RESET_B(net647),
    .Q(\mix1.data_o[86] ));
 sky130_fd_sc_hd__dfrtp_1 _18402_ (.CLK(clknet_leaf_25_clk),
    .D(_01832_),
    .RESET_B(net647),
    .Q(\mix1.data_o[87] ));
 sky130_fd_sc_hd__dfrtp_4 _18403_ (.CLK(clknet_leaf_25_clk),
    .D(_01833_),
    .RESET_B(net647),
    .Q(\mix1.data_o[88] ));
 sky130_fd_sc_hd__dfrtp_4 _18404_ (.CLK(clknet_leaf_25_clk),
    .D(_01834_),
    .RESET_B(net648),
    .Q(\mix1.data_o[89] ));
 sky130_fd_sc_hd__dfrtp_4 _18405_ (.CLK(clknet_leaf_25_clk),
    .D(_01835_),
    .RESET_B(net648),
    .Q(\mix1.data_o[90] ));
 sky130_fd_sc_hd__dfrtp_4 _18406_ (.CLK(clknet_leaf_25_clk),
    .D(_01836_),
    .RESET_B(net648),
    .Q(\mix1.data_o[91] ));
 sky130_fd_sc_hd__dfrtp_4 _18407_ (.CLK(clknet_leaf_25_clk),
    .D(_01837_),
    .RESET_B(net650),
    .Q(\mix1.data_o[92] ));
 sky130_fd_sc_hd__dfrtp_4 _18408_ (.CLK(clknet_leaf_10_clk),
    .D(_01838_),
    .RESET_B(net623),
    .Q(\mix1.data_o[93] ));
 sky130_fd_sc_hd__dfrtp_4 _18409_ (.CLK(clknet_leaf_10_clk),
    .D(_01839_),
    .RESET_B(net623),
    .Q(\mix1.data_o[94] ));
 sky130_fd_sc_hd__dfrtp_4 _18410_ (.CLK(clknet_leaf_0_clk),
    .D(_01840_),
    .RESET_B(net622),
    .Q(\mix1.data_o[95] ));
 sky130_fd_sc_hd__dfrtp_4 _18411_ (.CLK(clknet_leaf_13_clk),
    .D(_01841_),
    .RESET_B(net628),
    .Q(\mix1.data_o[96] ));
 sky130_fd_sc_hd__dfrtp_2 _18412_ (.CLK(clknet_leaf_14_clk),
    .D(_01842_),
    .RESET_B(net630),
    .Q(\mix1.data_o[97] ));
 sky130_fd_sc_hd__dfrtp_4 _18413_ (.CLK(clknet_leaf_16_clk),
    .D(_01843_),
    .RESET_B(net630),
    .Q(\mix1.data_o[98] ));
 sky130_fd_sc_hd__dfrtp_2 _18414_ (.CLK(clknet_leaf_13_clk),
    .D(_01844_),
    .RESET_B(net628),
    .Q(\mix1.data_o[99] ));
 sky130_fd_sc_hd__dfrtp_4 _18415_ (.CLK(clknet_leaf_13_clk),
    .D(_01845_),
    .RESET_B(net627),
    .Q(\mix1.data_o[100] ));
 sky130_fd_sc_hd__dfrtp_2 _18416_ (.CLK(clknet_leaf_13_clk),
    .D(_01846_),
    .RESET_B(net627),
    .Q(\mix1.data_o[101] ));
 sky130_fd_sc_hd__dfrtp_2 _18417_ (.CLK(clknet_leaf_11_clk),
    .D(_01847_),
    .RESET_B(net628),
    .Q(\mix1.data_o[102] ));
 sky130_fd_sc_hd__dfrtp_4 _18418_ (.CLK(clknet_leaf_13_clk),
    .D(_01848_),
    .RESET_B(net627),
    .Q(\mix1.data_o[103] ));
 sky130_fd_sc_hd__dfrtp_4 _18419_ (.CLK(clknet_leaf_12_clk),
    .D(_01849_),
    .RESET_B(net621),
    .Q(\mix1.data_o[104] ));
 sky130_fd_sc_hd__dfrtp_4 _18420_ (.CLK(clknet_leaf_11_clk),
    .D(_01850_),
    .RESET_B(net622),
    .Q(\mix1.data_o[105] ));
 sky130_fd_sc_hd__dfrtp_2 _18421_ (.CLK(clknet_leaf_84_clk),
    .D(_01851_),
    .RESET_B(net582),
    .Q(\mix1.data_o[106] ));
 sky130_fd_sc_hd__dfrtp_2 _18422_ (.CLK(clknet_leaf_83_clk),
    .D(_01852_),
    .RESET_B(net582),
    .Q(\mix1.data_o[107] ));
 sky130_fd_sc_hd__dfrtp_2 _18423_ (.CLK(clknet_leaf_83_clk),
    .D(_01853_),
    .RESET_B(net582),
    .Q(\mix1.data_o[108] ));
 sky130_fd_sc_hd__dfrtp_2 _18424_ (.CLK(clknet_leaf_83_clk),
    .D(_01854_),
    .RESET_B(net584),
    .Q(\mix1.data_o[109] ));
 sky130_fd_sc_hd__dfrtp_2 _18425_ (.CLK(clknet_leaf_3_clk),
    .D(_01855_),
    .RESET_B(net583),
    .Q(\mix1.data_o[110] ));
 sky130_fd_sc_hd__dfrtp_2 _18426_ (.CLK(clknet_leaf_0_clk),
    .D(_01856_),
    .RESET_B(net620),
    .Q(\mix1.data_o[111] ));
 sky130_fd_sc_hd__dfrtp_4 _18427_ (.CLK(clknet_leaf_15_clk),
    .D(_01857_),
    .RESET_B(net636),
    .Q(\mix1.data_o[112] ));
 sky130_fd_sc_hd__dfrtp_4 _18428_ (.CLK(clknet_leaf_15_clk),
    .D(_01858_),
    .RESET_B(net637),
    .Q(\mix1.data_o[113] ));
 sky130_fd_sc_hd__dfrtp_2 _18429_ (.CLK(clknet_leaf_16_clk),
    .D(_01859_),
    .RESET_B(net630),
    .Q(\mix1.data_o[114] ));
 sky130_fd_sc_hd__dfrtp_2 _18430_ (.CLK(clknet_leaf_23_clk),
    .D(_01860_),
    .RESET_B(net644),
    .Q(\mix1.data_o[115] ));
 sky130_fd_sc_hd__dfrtp_2 _18431_ (.CLK(clknet_leaf_24_clk),
    .D(_01861_),
    .RESET_B(net644),
    .Q(\mix1.data_o[116] ));
 sky130_fd_sc_hd__dfrtp_2 _18432_ (.CLK(clknet_leaf_24_clk),
    .D(_01862_),
    .RESET_B(net644),
    .Q(\mix1.data_o[117] ));
 sky130_fd_sc_hd__dfrtp_2 _18433_ (.CLK(clknet_leaf_23_clk),
    .D(_01863_),
    .RESET_B(net644),
    .Q(\mix1.data_o[118] ));
 sky130_fd_sc_hd__dfrtp_2 _18434_ (.CLK(clknet_leaf_24_clk),
    .D(_01864_),
    .RESET_B(net644),
    .Q(\mix1.data_o[119] ));
 sky130_fd_sc_hd__dfrtp_4 _18435_ (.CLK(clknet_leaf_23_clk),
    .D(_01865_),
    .RESET_B(net645),
    .Q(\mix1.data_o[120] ));
 sky130_fd_sc_hd__dfrtp_4 _18436_ (.CLK(clknet_leaf_25_clk),
    .D(_01866_),
    .RESET_B(net650),
    .Q(\mix1.data_o[121] ));
 sky130_fd_sc_hd__dfrtp_4 _18437_ (.CLK(clknet_leaf_24_clk),
    .D(_01867_),
    .RESET_B(net645),
    .Q(\mix1.data_o[122] ));
 sky130_fd_sc_hd__dfrtp_4 _18438_ (.CLK(clknet_leaf_36_clk),
    .D(_01868_),
    .RESET_B(net665),
    .Q(\mix1.data_o[123] ));
 sky130_fd_sc_hd__dfrtp_4 _18439_ (.CLK(clknet_leaf_36_clk),
    .D(_01869_),
    .RESET_B(net666),
    .Q(\mix1.data_o[124] ));
 sky130_fd_sc_hd__dfrtp_4 _18440_ (.CLK(clknet_leaf_35_clk),
    .D(_01870_),
    .RESET_B(net665),
    .Q(\mix1.data_o[125] ));
 sky130_fd_sc_hd__dfrtp_4 _18441_ (.CLK(clknet_leaf_1_clk),
    .D(_01871_),
    .RESET_B(net624),
    .Q(\mix1.data_o[126] ));
 sky130_fd_sc_hd__dfrtp_4 _18442_ (.CLK(clknet_leaf_1_clk),
    .D(_01872_),
    .RESET_B(net620),
    .Q(\mix1.data_o[127] ));
 sky130_fd_sc_hd__dfrtp_1 _18443_ (.CLK(clknet_leaf_9_clk),
    .D(_01873_),
    .RESET_B(net632),
    .Q(\sub1.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _18444_ (.CLK(clknet_leaf_8_clk),
    .D(_01874_),
    .RESET_B(net632),
    .Q(\sub1.state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _18445_ (.CLK(clknet_leaf_9_clk),
    .D(_01875_),
    .RESET_B(net632),
    .Q(\sub1.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _18446_ (.CLK(clknet_leaf_10_clk),
    .D(_01876_),
    .RESET_B(net623),
    .Q(\sub1.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _18447_ (.CLK(clknet_leaf_9_clk),
    .D(_01877_),
    .RESET_B(net631),
    .Q(\sub1.state[4] ));
 sky130_fd_sc_hd__dfrtp_1 _18448_ (.CLK(clknet_leaf_74_clk),
    .D(_01878_),
    .RESET_B(net593),
    .Q(\sub1.data_o[88] ));
 sky130_fd_sc_hd__dfrtp_1 _18449_ (.CLK(clknet_leaf_73_clk),
    .D(_01879_),
    .RESET_B(net593),
    .Q(\sub1.data_o[89] ));
 sky130_fd_sc_hd__dfrtp_1 _18450_ (.CLK(clknet_leaf_70_clk),
    .D(_01880_),
    .RESET_B(net609),
    .Q(\sub1.data_o[90] ));
 sky130_fd_sc_hd__dfrtp_1 _18451_ (.CLK(clknet_leaf_73_clk),
    .D(_01881_),
    .RESET_B(net593),
    .Q(\sub1.data_o[91] ));
 sky130_fd_sc_hd__dfrtp_2 _18452_ (.CLK(clknet_leaf_70_clk),
    .D(_01882_),
    .RESET_B(net608),
    .Q(\sub1.data_o[92] ));
 sky130_fd_sc_hd__dfrtp_2 _18453_ (.CLK(clknet_leaf_70_clk),
    .D(_01883_),
    .RESET_B(net609),
    .Q(\sub1.data_o[93] ));
 sky130_fd_sc_hd__dfrtp_1 _18454_ (.CLK(clknet_leaf_72_clk),
    .D(_01884_),
    .RESET_B(net594),
    .Q(\sub1.data_o[94] ));
 sky130_fd_sc_hd__dfrtp_2 _18455_ (.CLK(clknet_leaf_70_clk),
    .D(_01885_),
    .RESET_B(net609),
    .Q(\sub1.data_o[95] ));
 sky130_fd_sc_hd__dfrtp_4 _18456_ (.CLK(clknet_leaf_27_clk),
    .D(_01886_),
    .RESET_B(net642),
    .Q(\sub1.data_o[96] ));
 sky130_fd_sc_hd__dfrtp_4 _18457_ (.CLK(clknet_leaf_30_clk),
    .D(_01887_),
    .RESET_B(net642),
    .Q(\sub1.data_o[97] ));
 sky130_fd_sc_hd__dfrtp_4 _18458_ (.CLK(clknet_leaf_32_clk),
    .D(_01888_),
    .RESET_B(net653),
    .Q(\sub1.data_o[98] ));
 sky130_fd_sc_hd__dfrtp_4 _18459_ (.CLK(clknet_leaf_27_clk),
    .D(_01889_),
    .RESET_B(net642),
    .Q(\sub1.data_o[99] ));
 sky130_fd_sc_hd__dfrtp_4 _18460_ (.CLK(clknet_leaf_32_clk),
    .D(_01890_),
    .RESET_B(net661),
    .Q(\sub1.data_o[100] ));
 sky130_fd_sc_hd__dfrtp_4 _18461_ (.CLK(clknet_leaf_32_clk),
    .D(_01891_),
    .RESET_B(net661),
    .Q(\sub1.data_o[101] ));
 sky130_fd_sc_hd__dfrtp_4 _18462_ (.CLK(clknet_leaf_34_clk),
    .D(_01892_),
    .RESET_B(net662),
    .Q(\sub1.data_o[102] ));
 sky130_fd_sc_hd__dfrtp_4 _18463_ (.CLK(clknet_leaf_34_clk),
    .D(_01893_),
    .RESET_B(net662),
    .Q(\sub1.data_o[103] ));
 sky130_fd_sc_hd__dfrtp_4 _18464_ (.CLK(clknet_leaf_3_clk),
    .D(_01894_),
    .RESET_B(net583),
    .Q(\sub1.data_o[104] ));
 sky130_fd_sc_hd__dfrtp_4 _18465_ (.CLK(clknet_leaf_83_clk),
    .D(_01895_),
    .RESET_B(net584),
    .Q(\sub1.data_o[105] ));
 sky130_fd_sc_hd__dfrtp_2 _18466_ (.CLK(clknet_leaf_3_clk),
    .D(_01896_),
    .RESET_B(net583),
    .Q(\sub1.data_o[106] ));
 sky130_fd_sc_hd__dfrtp_4 _18467_ (.CLK(clknet_leaf_3_clk),
    .D(_01897_),
    .RESET_B(net584),
    .Q(\sub1.data_o[107] ));
 sky130_fd_sc_hd__dfrtp_2 _18468_ (.CLK(clknet_leaf_3_clk),
    .D(_01898_),
    .RESET_B(net584),
    .Q(\sub1.data_o[108] ));
 sky130_fd_sc_hd__dfrtp_2 _18469_ (.CLK(clknet_leaf_4_clk),
    .D(_01899_),
    .RESET_B(net592),
    .Q(\sub1.data_o[109] ));
 sky130_fd_sc_hd__dfrtp_4 _18470_ (.CLK(clknet_leaf_3_clk),
    .D(_01900_),
    .RESET_B(net583),
    .Q(\sub1.data_o[110] ));
 sky130_fd_sc_hd__dfrtp_4 _18471_ (.CLK(clknet_leaf_83_clk),
    .D(_01901_),
    .RESET_B(net584),
    .Q(\sub1.data_o[111] ));
 sky130_fd_sc_hd__dfrtp_2 _18472_ (.CLK(clknet_leaf_33_clk),
    .D(\mix1.next_ready_o ),
    .RESET_B(net660),
    .Q(\mix1.ready_o ));
 sky130_fd_sc_hd__dfrtp_1 _18473_ (.CLK(clknet_leaf_57_clk),
    .D(_01902_),
    .RESET_B(net602),
    .Q(\ks1.key_reg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _18474_ (.CLK(clknet_leaf_56_clk),
    .D(_01903_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _18475_ (.CLK(clknet_leaf_58_clk),
    .D(_01904_),
    .RESET_B(net602),
    .Q(\ks1.key_reg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _18476_ (.CLK(clknet_leaf_54_clk),
    .D(_01905_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _18477_ (.CLK(clknet_leaf_58_clk),
    .D(_01906_),
    .RESET_B(net602),
    .Q(\ks1.key_reg[4] ));
 sky130_fd_sc_hd__dfrtp_1 _18478_ (.CLK(clknet_leaf_57_clk),
    .D(_01907_),
    .RESET_B(net602),
    .Q(\ks1.key_reg[5] ));
 sky130_fd_sc_hd__dfrtp_1 _18479_ (.CLK(clknet_leaf_55_clk),
    .D(_01908_),
    .RESET_B(net615),
    .Q(\ks1.key_reg[6] ));
 sky130_fd_sc_hd__dfrtp_1 _18480_ (.CLK(clknet_leaf_59_clk),
    .D(_01909_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[7] ));
 sky130_fd_sc_hd__dfrtp_1 _18481_ (.CLK(clknet_leaf_59_clk),
    .D(_01910_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[8] ));
 sky130_fd_sc_hd__dfrtp_1 _18482_ (.CLK(clknet_leaf_57_clk),
    .D(_01911_),
    .RESET_B(net602),
    .Q(\ks1.key_reg[9] ));
 sky130_fd_sc_hd__dfrtp_1 _18483_ (.CLK(clknet_leaf_55_clk),
    .D(_01912_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[10] ));
 sky130_fd_sc_hd__dfrtp_1 _18484_ (.CLK(clknet_leaf_56_clk),
    .D(_01913_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[11] ));
 sky130_fd_sc_hd__dfrtp_1 _18485_ (.CLK(clknet_leaf_57_clk),
    .D(_01914_),
    .RESET_B(net602),
    .Q(\ks1.key_reg[12] ));
 sky130_fd_sc_hd__dfrtp_1 _18486_ (.CLK(clknet_leaf_58_clk),
    .D(_01915_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[13] ));
 sky130_fd_sc_hd__dfrtp_1 _18487_ (.CLK(clknet_leaf_54_clk),
    .D(_01916_),
    .RESET_B(net615),
    .Q(\ks1.key_reg[14] ));
 sky130_fd_sc_hd__dfrtp_1 _18488_ (.CLK(clknet_leaf_56_clk),
    .D(_01917_),
    .RESET_B(net614),
    .Q(\ks1.key_reg[15] ));
 sky130_fd_sc_hd__dfrtp_1 _18489_ (.CLK(clknet_leaf_59_clk),
    .D(_01918_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[16] ));
 sky130_fd_sc_hd__dfrtp_1 _18490_ (.CLK(clknet_leaf_54_clk),
    .D(_01919_),
    .RESET_B(net615),
    .Q(\ks1.key_reg[17] ));
 sky130_fd_sc_hd__dfrtp_1 _18491_ (.CLK(clknet_leaf_55_clk),
    .D(_01920_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[18] ));
 sky130_fd_sc_hd__dfrtp_1 _18492_ (.CLK(clknet_leaf_54_clk),
    .D(_01921_),
    .RESET_B(net614),
    .Q(\ks1.key_reg[19] ));
 sky130_fd_sc_hd__dfrtp_1 _18493_ (.CLK(clknet_leaf_54_clk),
    .D(_01922_),
    .RESET_B(net615),
    .Q(\ks1.key_reg[20] ));
 sky130_fd_sc_hd__dfrtp_1 _18494_ (.CLK(clknet_leaf_56_clk),
    .D(_01923_),
    .RESET_B(net614),
    .Q(\ks1.key_reg[21] ));
 sky130_fd_sc_hd__dfrtp_1 _18495_ (.CLK(clknet_leaf_59_clk),
    .D(_01924_),
    .RESET_B(net613),
    .Q(\ks1.key_reg[22] ));
 sky130_fd_sc_hd__dfrtp_1 _18496_ (.CLK(clknet_leaf_58_clk),
    .D(_01925_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[23] ));
 sky130_fd_sc_hd__dfrtp_1 _18497_ (.CLK(clknet_leaf_59_clk),
    .D(_01926_),
    .RESET_B(net606),
    .Q(\ks1.key_reg[24] ));
 sky130_fd_sc_hd__dfrtp_1 _18498_ (.CLK(clknet_leaf_58_clk),
    .D(_01927_),
    .RESET_B(net602),
    .Q(\ks1.key_reg[25] ));
 sky130_fd_sc_hd__dfrtp_1 _18499_ (.CLK(clknet_leaf_57_clk),
    .D(_01928_),
    .RESET_B(net618),
    .Q(\ks1.key_reg[26] ));
 sky130_fd_sc_hd__dfrtp_1 _18500_ (.CLK(clknet_leaf_55_clk),
    .D(_01929_),
    .RESET_B(net614),
    .Q(\ks1.key_reg[27] ));
 sky130_fd_sc_hd__dfrtp_1 _18501_ (.CLK(clknet_leaf_58_clk),
    .D(_01930_),
    .RESET_B(net618),
    .Q(\ks1.key_reg[28] ));
 sky130_fd_sc_hd__dfrtp_1 _18502_ (.CLK(clknet_leaf_58_clk),
    .D(_01931_),
    .RESET_B(net618),
    .Q(\ks1.key_reg[29] ));
 sky130_fd_sc_hd__dfrtp_1 _18503_ (.CLK(clknet_leaf_59_clk),
    .D(_01932_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[30] ));
 sky130_fd_sc_hd__dfrtp_1 _18504_ (.CLK(clknet_leaf_61_clk),
    .D(_01933_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[31] ));
 sky130_fd_sc_hd__dfrtp_1 _18505_ (.CLK(clknet_leaf_58_clk),
    .D(_01934_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[32] ));
 sky130_fd_sc_hd__dfrtp_1 _18506_ (.CLK(clknet_leaf_59_clk),
    .D(_01935_),
    .RESET_B(net606),
    .Q(\ks1.key_reg[33] ));
 sky130_fd_sc_hd__dfrtp_1 _18507_ (.CLK(clknet_leaf_61_clk),
    .D(_01936_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[34] ));
 sky130_fd_sc_hd__dfrtp_1 _18508_ (.CLK(clknet_leaf_67_clk),
    .D(_01937_),
    .RESET_B(net606),
    .Q(\ks1.key_reg[35] ));
 sky130_fd_sc_hd__dfrtp_1 _18509_ (.CLK(clknet_leaf_62_clk),
    .D(_01938_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[36] ));
 sky130_fd_sc_hd__dfrtp_1 _18510_ (.CLK(clknet_leaf_62_clk),
    .D(_01939_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[37] ));
 sky130_fd_sc_hd__dfrtp_1 _18511_ (.CLK(clknet_leaf_62_clk),
    .D(_01940_),
    .RESET_B(net598),
    .Q(\ks1.key_reg[38] ));
 sky130_fd_sc_hd__dfrtp_1 _18512_ (.CLK(clknet_leaf_66_clk),
    .D(_01941_),
    .RESET_B(net604),
    .Q(\ks1.key_reg[39] ));
 sky130_fd_sc_hd__dfrtp_1 _18513_ (.CLK(clknet_leaf_59_clk),
    .D(_01942_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[40] ));
 sky130_fd_sc_hd__dfrtp_1 _18514_ (.CLK(clknet_leaf_62_clk),
    .D(_01943_),
    .RESET_B(net598),
    .Q(\ks1.key_reg[41] ));
 sky130_fd_sc_hd__dfrtp_1 _18515_ (.CLK(clknet_leaf_65_clk),
    .D(_01944_),
    .RESET_B(net604),
    .Q(\ks1.key_reg[42] ));
 sky130_fd_sc_hd__dfrtp_1 _18516_ (.CLK(clknet_leaf_62_clk),
    .D(_01945_),
    .RESET_B(net599),
    .Q(\ks1.key_reg[43] ));
 sky130_fd_sc_hd__dfrtp_1 _18517_ (.CLK(clknet_leaf_63_clk),
    .D(_01946_),
    .RESET_B(net599),
    .Q(\ks1.key_reg[44] ));
 sky130_fd_sc_hd__dfrtp_1 _18518_ (.CLK(clknet_leaf_64_clk),
    .D(_01947_),
    .RESET_B(net603),
    .Q(\ks1.key_reg[45] ));
 sky130_fd_sc_hd__dfrtp_1 _18519_ (.CLK(clknet_leaf_64_clk),
    .D(_01948_),
    .RESET_B(net607),
    .Q(\ks1.key_reg[46] ));
 sky130_fd_sc_hd__dfrtp_1 _18520_ (.CLK(clknet_leaf_66_clk),
    .D(_01949_),
    .RESET_B(net606),
    .Q(\ks1.key_reg[47] ));
 sky130_fd_sc_hd__dfrtp_1 _18521_ (.CLK(clknet_leaf_66_clk),
    .D(_01950_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[48] ));
 sky130_fd_sc_hd__dfrtp_1 _18522_ (.CLK(clknet_leaf_67_clk),
    .D(_01951_),
    .RESET_B(net606),
    .Q(\ks1.key_reg[49] ));
 sky130_fd_sc_hd__dfrtp_1 _18523_ (.CLK(clknet_leaf_67_clk),
    .D(_01952_),
    .RESET_B(net606),
    .Q(\ks1.key_reg[50] ));
 sky130_fd_sc_hd__dfrtp_1 _18524_ (.CLK(clknet_leaf_67_clk),
    .D(_01953_),
    .RESET_B(net610),
    .Q(\ks1.key_reg[51] ));
 sky130_fd_sc_hd__dfrtp_1 _18525_ (.CLK(clknet_leaf_67_clk),
    .D(_01954_),
    .RESET_B(net606),
    .Q(\ks1.key_reg[52] ));
 sky130_fd_sc_hd__dfrtp_1 _18526_ (.CLK(clknet_leaf_66_clk),
    .D(_01955_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[53] ));
 sky130_fd_sc_hd__dfrtp_1 _18527_ (.CLK(clknet_leaf_60_clk),
    .D(_01956_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[54] ));
 sky130_fd_sc_hd__dfrtp_1 _18528_ (.CLK(clknet_leaf_60_clk),
    .D(_01957_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[55] ));
 sky130_fd_sc_hd__dfrtp_1 _18529_ (.CLK(clknet_leaf_66_clk),
    .D(_01958_),
    .RESET_B(net606),
    .Q(\ks1.key_reg[56] ));
 sky130_fd_sc_hd__dfrtp_1 _18530_ (.CLK(clknet_leaf_60_clk),
    .D(_01959_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[57] ));
 sky130_fd_sc_hd__dfrtp_1 _18531_ (.CLK(clknet_leaf_62_clk),
    .D(_01960_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[58] ));
 sky130_fd_sc_hd__dfrtp_1 _18532_ (.CLK(clknet_leaf_59_clk),
    .D(_01961_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[59] ));
 sky130_fd_sc_hd__dfrtp_1 _18533_ (.CLK(clknet_leaf_61_clk),
    .D(_01962_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[60] ));
 sky130_fd_sc_hd__dfrtp_1 _18534_ (.CLK(clknet_leaf_61_clk),
    .D(_01963_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[61] ));
 sky130_fd_sc_hd__dfrtp_1 _18535_ (.CLK(clknet_leaf_60_clk),
    .D(_01964_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[62] ));
 sky130_fd_sc_hd__dfrtp_1 _18536_ (.CLK(clknet_leaf_61_clk),
    .D(_01965_),
    .RESET_B(net600),
    .Q(\ks1.key_reg[63] ));
 sky130_fd_sc_hd__dfrtp_1 _18537_ (.CLK(clknet_leaf_60_clk),
    .D(_01966_),
    .RESET_B(net601),
    .Q(\ks1.key_reg[64] ));
 sky130_fd_sc_hd__dfrtp_1 _18538_ (.CLK(clknet_leaf_60_clk),
    .D(_01967_),
    .RESET_B(net601),
    .Q(\ks1.key_reg[65] ));
 sky130_fd_sc_hd__dfrtp_1 _18539_ (.CLK(clknet_leaf_60_clk),
    .D(_01968_),
    .RESET_B(net605),
    .Q(\ks1.key_reg[66] ));
 sky130_fd_sc_hd__dfrtp_1 _18540_ (.CLK(clknet_leaf_66_clk),
    .D(_01969_),
    .RESET_B(net606),
    .Q(\ks1.key_reg[67] ));
 sky130_fd_sc_hd__dfrtp_1 _18541_ (.CLK(clknet_leaf_62_clk),
    .D(_01970_),
    .RESET_B(net601),
    .Q(\ks1.key_reg[68] ));
 sky130_fd_sc_hd__dfrtp_1 _18542_ (.CLK(clknet_leaf_79_clk),
    .D(_01971_),
    .RESET_B(net579),
    .Q(\ks1.key_reg[69] ));
 sky130_fd_sc_hd__dfrtp_1 _18543_ (.CLK(clknet_leaf_79_clk),
    .D(_01972_),
    .RESET_B(net579),
    .Q(\ks1.key_reg[70] ));
 sky130_fd_sc_hd__dfrtp_1 _18544_ (.CLK(clknet_leaf_63_clk),
    .D(_01973_),
    .RESET_B(net599),
    .Q(\ks1.key_reg[71] ));
 sky130_fd_sc_hd__dfrtp_1 _18545_ (.CLK(clknet_leaf_65_clk),
    .D(_01974_),
    .RESET_B(net603),
    .Q(\ks1.key_reg[72] ));
 sky130_fd_sc_hd__dfrtp_1 _18546_ (.CLK(clknet_leaf_63_clk),
    .D(_01975_),
    .RESET_B(net599),
    .Q(\ks1.key_reg[73] ));
 sky130_fd_sc_hd__dfrtp_1 _18547_ (.CLK(clknet_leaf_77_clk),
    .D(_01976_),
    .RESET_B(net589),
    .Q(\ks1.key_reg[74] ));
 sky130_fd_sc_hd__dfrtp_1 _18548_ (.CLK(clknet_leaf_64_clk),
    .D(_01977_),
    .RESET_B(net599),
    .Q(\ks1.key_reg[75] ));
 sky130_fd_sc_hd__dfrtp_1 _18549_ (.CLK(clknet_leaf_78_clk),
    .D(_01978_),
    .RESET_B(net579),
    .Q(\ks1.key_reg[76] ));
 sky130_fd_sc_hd__dfrtp_1 _18550_ (.CLK(clknet_leaf_64_clk),
    .D(_01979_),
    .RESET_B(net603),
    .Q(\ks1.key_reg[77] ));
 sky130_fd_sc_hd__dfrtp_1 _18551_ (.CLK(clknet_leaf_78_clk),
    .D(_01980_),
    .RESET_B(net580),
    .Q(\ks1.key_reg[78] ));
 sky130_fd_sc_hd__dfrtp_1 _18552_ (.CLK(clknet_leaf_64_clk),
    .D(_01981_),
    .RESET_B(net599),
    .Q(\ks1.key_reg[79] ));
 sky130_fd_sc_hd__dfrtp_1 _18553_ (.CLK(clknet_leaf_78_clk),
    .D(_01982_),
    .RESET_B(net589),
    .Q(\ks1.key_reg[80] ));
 sky130_fd_sc_hd__dfrtp_1 _18554_ (.CLK(clknet_leaf_77_clk),
    .D(_01983_),
    .RESET_B(net589),
    .Q(\ks1.key_reg[81] ));
 sky130_fd_sc_hd__dfrtp_1 _18555_ (.CLK(clknet_leaf_77_clk),
    .D(_01984_),
    .RESET_B(net590),
    .Q(\ks1.key_reg[82] ));
 sky130_fd_sc_hd__dfrtp_1 _18556_ (.CLK(clknet_leaf_77_clk),
    .D(_01985_),
    .RESET_B(net590),
    .Q(\ks1.key_reg[83] ));
 sky130_fd_sc_hd__dfrtp_1 _18557_ (.CLK(clknet_leaf_78_clk),
    .D(_01986_),
    .RESET_B(net589),
    .Q(\ks1.key_reg[84] ));
 sky130_fd_sc_hd__dfrtp_1 _18558_ (.CLK(clknet_leaf_65_clk),
    .D(_01987_),
    .RESET_B(net589),
    .Q(\ks1.key_reg[85] ));
 sky130_fd_sc_hd__dfrtp_1 _18559_ (.CLK(clknet_leaf_76_clk),
    .D(_01988_),
    .RESET_B(net590),
    .Q(\ks1.key_reg[86] ));
 sky130_fd_sc_hd__dfrtp_1 _18560_ (.CLK(clknet_leaf_64_clk),
    .D(_01989_),
    .RESET_B(net603),
    .Q(\ks1.key_reg[87] ));
 sky130_fd_sc_hd__dfrtp_1 _18561_ (.CLK(clknet_leaf_65_clk),
    .D(_01990_),
    .RESET_B(net604),
    .Q(\ks1.key_reg[88] ));
 sky130_fd_sc_hd__dfrtp_1 _18562_ (.CLK(clknet_leaf_63_clk),
    .D(_01991_),
    .RESET_B(net598),
    .Q(\ks1.key_reg[89] ));
 sky130_fd_sc_hd__dfrtp_1 _18563_ (.CLK(clknet_leaf_63_clk),
    .D(_01992_),
    .RESET_B(net598),
    .Q(\ks1.key_reg[90] ));
 sky130_fd_sc_hd__dfrtp_1 _18564_ (.CLK(clknet_leaf_63_clk),
    .D(_01993_),
    .RESET_B(net598),
    .Q(\ks1.key_reg[91] ));
 sky130_fd_sc_hd__dfrtp_1 _18565_ (.CLK(clknet_leaf_63_clk),
    .D(_01994_),
    .RESET_B(net598),
    .Q(\ks1.key_reg[92] ));
 sky130_fd_sc_hd__dfrtp_1 _18566_ (.CLK(clknet_leaf_62_clk),
    .D(_01995_),
    .RESET_B(net598),
    .Q(\ks1.key_reg[93] ));
 sky130_fd_sc_hd__dfrtp_1 _18567_ (.CLK(clknet_leaf_66_clk),
    .D(_01996_),
    .RESET_B(net604),
    .Q(\ks1.key_reg[94] ));
 sky130_fd_sc_hd__dfrtp_1 _18568_ (.CLK(clknet_leaf_63_clk),
    .D(_01997_),
    .RESET_B(net598),
    .Q(\ks1.key_reg[95] ));
 sky130_fd_sc_hd__dfrtp_1 _18569_ (.CLK(clknet_leaf_64_clk),
    .D(_01998_),
    .RESET_B(net599),
    .Q(\ks1.key_reg[96] ));
 sky130_fd_sc_hd__dfrtp_1 _18570_ (.CLK(clknet_leaf_80_clk),
    .D(_01999_),
    .RESET_B(net580),
    .Q(\ks1.key_reg[97] ));
 sky130_fd_sc_hd__dfrtp_1 _18571_ (.CLK(clknet_leaf_81_clk),
    .D(_02000_),
    .RESET_B(net586),
    .Q(\ks1.key_reg[98] ));
 sky130_fd_sc_hd__dfrtp_1 _18572_ (.CLK(clknet_leaf_82_clk),
    .D(_02001_),
    .RESET_B(net587),
    .Q(\ks1.key_reg[99] ));
 sky130_fd_sc_hd__dfrtp_1 _18573_ (.CLK(clknet_leaf_81_clk),
    .D(_02002_),
    .RESET_B(net578),
    .Q(\ks1.key_reg[100] ));
 sky130_fd_sc_hd__dfrtp_1 _18574_ (.CLK(clknet_leaf_81_clk),
    .D(_02003_),
    .RESET_B(net578),
    .Q(\ks1.key_reg[101] ));
 sky130_fd_sc_hd__dfrtp_1 _18575_ (.CLK(clknet_leaf_75_clk),
    .D(_02004_),
    .RESET_B(net587),
    .Q(\ks1.key_reg[102] ));
 sky130_fd_sc_hd__dfrtp_1 _18576_ (.CLK(clknet_leaf_80_clk),
    .D(_02005_),
    .RESET_B(net580),
    .Q(\ks1.key_reg[103] ));
 sky130_fd_sc_hd__dfrtp_1 _18577_ (.CLK(clknet_leaf_75_clk),
    .D(_02006_),
    .RESET_B(net587),
    .Q(\ks1.key_reg[104] ));
 sky130_fd_sc_hd__dfrtp_1 _18578_ (.CLK(clknet_leaf_64_clk),
    .D(_02007_),
    .RESET_B(net603),
    .Q(\ks1.key_reg[105] ));
 sky130_fd_sc_hd__dfrtp_1 _18579_ (.CLK(clknet_leaf_77_clk),
    .D(_02008_),
    .RESET_B(net589),
    .Q(\ks1.key_reg[106] ));
 sky130_fd_sc_hd__dfrtp_1 _18580_ (.CLK(clknet_leaf_75_clk),
    .D(_02009_),
    .RESET_B(net588),
    .Q(\ks1.key_reg[107] ));
 sky130_fd_sc_hd__dfrtp_1 _18581_ (.CLK(clknet_leaf_65_clk),
    .D(_02010_),
    .RESET_B(net590),
    .Q(\ks1.key_reg[108] ));
 sky130_fd_sc_hd__dfrtp_1 _18582_ (.CLK(clknet_leaf_65_clk),
    .D(_02011_),
    .RESET_B(net590),
    .Q(\ks1.key_reg[109] ));
 sky130_fd_sc_hd__dfrtp_1 _18583_ (.CLK(clknet_leaf_78_clk),
    .D(_02012_),
    .RESET_B(net580),
    .Q(\ks1.key_reg[110] ));
 sky130_fd_sc_hd__dfrtp_1 _18584_ (.CLK(clknet_leaf_81_clk),
    .D(_02013_),
    .RESET_B(net578),
    .Q(\ks1.key_reg[111] ));
 sky130_fd_sc_hd__dfrtp_1 _18585_ (.CLK(clknet_leaf_81_clk),
    .D(_02014_),
    .RESET_B(net588),
    .Q(\ks1.key_reg[112] ));
 sky130_fd_sc_hd__dfrtp_1 _18586_ (.CLK(clknet_leaf_76_clk),
    .D(_02015_),
    .RESET_B(net589),
    .Q(\ks1.key_reg[113] ));
 sky130_fd_sc_hd__dfrtp_1 _18587_ (.CLK(clknet_leaf_75_clk),
    .D(_02016_),
    .RESET_B(net587),
    .Q(\ks1.key_reg[114] ));
 sky130_fd_sc_hd__dfrtp_1 _18588_ (.CLK(clknet_leaf_74_clk),
    .D(_02017_),
    .RESET_B(net588),
    .Q(\ks1.key_reg[115] ));
 sky130_fd_sc_hd__dfrtp_1 _18589_ (.CLK(clknet_leaf_81_clk),
    .D(_02018_),
    .RESET_B(net586),
    .Q(\ks1.key_reg[116] ));
 sky130_fd_sc_hd__dfrtp_1 _18590_ (.CLK(clknet_leaf_76_clk),
    .D(_02019_),
    .RESET_B(net588),
    .Q(\ks1.key_reg[117] ));
 sky130_fd_sc_hd__dfrtp_1 _18591_ (.CLK(clknet_leaf_75_clk),
    .D(_02020_),
    .RESET_B(net587),
    .Q(\ks1.key_reg[118] ));
 sky130_fd_sc_hd__dfrtp_1 _18592_ (.CLK(clknet_leaf_77_clk),
    .D(_02021_),
    .RESET_B(net589),
    .Q(\ks1.key_reg[119] ));
 sky130_fd_sc_hd__dfrtp_1 _18593_ (.CLK(clknet_leaf_65_clk),
    .D(_02022_),
    .RESET_B(net604),
    .Q(\ks1.key_reg[120] ));
 sky130_fd_sc_hd__dfrtp_1 _18594_ (.CLK(clknet_leaf_69_clk),
    .D(_02023_),
    .RESET_B(net608),
    .Q(\ks1.key_reg[121] ));
 sky130_fd_sc_hd__dfrtp_1 _18595_ (.CLK(clknet_leaf_69_clk),
    .D(_02024_),
    .RESET_B(net607),
    .Q(\ks1.key_reg[122] ));
 sky130_fd_sc_hd__dfrtp_1 _18596_ (.CLK(clknet_leaf_65_clk),
    .D(_02025_),
    .RESET_B(net604),
    .Q(\ks1.key_reg[123] ));
 sky130_fd_sc_hd__dfrtp_1 _18597_ (.CLK(clknet_leaf_67_clk),
    .D(_02026_),
    .RESET_B(net610),
    .Q(\ks1.key_reg[124] ));
 sky130_fd_sc_hd__dfrtp_1 _18598_ (.CLK(clknet_leaf_68_clk),
    .D(_02027_),
    .RESET_B(net608),
    .Q(\ks1.key_reg[125] ));
 sky130_fd_sc_hd__dfrtp_1 _18599_ (.CLK(clknet_leaf_68_clk),
    .D(_02028_),
    .RESET_B(net608),
    .Q(\ks1.key_reg[126] ));
 sky130_fd_sc_hd__dfrtp_1 _18600_ (.CLK(clknet_leaf_69_clk),
    .D(_02029_),
    .RESET_B(net604),
    .Q(\ks1.key_reg[127] ));
 sky130_fd_sc_hd__dfrtp_2 _18601_ (.CLK(clknet_leaf_33_clk),
    .D(_02030_),
    .RESET_B(net660),
    .Q(\mix1.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _18602_ (.CLK(clknet_leaf_14_clk),
    .D(_02031_),
    .RESET_B(net629),
    .Q(\mix1.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _18603_ (.CLK(clknet_leaf_13_clk),
    .D(_02032_),
    .RESET_B(net628),
    .Q(\mix1.data_reg[96] ));
 sky130_fd_sc_hd__dfrtp_1 _18604_ (.CLK(clknet_leaf_14_clk),
    .D(_02033_),
    .RESET_B(net630),
    .Q(\mix1.data_reg[97] ));
 sky130_fd_sc_hd__dfrtp_1 _18605_ (.CLK(clknet_leaf_14_clk),
    .D(_02034_),
    .RESET_B(net630),
    .Q(\mix1.data_reg[98] ));
 sky130_fd_sc_hd__dfrtp_1 _18606_ (.CLK(clknet_leaf_14_clk),
    .D(_02035_),
    .RESET_B(net630),
    .Q(\mix1.data_reg[99] ));
 sky130_fd_sc_hd__dfrtp_1 _18607_ (.CLK(clknet_leaf_14_clk),
    .D(_02036_),
    .RESET_B(net629),
    .Q(\mix1.data_reg[100] ));
 sky130_fd_sc_hd__dfrtp_1 _18608_ (.CLK(clknet_leaf_13_clk),
    .D(_02037_),
    .RESET_B(net627),
    .Q(\mix1.data_reg[101] ));
 sky130_fd_sc_hd__dfrtp_1 _18609_ (.CLK(clknet_leaf_13_clk),
    .D(_02038_),
    .RESET_B(net627),
    .Q(\mix1.data_reg[102] ));
 sky130_fd_sc_hd__dfrtp_1 _18610_ (.CLK(clknet_leaf_13_clk),
    .D(_02039_),
    .RESET_B(net627),
    .Q(\mix1.data_reg[103] ));
 sky130_fd_sc_hd__dfrtp_1 _18611_ (.CLK(clknet_leaf_12_clk),
    .D(_02040_),
    .RESET_B(net621),
    .Q(\mix1.data_reg[104] ));
 sky130_fd_sc_hd__dfrtp_1 _18612_ (.CLK(clknet_leaf_12_clk),
    .D(_02041_),
    .RESET_B(net628),
    .Q(\mix1.data_reg[105] ));
 sky130_fd_sc_hd__dfrtp_1 _18613_ (.CLK(clknet_leaf_84_clk),
    .D(_02042_),
    .RESET_B(net581),
    .Q(\mix1.data_reg[106] ));
 sky130_fd_sc_hd__dfrtp_1 _18614_ (.CLK(clknet_leaf_83_clk),
    .D(_02043_),
    .RESET_B(net582),
    .Q(\mix1.data_reg[107] ));
 sky130_fd_sc_hd__dfrtp_1 _18615_ (.CLK(clknet_leaf_83_clk),
    .D(_02044_),
    .RESET_B(net582),
    .Q(\mix1.data_reg[108] ));
 sky130_fd_sc_hd__dfrtp_1 _18616_ (.CLK(clknet_leaf_83_clk),
    .D(_02045_),
    .RESET_B(net584),
    .Q(\mix1.data_reg[109] ));
 sky130_fd_sc_hd__dfrtp_1 _18617_ (.CLK(clknet_leaf_83_clk),
    .D(_02046_),
    .RESET_B(net583),
    .Q(\mix1.data_reg[110] ));
 sky130_fd_sc_hd__dfrtp_1 _18618_ (.CLK(clknet_leaf_0_clk),
    .D(_02047_),
    .RESET_B(net619),
    .Q(\mix1.data_reg[111] ));
 sky130_fd_sc_hd__dfrtp_1 _18619_ (.CLK(clknet_leaf_15_clk),
    .D(_02048_),
    .RESET_B(net636),
    .Q(\mix1.data_reg[112] ));
 sky130_fd_sc_hd__dfrtp_1 _18620_ (.CLK(clknet_leaf_15_clk),
    .D(_02049_),
    .RESET_B(net636),
    .Q(\mix1.data_reg[113] ));
 sky130_fd_sc_hd__dfrtp_1 _18621_ (.CLK(clknet_leaf_16_clk),
    .D(_02050_),
    .RESET_B(net634),
    .Q(\mix1.data_reg[114] ));
 sky130_fd_sc_hd__dfrtp_1 _18622_ (.CLK(clknet_leaf_20_clk),
    .D(_02051_),
    .RESET_B(net640),
    .Q(\mix1.data_reg[115] ));
 sky130_fd_sc_hd__dfrtp_1 _18623_ (.CLK(clknet_leaf_23_clk),
    .D(_02052_),
    .RESET_B(net644),
    .Q(\mix1.data_reg[116] ));
 sky130_fd_sc_hd__dfrtp_1 _18624_ (.CLK(clknet_leaf_24_clk),
    .D(_02053_),
    .RESET_B(net645),
    .Q(\mix1.data_reg[117] ));
 sky130_fd_sc_hd__dfrtp_1 _18625_ (.CLK(clknet_leaf_23_clk),
    .D(_02054_),
    .RESET_B(net644),
    .Q(\mix1.data_reg[118] ));
 sky130_fd_sc_hd__dfrtp_1 _18626_ (.CLK(clknet_leaf_24_clk),
    .D(_02055_),
    .RESET_B(net645),
    .Q(\mix1.data_reg[119] ));
 sky130_fd_sc_hd__dfrtp_1 _18627_ (.CLK(clknet_leaf_23_clk),
    .D(_02056_),
    .RESET_B(net645),
    .Q(\mix1.data_reg[120] ));
 sky130_fd_sc_hd__dfrtp_1 _18628_ (.CLK(clknet_leaf_25_clk),
    .D(_02057_),
    .RESET_B(net648),
    .Q(\mix1.data_reg[121] ));
 sky130_fd_sc_hd__dfrtp_1 _18629_ (.CLK(clknet_leaf_23_clk),
    .D(_02058_),
    .RESET_B(net644),
    .Q(\mix1.data_reg[122] ));
 sky130_fd_sc_hd__dfrtp_1 _18630_ (.CLK(clknet_leaf_36_clk),
    .D(_02059_),
    .RESET_B(net666),
    .Q(\mix1.data_reg[123] ));
 sky130_fd_sc_hd__dfrtp_1 _18631_ (.CLK(clknet_leaf_36_clk),
    .D(_02060_),
    .RESET_B(net666),
    .Q(\mix1.data_reg[124] ));
 sky130_fd_sc_hd__dfrtp_1 _18632_ (.CLK(clknet_leaf_36_clk),
    .D(_02061_),
    .RESET_B(net665),
    .Q(\mix1.data_reg[125] ));
 sky130_fd_sc_hd__dfrtp_1 _18633_ (.CLK(clknet_leaf_1_clk),
    .D(_02062_),
    .RESET_B(net622),
    .Q(\mix1.data_reg[126] ));
 sky130_fd_sc_hd__dfrtp_1 _18634_ (.CLK(clknet_leaf_0_clk),
    .D(_02063_),
    .RESET_B(net620),
    .Q(\mix1.data_reg[127] ));
 sky130_fd_sc_hd__dfrtp_4 _18635_ (.CLK(clknet_leaf_21_clk),
    .D(_02064_),
    .RESET_B(net639),
    .Q(\sub1.data_o[112] ));
 sky130_fd_sc_hd__dfrtp_4 _18636_ (.CLK(clknet_leaf_21_clk),
    .D(_02065_),
    .RESET_B(net639),
    .Q(\sub1.data_o[113] ));
 sky130_fd_sc_hd__dfrtp_4 _18637_ (.CLK(clknet_leaf_21_clk),
    .D(_02066_),
    .RESET_B(net639),
    .Q(\sub1.data_o[114] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_2 fanout389 (.A(net391),
    .X(net389));
 sky130_fd_sc_hd__buf_1 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_2 fanout391 (.A(net444),
    .X(net391));
 sky130_fd_sc_hd__buf_2 fanout392 (.A(net397),
    .X(net392));
 sky130_fd_sc_hd__buf_2 fanout393 (.A(net397),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_2 fanout394 (.A(net397),
    .X(net394));
 sky130_fd_sc_hd__buf_2 fanout395 (.A(net397),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_2 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__buf_2 fanout397 (.A(net444),
    .X(net397));
 sky130_fd_sc_hd__buf_2 fanout398 (.A(net404),
    .X(net398));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout399 (.A(net404),
    .X(net399));
 sky130_fd_sc_hd__buf_2 fanout400 (.A(net404),
    .X(net400));
 sky130_fd_sc_hd__buf_2 fanout401 (.A(net404),
    .X(net401));
 sky130_fd_sc_hd__buf_2 fanout402 (.A(net404),
    .X(net402));
 sky130_fd_sc_hd__buf_1 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_2 fanout404 (.A(net444),
    .X(net404));
 sky130_fd_sc_hd__buf_2 fanout405 (.A(net413),
    .X(net405));
 sky130_fd_sc_hd__buf_1 fanout406 (.A(net413),
    .X(net406));
 sky130_fd_sc_hd__buf_2 fanout407 (.A(net413),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 fanout408 (.A(net413),
    .X(net408));
 sky130_fd_sc_hd__buf_2 fanout409 (.A(net413),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_2 fanout410 (.A(net413),
    .X(net410));
 sky130_fd_sc_hd__buf_2 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__buf_2 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__buf_2 fanout413 (.A(net444),
    .X(net413));
 sky130_fd_sc_hd__buf_2 fanout414 (.A(net419),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_2 fanout415 (.A(net419),
    .X(net415));
 sky130_fd_sc_hd__buf_2 fanout416 (.A(net419),
    .X(net416));
 sky130_fd_sc_hd__buf_2 fanout417 (.A(net419),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_2 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__buf_2 fanout419 (.A(net444),
    .X(net419));
 sky130_fd_sc_hd__buf_2 fanout420 (.A(net427),
    .X(net420));
 sky130_fd_sc_hd__buf_1 fanout421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__buf_2 fanout422 (.A(net427),
    .X(net422));
 sky130_fd_sc_hd__buf_2 fanout423 (.A(net427),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 fanout424 (.A(net427),
    .X(net424));
 sky130_fd_sc_hd__buf_2 fanout425 (.A(net427),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_2 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_2 fanout427 (.A(net444),
    .X(net427));
 sky130_fd_sc_hd__buf_2 fanout428 (.A(net431),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 fanout429 (.A(net431),
    .X(net429));
 sky130_fd_sc_hd__buf_2 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 fanout431 (.A(net436),
    .X(net431));
 sky130_fd_sc_hd__buf_2 fanout432 (.A(net436),
    .X(net432));
 sky130_fd_sc_hd__buf_1 fanout433 (.A(net436),
    .X(net433));
 sky130_fd_sc_hd__buf_2 fanout434 (.A(net436),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_2 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 fanout436 (.A(net444),
    .X(net436));
 sky130_fd_sc_hd__buf_2 fanout437 (.A(net443),
    .X(net437));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout438 (.A(net443),
    .X(net438));
 sky130_fd_sc_hd__buf_2 fanout439 (.A(net443),
    .X(net439));
 sky130_fd_sc_hd__buf_1 fanout440 (.A(net443),
    .X(net440));
 sky130_fd_sc_hd__buf_2 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__buf_2 fanout442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_2 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_4 fanout444 (.A(\fifo_bank_register.clk ),
    .X(net444));
 sky130_fd_sc_hd__buf_2 fanout445 (.A(net449),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_2 fanout446 (.A(net449),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_2 fanout447 (.A(net449),
    .X(net447));
 sky130_fd_sc_hd__buf_2 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_2 fanout449 (.A(net461),
    .X(net449));
 sky130_fd_sc_hd__buf_2 fanout450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_2 fanout451 (.A(net461),
    .X(net451));
 sky130_fd_sc_hd__buf_2 fanout452 (.A(net461),
    .X(net452));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout453 (.A(net461),
    .X(net453));
 sky130_fd_sc_hd__buf_2 fanout454 (.A(net460),
    .X(net454));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout455 (.A(net460),
    .X(net455));
 sky130_fd_sc_hd__buf_2 fanout456 (.A(net460),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_2 fanout457 (.A(net460),
    .X(net457));
 sky130_fd_sc_hd__buf_2 fanout458 (.A(net460),
    .X(net458));
 sky130_fd_sc_hd__buf_1 fanout459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_2 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_2 fanout461 (.A(net472),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_2 fanout462 (.A(net466),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_2 fanout463 (.A(net466),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_2 fanout464 (.A(net466),
    .X(net464));
 sky130_fd_sc_hd__buf_2 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__buf_2 fanout466 (.A(net472),
    .X(net466));
 sky130_fd_sc_hd__buf_2 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout468 (.A(net472),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_2 fanout469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__buf_2 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_2 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_2 fanout472 (.A(\fifo_bank_register.clk ),
    .X(net472));
 sky130_fd_sc_hd__buf_2 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__buf_2 fanout474 (.A(net481),
    .X(net474));
 sky130_fd_sc_hd__buf_2 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_2 fanout476 (.A(net481),
    .X(net476));
 sky130_fd_sc_hd__buf_2 fanout477 (.A(net481),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_2 fanout478 (.A(net481),
    .X(net478));
 sky130_fd_sc_hd__buf_2 fanout479 (.A(net481),
    .X(net479));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_2 fanout481 (.A(net530),
    .X(net481));
 sky130_fd_sc_hd__buf_2 fanout482 (.A(net484),
    .X(net482));
 sky130_fd_sc_hd__buf_2 fanout483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_2 fanout484 (.A(net489),
    .X(net484));
 sky130_fd_sc_hd__buf_2 fanout485 (.A(net489),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_2 fanout486 (.A(net489),
    .X(net486));
 sky130_fd_sc_hd__buf_2 fanout487 (.A(net489),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_2 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_2 fanout489 (.A(net530),
    .X(net489));
 sky130_fd_sc_hd__buf_2 fanout490 (.A(net498),
    .X(net490));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout491 (.A(net498),
    .X(net491));
 sky130_fd_sc_hd__buf_2 fanout492 (.A(net498),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_2 fanout493 (.A(net498),
    .X(net493));
 sky130_fd_sc_hd__buf_2 fanout494 (.A(net498),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_2 fanout495 (.A(net498),
    .X(net495));
 sky130_fd_sc_hd__buf_2 fanout496 (.A(net498),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_2 fanout497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__buf_2 fanout498 (.A(net530),
    .X(net498));
 sky130_fd_sc_hd__buf_2 fanout499 (.A(net507),
    .X(net499));
 sky130_fd_sc_hd__buf_2 fanout500 (.A(net507),
    .X(net500));
 sky130_fd_sc_hd__buf_2 fanout501 (.A(net507),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_2 fanout502 (.A(net507),
    .X(net502));
 sky130_fd_sc_hd__buf_2 fanout503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__buf_2 fanout504 (.A(net507),
    .X(net504));
 sky130_fd_sc_hd__buf_2 fanout505 (.A(net507),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_2 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__buf_2 fanout507 (.A(net530),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_2 fanout508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__clkbuf_2 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout510 (.A(net511),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_2 fanout511 (.A(net530),
    .X(net511));
 sky130_fd_sc_hd__buf_2 fanout512 (.A(net520),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_2 fanout513 (.A(net520),
    .X(net513));
 sky130_fd_sc_hd__buf_2 fanout514 (.A(net520),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_2 fanout515 (.A(net520),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_2 fanout516 (.A(net520),
    .X(net516));
 sky130_fd_sc_hd__buf_2 fanout517 (.A(net520),
    .X(net517));
 sky130_fd_sc_hd__buf_2 fanout518 (.A(net520),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_2 fanout519 (.A(net520),
    .X(net519));
 sky130_fd_sc_hd__buf_2 fanout520 (.A(net530),
    .X(net520));
 sky130_fd_sc_hd__buf_2 fanout521 (.A(net529),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_2 fanout522 (.A(net529),
    .X(net522));
 sky130_fd_sc_hd__buf_2 fanout523 (.A(net529),
    .X(net523));
 sky130_fd_sc_hd__clkbuf_2 fanout524 (.A(net529),
    .X(net524));
 sky130_fd_sc_hd__buf_2 fanout525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__buf_2 fanout526 (.A(net528),
    .X(net526));
 sky130_fd_sc_hd__buf_2 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_2 fanout528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_4 fanout530 (.A(\fifo_bank_register.clk ),
    .X(net530));
 sky130_fd_sc_hd__buf_2 fanout531 (.A(net537),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_2 fanout532 (.A(net537),
    .X(net532));
 sky130_fd_sc_hd__buf_2 fanout533 (.A(net535),
    .X(net533));
 sky130_fd_sc_hd__buf_2 fanout534 (.A(net535),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_2 fanout535 (.A(net537),
    .X(net535));
 sky130_fd_sc_hd__buf_2 fanout536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__buf_2 fanout537 (.A(net577),
    .X(net537));
 sky130_fd_sc_hd__buf_2 fanout538 (.A(net542),
    .X(net538));
 sky130_fd_sc_hd__buf_1 fanout539 (.A(net542),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_2 fanout540 (.A(net542),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_2 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_2 fanout542 (.A(net577),
    .X(net542));
 sky130_fd_sc_hd__buf_2 fanout543 (.A(net551),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_2 fanout544 (.A(net551),
    .X(net544));
 sky130_fd_sc_hd__buf_2 fanout545 (.A(net551),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_2 fanout546 (.A(net551),
    .X(net546));
 sky130_fd_sc_hd__buf_2 fanout547 (.A(net551),
    .X(net547));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout548 (.A(net551),
    .X(net548));
 sky130_fd_sc_hd__buf_2 fanout549 (.A(net551),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_2 fanout550 (.A(net551),
    .X(net550));
 sky130_fd_sc_hd__buf_2 fanout551 (.A(net577),
    .X(net551));
 sky130_fd_sc_hd__buf_2 fanout552 (.A(net554),
    .X(net552));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_2 fanout554 (.A(net559),
    .X(net554));
 sky130_fd_sc_hd__buf_2 fanout555 (.A(net559),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_2 fanout556 (.A(net559),
    .X(net556));
 sky130_fd_sc_hd__buf_2 fanout557 (.A(net559),
    .X(net557));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout558 (.A(net559),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_2 fanout559 (.A(net577),
    .X(net559));
 sky130_fd_sc_hd__buf_2 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__buf_2 fanout561 (.A(net564),
    .X(net561));
 sky130_fd_sc_hd__buf_2 fanout562 (.A(net564),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_2 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_2 fanout564 (.A(net569),
    .X(net564));
 sky130_fd_sc_hd__buf_2 fanout565 (.A(net569),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_2 fanout566 (.A(net569),
    .X(net566));
 sky130_fd_sc_hd__buf_2 fanout567 (.A(net569),
    .X(net567));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_2 fanout569 (.A(net577),
    .X(net569));
 sky130_fd_sc_hd__buf_2 fanout570 (.A(net576),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_2 fanout571 (.A(net576),
    .X(net571));
 sky130_fd_sc_hd__buf_2 fanout572 (.A(net576),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_2 fanout573 (.A(net576),
    .X(net573));
 sky130_fd_sc_hd__buf_2 fanout574 (.A(net576),
    .X(net574));
 sky130_fd_sc_hd__buf_1 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_2 fanout576 (.A(net577),
    .X(net576));
 sky130_fd_sc_hd__clkbuf_4 fanout577 (.A(\fifo_bank_register.clk ),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_4 fanout578 (.A(net580),
    .X(net578));
 sky130_fd_sc_hd__buf_4 fanout579 (.A(net580),
    .X(net579));
 sky130_fd_sc_hd__buf_2 fanout580 (.A(net596),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_4 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__buf_2 fanout582 (.A(net585),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_4 fanout583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_4 fanout584 (.A(net585),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_2 fanout585 (.A(net596),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_4 fanout586 (.A(net588),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_4 fanout587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__buf_2 fanout588 (.A(net595),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_4 fanout589 (.A(net595),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_4 fanout590 (.A(net595),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_4 fanout591 (.A(net595),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_2 fanout592 (.A(net595),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_4 fanout593 (.A(net595),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_2 fanout594 (.A(net595),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_4 fanout595 (.A(net596),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_4 fanout596 (.A(net259),
    .X(net596));
 sky130_fd_sc_hd__buf_2 fanout597 (.A(net602),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_4 fanout598 (.A(net601),
    .X(net598));
 sky130_fd_sc_hd__buf_2 fanout599 (.A(net601),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_4 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_2 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_4 fanout602 (.A(net618),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_4 fanout603 (.A(net607),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_4 fanout604 (.A(net607),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_4 fanout605 (.A(net607),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_4 fanout606 (.A(net607),
    .X(net606));
 sky130_fd_sc_hd__buf_2 fanout607 (.A(net617),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_4 fanout608 (.A(net612),
    .X(net608));
 sky130_fd_sc_hd__buf_2 fanout609 (.A(net612),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_4 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_4 fanout611 (.A(net612),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_2 fanout612 (.A(net617),
    .X(net612));
 sky130_fd_sc_hd__buf_4 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_2 fanout614 (.A(net617),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_4 fanout615 (.A(net617),
    .X(net615));
 sky130_fd_sc_hd__buf_2 fanout616 (.A(net617),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_2 fanout617 (.A(net618),
    .X(net617));
 sky130_fd_sc_hd__buf_2 fanout618 (.A(net259),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_4 fanout619 (.A(net626),
    .X(net619));
 sky130_fd_sc_hd__buf_2 fanout620 (.A(net626),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_4 fanout621 (.A(net626),
    .X(net621));
 sky130_fd_sc_hd__buf_2 fanout622 (.A(net626),
    .X(net622));
 sky130_fd_sc_hd__clkbuf_4 fanout623 (.A(net625),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_4 fanout624 (.A(net626),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_2 fanout625 (.A(net626),
    .X(net625));
 sky130_fd_sc_hd__buf_2 fanout626 (.A(net635),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_4 fanout627 (.A(net634),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_4 fanout628 (.A(net634),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_4 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_4 fanout630 (.A(net634),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_4 fanout631 (.A(net633),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_2 fanout632 (.A(net633),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_4 fanout633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__buf_2 fanout634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_4 fanout635 (.A(net670),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_4 fanout636 (.A(net638),
    .X(net636));
 sky130_fd_sc_hd__buf_2 fanout637 (.A(net638),
    .X(net637));
 sky130_fd_sc_hd__buf_2 fanout638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_2 fanout639 (.A(net640),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_4 fanout640 (.A(net670),
    .X(net640));
 sky130_fd_sc_hd__buf_4 fanout641 (.A(net650),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_4 fanout642 (.A(net650),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_4 fanout643 (.A(net646),
    .X(net643));
 sky130_fd_sc_hd__clkbuf_4 fanout644 (.A(net646),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_2 fanout645 (.A(net646),
    .X(net645));
 sky130_fd_sc_hd__buf_2 fanout646 (.A(net650),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_4 fanout647 (.A(net648),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_4 fanout648 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_4 fanout649 (.A(net650),
    .X(net649));
 sky130_fd_sc_hd__buf_2 fanout650 (.A(net670),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 fanout651 (.A(net652),
    .X(net651));
 sky130_fd_sc_hd__buf_4 fanout652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__buf_4 fanout653 (.A(net660),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_4 fanout654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_4 fanout655 (.A(net657),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_4 fanout656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_2 fanout657 (.A(net660),
    .X(net657));
 sky130_fd_sc_hd__buf_4 fanout658 (.A(net659),
    .X(net658));
 sky130_fd_sc_hd__buf_2 fanout659 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_4 fanout660 (.A(net670),
    .X(net660));
 sky130_fd_sc_hd__clkbuf_4 fanout661 (.A(net663),
    .X(net661));
 sky130_fd_sc_hd__buf_2 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__clkbuf_4 fanout663 (.A(net669),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_4 fanout664 (.A(net667),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_4 fanout665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_4 fanout666 (.A(net667),
    .X(net666));
 sky130_fd_sc_hd__buf_2 fanout667 (.A(net669),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_4 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_4 fanout669 (.A(net670),
    .X(net669));
 sky130_fd_sc_hd__buf_4 fanout670 (.A(net259),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(first_round_reg),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\ks1.key_reg[58] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\mix1.data_reg[73] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\mix1.data_reg[112] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\mix1.data_reg[33] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\mix1.data_reg[93] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\mix1.data_reg[123] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\mix1.data_reg[85] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\mix1.data_reg[117] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\mix1.data_reg[76] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\mix1.data_reg[80] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\mix1.data_reg[118] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\ks1.key_reg[120] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\mix1.data_reg[77] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\mix1.data_reg[104] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\mix1.data_reg[92] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\mix1.data_reg[84] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\mix1.data_reg[101] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\mix1.data_reg[89] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\mix1.data_reg[83] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\mix1.data_reg[109] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\mix1.data_reg[49] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\mix1.data_reg[37] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\ks1.key_reg[123] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\mix1.data_reg[119] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\mix1.data_reg[39] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\mix1.data_reg[86] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\ks1.key_reg[115] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\ks1.key_reg[114] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\ks1.key_reg[27] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\ks1.key_reg[76] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\ks1.key_reg[107] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\mix1.data_reg[58] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\ks1.key_reg[99] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\ks1.key_reg[41] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\ks1.key_reg[85] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\ks1.key_reg[119] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\ks1.key_reg[70] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\ks1.key_reg[84] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\ks1.key_reg[102] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\ks1.key_reg[86] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\ks1.col[0] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\ks1.key_reg[56] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\ks1.key_reg[83] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\ks1.key_reg[55] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\mix1.data_reg[122] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\ks1.key_reg[53] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\ks1.key_reg[48] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\ks1.key_reg[104] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\ks1.key_reg[33] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\ks1.key_reg[113] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\ks1.key_reg[122] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\ks1.key_reg[51] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\ks1.key_reg[78] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\ks1.key_reg[45] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\ks1.key_reg[124] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\ks1.key_reg[79] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\ks1.key_reg[34] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\ks1.key_reg[54] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\ks1.key_reg[88] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\ks1.key_reg[69] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\ks1.key_reg[32] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\ks1.key_reg[36] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\ks1.key_reg[103] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\ks1.key_reg[97] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\ks1.key_reg[98] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\ks1.key_reg[71] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\ks1.key_reg[109] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\ks1.key_reg[47] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\ks1.key_reg[87] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\ks1.key_reg[74] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\ks1.key_reg[50] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\ks1.key_reg[49] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\ks1.key_reg[118] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\ks1.key_reg[67] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\ks1.key_reg[80] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\ks1.key_reg[65] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\mix1.data_reg[68] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\mix1.data_reg[105] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\ks1.key_reg[125] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\ks1.key_reg[46] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\ks1.key_reg[116] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\ks1.key_reg[82] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\ks1.key_reg[91] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\ks1.key_reg[64] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\ks1.key_reg[117] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\ks1.key_reg[68] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\ks1.key_reg[89] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\ks1.key_reg[127] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\mix1.data_reg[116] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\ks1.key_reg[30] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\ks1.key_reg[61] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\ks1.key_reg[59] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\ks1.key_reg[2] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\ks1.key_reg[75] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\mix1.data_reg[34] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\mix1.data_reg[32] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\ks1.key_reg[13] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\mix1.data_reg[115] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\mix1.data_reg[70] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\ks1.key_reg[21] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\ks1.key_reg[14] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\ks1.key_reg[57] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\mix1.data_reg[36] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\ks1.key_reg[16] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\ks1.key_reg[6] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\ks1.key_reg[1] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\ks1.key_reg[0] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\mix1.state[0] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\mix1.data_reg[127] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\ks1.key_reg[11] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\ks1.key_reg[10] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\mix1.data_reg[100] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\ks1.key_reg[63] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\mix1.data_reg[54] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\mix1.data_reg[110] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\ks1.key_reg[25] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\ks1.key_reg[7] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\ks1.key_reg[26] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\mix1.data_reg[57] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\mix1.data_reg[94] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\mix1.data_reg[102] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\mix1.data_reg[45] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\mix1.data_reg[99] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\sub1.state[4] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\mix1.data_reg[71] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\ks1.key_reg[105] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\mix1.data_reg[98] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\mix1.data_reg[43] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\mix1.data_reg[61] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\mix1.data_reg[95] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\mix1.data_reg[40] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\mix1.data_reg[74] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\mix1.data_reg[103] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\mix1.data_reg[125] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\ks1.key_reg[60] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\mix1.data_reg[46] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\mix1.data_reg[79] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\mix1.data_reg[42] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\mix1.data_reg[65] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\mix1.data_reg[55] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\mix1.data_reg[35] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\mix1.data_reg[91] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\mix1.data_reg[78] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\mix1.data_reg[113] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\mix1.data_reg[96] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\ks1.key_reg[40] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\mix1.data_reg[53] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\mix1.data_reg[48] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\mix1.data_reg[60] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\mix1.data_reg[59] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\mix1.data_reg[120] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\mix1.data_reg[111] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\mix1.data_reg[107] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\mix1.data_reg[87] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\mix1.data_reg[82] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\mix1.data_reg[114] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\ks1.key_reg[108] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\mix1.data_reg[69] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\mix1.data_reg[106] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\mix1.data_reg[90] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\mix1.data_reg[50] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\mix1.data_reg[41] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\mix1.data_reg[81] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\mix1.data_reg[56] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\mix1.data_reg[121] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\mix1.data_reg[108] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\mix1.data_reg[97] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\ks1.key_reg[44] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\mix1.data_reg[75] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\mix1.data_reg[88] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\mix1.data_reg[38] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\mix1.data_reg[51] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\mix1.data_reg[52] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\mix1.data_reg[126] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\mix1.data_reg[124] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\mix1.data_reg[44] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\mix1.data_reg[47] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\mix1.data_reg[72] ),
    .X(net769));
 sky130_fd_sc_hd__buf_4 input1 (.A(data_i[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(data_i[108]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input100 (.A(data_i[74]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(data_i[75]),
    .X(net101));
 sky130_fd_sc_hd__buf_2 input102 (.A(data_i[76]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 input103 (.A(data_i[77]),
    .X(net103));
 sky130_fd_sc_hd__buf_4 input104 (.A(data_i[78]),
    .X(net104));
 sky130_fd_sc_hd__buf_2 input105 (.A(data_i[79]),
    .X(net105));
 sky130_fd_sc_hd__buf_4 input106 (.A(data_i[7]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 input107 (.A(data_i[80]),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(data_i[81]),
    .X(net108));
 sky130_fd_sc_hd__buf_4 input109 (.A(data_i[82]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(data_i[109]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input110 (.A(data_i[83]),
    .X(net110));
 sky130_fd_sc_hd__buf_4 input111 (.A(data_i[84]),
    .X(net111));
 sky130_fd_sc_hd__buf_2 input112 (.A(data_i[85]),
    .X(net112));
 sky130_fd_sc_hd__buf_4 input113 (.A(data_i[86]),
    .X(net113));
 sky130_fd_sc_hd__buf_4 input114 (.A(data_i[87]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(data_i[88]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 input116 (.A(data_i[89]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(data_i[8]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 input118 (.A(data_i[90]),
    .X(net118));
 sky130_fd_sc_hd__buf_4 input119 (.A(data_i[91]),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input12 (.A(data_i[10]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input120 (.A(data_i[92]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(data_i[93]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 input122 (.A(data_i[94]),
    .X(net122));
 sky130_fd_sc_hd__buf_2 input123 (.A(data_i[95]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_8 input124 (.A(data_i[96]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_8 input125 (.A(data_i[97]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 input126 (.A(data_i[98]),
    .X(net126));
 sky130_fd_sc_hd__buf_4 input127 (.A(data_i[99]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 input128 (.A(data_i[9]),
    .X(net128));
 sky130_fd_sc_hd__buf_4 input129 (.A(decrypt_i),
    .X(net129));
 sky130_fd_sc_hd__buf_4 input13 (.A(data_i[110]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input130 (.A(key_i[0]),
    .X(net130));
 sky130_fd_sc_hd__buf_4 input131 (.A(key_i[100]),
    .X(net131));
 sky130_fd_sc_hd__buf_4 input132 (.A(key_i[101]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 input133 (.A(key_i[102]),
    .X(net133));
 sky130_fd_sc_hd__buf_4 input134 (.A(key_i[103]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 input135 (.A(key_i[104]),
    .X(net135));
 sky130_fd_sc_hd__buf_4 input136 (.A(key_i[105]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 input137 (.A(key_i[106]),
    .X(net137));
 sky130_fd_sc_hd__buf_4 input138 (.A(key_i[107]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_8 input139 (.A(key_i[108]),
    .X(net139));
 sky130_fd_sc_hd__buf_2 input14 (.A(data_i[111]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 input140 (.A(key_i[109]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 input141 (.A(key_i[10]),
    .X(net141));
 sky130_fd_sc_hd__buf_4 input142 (.A(key_i[110]),
    .X(net142));
 sky130_fd_sc_hd__buf_4 input143 (.A(key_i[111]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 input144 (.A(key_i[112]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 input145 (.A(key_i[113]),
    .X(net145));
 sky130_fd_sc_hd__buf_4 input146 (.A(key_i[114]),
    .X(net146));
 sky130_fd_sc_hd__buf_4 input147 (.A(key_i[115]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 input148 (.A(key_i[116]),
    .X(net148));
 sky130_fd_sc_hd__buf_4 input149 (.A(key_i[117]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(data_i[112]),
    .X(net15));
 sky130_fd_sc_hd__buf_4 input150 (.A(key_i[118]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_8 input151 (.A(key_i[119]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 input152 (.A(key_i[11]),
    .X(net152));
 sky130_fd_sc_hd__buf_4 input153 (.A(key_i[120]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(key_i[121]),
    .X(net154));
 sky130_fd_sc_hd__buf_4 input155 (.A(key_i[122]),
    .X(net155));
 sky130_fd_sc_hd__buf_4 input156 (.A(key_i[123]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(key_i[124]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 input158 (.A(key_i[125]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(key_i[126]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(data_i[113]),
    .X(net16));
 sky130_fd_sc_hd__buf_4 input160 (.A(key_i[127]),
    .X(net160));
 sky130_fd_sc_hd__buf_4 input161 (.A(key_i[12]),
    .X(net161));
 sky130_fd_sc_hd__buf_4 input162 (.A(key_i[13]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 input163 (.A(key_i[14]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 input164 (.A(key_i[15]),
    .X(net164));
 sky130_fd_sc_hd__buf_2 input165 (.A(key_i[16]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_4 input166 (.A(key_i[17]),
    .X(net166));
 sky130_fd_sc_hd__buf_4 input167 (.A(key_i[18]),
    .X(net167));
 sky130_fd_sc_hd__buf_4 input168 (.A(key_i[19]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 input169 (.A(key_i[1]),
    .X(net169));
 sky130_fd_sc_hd__buf_2 input17 (.A(data_i[114]),
    .X(net17));
 sky130_fd_sc_hd__buf_4 input170 (.A(key_i[20]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 input171 (.A(key_i[21]),
    .X(net171));
 sky130_fd_sc_hd__buf_4 input172 (.A(key_i[22]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 input173 (.A(key_i[23]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_8 input174 (.A(key_i[24]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 input175 (.A(key_i[25]),
    .X(net175));
 sky130_fd_sc_hd__buf_4 input176 (.A(key_i[26]),
    .X(net176));
 sky130_fd_sc_hd__buf_4 input177 (.A(key_i[27]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 input178 (.A(key_i[28]),
    .X(net178));
 sky130_fd_sc_hd__buf_4 input179 (.A(key_i[29]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(data_i[115]),
    .X(net18));
 sky130_fd_sc_hd__buf_4 input180 (.A(key_i[2]),
    .X(net180));
 sky130_fd_sc_hd__buf_4 input181 (.A(key_i[30]),
    .X(net181));
 sky130_fd_sc_hd__buf_2 input182 (.A(key_i[31]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 input183 (.A(key_i[32]),
    .X(net183));
 sky130_fd_sc_hd__buf_4 input184 (.A(key_i[33]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_4 input185 (.A(key_i[34]),
    .X(net185));
 sky130_fd_sc_hd__buf_4 input186 (.A(key_i[35]),
    .X(net186));
 sky130_fd_sc_hd__buf_4 input187 (.A(key_i[36]),
    .X(net187));
 sky130_fd_sc_hd__buf_4 input188 (.A(key_i[37]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 input189 (.A(key_i[38]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_8 input19 (.A(data_i[116]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_8 input190 (.A(key_i[39]),
    .X(net190));
 sky130_fd_sc_hd__buf_4 input191 (.A(key_i[3]),
    .X(net191));
 sky130_fd_sc_hd__buf_4 input192 (.A(key_i[40]),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 input193 (.A(key_i[41]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_8 input194 (.A(key_i[42]),
    .X(net194));
 sky130_fd_sc_hd__buf_4 input195 (.A(key_i[43]),
    .X(net195));
 sky130_fd_sc_hd__buf_4 input196 (.A(key_i[44]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_4 input197 (.A(key_i[45]),
    .X(net197));
 sky130_fd_sc_hd__buf_2 input198 (.A(key_i[46]),
    .X(net198));
 sky130_fd_sc_hd__buf_4 input199 (.A(key_i[47]),
    .X(net199));
 sky130_fd_sc_hd__buf_2 input2 (.A(data_i[100]),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input20 (.A(data_i[117]),
    .X(net20));
 sky130_fd_sc_hd__buf_4 input200 (.A(key_i[48]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_8 input201 (.A(key_i[49]),
    .X(net201));
 sky130_fd_sc_hd__buf_4 input202 (.A(key_i[4]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_4 input203 (.A(key_i[50]),
    .X(net203));
 sky130_fd_sc_hd__buf_4 input204 (.A(key_i[51]),
    .X(net204));
 sky130_fd_sc_hd__buf_4 input205 (.A(key_i[52]),
    .X(net205));
 sky130_fd_sc_hd__buf_4 input206 (.A(key_i[53]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 input207 (.A(key_i[54]),
    .X(net207));
 sky130_fd_sc_hd__buf_2 input208 (.A(key_i[55]),
    .X(net208));
 sky130_fd_sc_hd__buf_4 input209 (.A(key_i[56]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_8 input21 (.A(data_i[118]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_8 input210 (.A(key_i[57]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 input211 (.A(key_i[58]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 input212 (.A(key_i[59]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 input213 (.A(key_i[5]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 input214 (.A(key_i[60]),
    .X(net214));
 sky130_fd_sc_hd__buf_4 input215 (.A(key_i[61]),
    .X(net215));
 sky130_fd_sc_hd__buf_4 input216 (.A(key_i[62]),
    .X(net216));
 sky130_fd_sc_hd__buf_4 input217 (.A(key_i[63]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 input218 (.A(key_i[64]),
    .X(net218));
 sky130_fd_sc_hd__buf_2 input219 (.A(key_i[65]),
    .X(net219));
 sky130_fd_sc_hd__buf_4 input22 (.A(data_i[119]),
    .X(net22));
 sky130_fd_sc_hd__buf_4 input220 (.A(key_i[66]),
    .X(net220));
 sky130_fd_sc_hd__buf_4 input221 (.A(key_i[67]),
    .X(net221));
 sky130_fd_sc_hd__buf_4 input222 (.A(key_i[68]),
    .X(net222));
 sky130_fd_sc_hd__buf_4 input223 (.A(key_i[69]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 input224 (.A(key_i[6]),
    .X(net224));
 sky130_fd_sc_hd__buf_4 input225 (.A(key_i[70]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_8 input226 (.A(key_i[71]),
    .X(net226));
 sky130_fd_sc_hd__buf_4 input227 (.A(key_i[72]),
    .X(net227));
 sky130_fd_sc_hd__buf_4 input228 (.A(key_i[73]),
    .X(net228));
 sky130_fd_sc_hd__buf_4 input229 (.A(key_i[74]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(data_i[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input230 (.A(key_i[75]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 input231 (.A(key_i[76]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 input232 (.A(key_i[77]),
    .X(net232));
 sky130_fd_sc_hd__buf_4 input233 (.A(key_i[78]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 input234 (.A(key_i[79]),
    .X(net234));
 sky130_fd_sc_hd__buf_4 input235 (.A(key_i[7]),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_8 input236 (.A(key_i[80]),
    .X(net236));
 sky130_fd_sc_hd__buf_4 input237 (.A(key_i[81]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 input238 (.A(key_i[82]),
    .X(net238));
 sky130_fd_sc_hd__buf_4 input239 (.A(key_i[83]),
    .X(net239));
 sky130_fd_sc_hd__buf_4 input24 (.A(data_i[120]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input240 (.A(key_i[84]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 input241 (.A(key_i[85]),
    .X(net241));
 sky130_fd_sc_hd__buf_4 input242 (.A(key_i[86]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 input243 (.A(key_i[87]),
    .X(net243));
 sky130_fd_sc_hd__buf_4 input244 (.A(key_i[88]),
    .X(net244));
 sky130_fd_sc_hd__buf_4 input245 (.A(key_i[89]),
    .X(net245));
 sky130_fd_sc_hd__buf_4 input246 (.A(key_i[8]),
    .X(net246));
 sky130_fd_sc_hd__buf_4 input247 (.A(key_i[90]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_4 input248 (.A(key_i[91]),
    .X(net248));
 sky130_fd_sc_hd__buf_2 input249 (.A(key_i[92]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(data_i[121]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input250 (.A(key_i[93]),
    .X(net250));
 sky130_fd_sc_hd__buf_4 input251 (.A(key_i[94]),
    .X(net251));
 sky130_fd_sc_hd__buf_2 input252 (.A(key_i[95]),
    .X(net252));
 sky130_fd_sc_hd__buf_4 input253 (.A(key_i[96]),
    .X(net253));
 sky130_fd_sc_hd__buf_4 input254 (.A(key_i[97]),
    .X(net254));
 sky130_fd_sc_hd__buf_4 input255 (.A(key_i[98]),
    .X(net255));
 sky130_fd_sc_hd__buf_4 input256 (.A(key_i[99]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 input257 (.A(key_i[9]),
    .X(net257));
 sky130_fd_sc_hd__buf_6 input258 (.A(load_i),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 input259 (.A(reset),
    .X(net259));
 sky130_fd_sc_hd__buf_2 input26 (.A(data_i[122]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(data_i[123]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(data_i[124]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(data_i[125]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input3 (.A(data_i[101]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input30 (.A(data_i[126]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 input31 (.A(data_i[127]),
    .X(net31));
 sky130_fd_sc_hd__buf_4 input32 (.A(data_i[12]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(data_i[13]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(data_i[14]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(data_i[15]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(data_i[16]),
    .X(net36));
 sky130_fd_sc_hd__buf_4 input37 (.A(data_i[17]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(data_i[18]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(data_i[19]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input4 (.A(data_i[102]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input40 (.A(data_i[1]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_8 input41 (.A(data_i[20]),
    .X(net41));
 sky130_fd_sc_hd__buf_4 input42 (.A(data_i[21]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(data_i[22]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_8 input44 (.A(data_i[23]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(data_i[24]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(data_i[25]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_8 input47 (.A(data_i[26]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(data_i[27]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(data_i[28]),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input5 (.A(data_i[103]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(data_i[29]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 input51 (.A(data_i[2]),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(data_i[30]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(data_i[31]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 input54 (.A(data_i[32]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 input55 (.A(data_i[33]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 input56 (.A(data_i[34]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(data_i[35]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(data_i[36]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_8 input59 (.A(data_i[37]),
    .X(net59));
 sky130_fd_sc_hd__buf_4 input6 (.A(data_i[104]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input60 (.A(data_i[38]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(data_i[39]),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input62 (.A(data_i[3]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(data_i[40]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(data_i[41]),
    .X(net64));
 sky130_fd_sc_hd__buf_4 input65 (.A(data_i[42]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 input66 (.A(data_i[43]),
    .X(net66));
 sky130_fd_sc_hd__buf_4 input67 (.A(data_i[44]),
    .X(net67));
 sky130_fd_sc_hd__buf_4 input68 (.A(data_i[45]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_4 input69 (.A(data_i[46]),
    .X(net69));
 sky130_fd_sc_hd__buf_4 input7 (.A(data_i[105]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input70 (.A(data_i[47]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input71 (.A(data_i[48]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input72 (.A(data_i[49]),
    .X(net72));
 sky130_fd_sc_hd__buf_4 input73 (.A(data_i[4]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 input74 (.A(data_i[50]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 input75 (.A(data_i[51]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 input76 (.A(data_i[52]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 input77 (.A(data_i[53]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input78 (.A(data_i[54]),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(data_i[55]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(data_i[106]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input80 (.A(data_i[56]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(data_i[57]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 input82 (.A(data_i[58]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(data_i[59]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 input84 (.A(data_i[5]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 input85 (.A(data_i[60]),
    .X(net85));
 sky130_fd_sc_hd__buf_4 input86 (.A(data_i[61]),
    .X(net86));
 sky130_fd_sc_hd__buf_4 input87 (.A(data_i[62]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 input88 (.A(data_i[63]),
    .X(net88));
 sky130_fd_sc_hd__buf_4 input89 (.A(data_i[64]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 input9 (.A(data_i[107]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 input90 (.A(data_i[65]),
    .X(net90));
 sky130_fd_sc_hd__buf_4 input91 (.A(data_i[66]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 input92 (.A(data_i[67]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(data_i[68]),
    .X(net93));
 sky130_fd_sc_hd__buf_4 input94 (.A(data_i[69]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(data_i[6]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 input96 (.A(data_i[70]),
    .X(net96));
 sky130_fd_sc_hd__buf_4 input97 (.A(data_i[71]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 input98 (.A(data_i[72]),
    .X(net98));
 sky130_fd_sc_hd__buf_4 input99 (.A(data_i[73]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net260),
    .X(data_o[0]));
 sky130_fd_sc_hd__clkbuf_4 output261 (.A(net261),
    .X(data_o[100]));
 sky130_fd_sc_hd__clkbuf_4 output262 (.A(net262),
    .X(data_o[101]));
 sky130_fd_sc_hd__clkbuf_4 output263 (.A(net263),
    .X(data_o[102]));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net264),
    .X(data_o[103]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(data_o[104]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(data_o[105]));
 sky130_fd_sc_hd__clkbuf_4 output267 (.A(net267),
    .X(data_o[106]));
 sky130_fd_sc_hd__clkbuf_4 output268 (.A(net268),
    .X(data_o[107]));
 sky130_fd_sc_hd__clkbuf_4 output269 (.A(net269),
    .X(data_o[108]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(data_o[109]));
 sky130_fd_sc_hd__clkbuf_4 output271 (.A(net271),
    .X(data_o[10]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(data_o[110]));
 sky130_fd_sc_hd__clkbuf_4 output273 (.A(net273),
    .X(data_o[111]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(data_o[112]));
 sky130_fd_sc_hd__clkbuf_4 output275 (.A(net275),
    .X(data_o[113]));
 sky130_fd_sc_hd__clkbuf_4 output276 (.A(net276),
    .X(data_o[114]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(data_o[115]));
 sky130_fd_sc_hd__clkbuf_4 output278 (.A(net278),
    .X(data_o[116]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(data_o[117]));
 sky130_fd_sc_hd__clkbuf_4 output280 (.A(net280),
    .X(data_o[118]));
 sky130_fd_sc_hd__clkbuf_4 output281 (.A(net281),
    .X(data_o[119]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(data_o[11]));
 sky130_fd_sc_hd__clkbuf_4 output283 (.A(net283),
    .X(data_o[120]));
 sky130_fd_sc_hd__clkbuf_4 output284 (.A(net284),
    .X(data_o[121]));
 sky130_fd_sc_hd__clkbuf_4 output285 (.A(net285),
    .X(data_o[122]));
 sky130_fd_sc_hd__clkbuf_4 output286 (.A(net286),
    .X(data_o[123]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(data_o[124]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(data_o[125]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(data_o[126]));
 sky130_fd_sc_hd__clkbuf_4 output290 (.A(net290),
    .X(data_o[127]));
 sky130_fd_sc_hd__clkbuf_4 output291 (.A(net291),
    .X(data_o[12]));
 sky130_fd_sc_hd__clkbuf_4 output292 (.A(net292),
    .X(data_o[13]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(data_o[14]));
 sky130_fd_sc_hd__clkbuf_4 output294 (.A(net294),
    .X(data_o[15]));
 sky130_fd_sc_hd__clkbuf_4 output295 (.A(net295),
    .X(data_o[16]));
 sky130_fd_sc_hd__clkbuf_4 output296 (.A(net296),
    .X(data_o[17]));
 sky130_fd_sc_hd__clkbuf_4 output297 (.A(net297),
    .X(data_o[18]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(data_o[19]));
 sky130_fd_sc_hd__clkbuf_4 output299 (.A(net299),
    .X(data_o[1]));
 sky130_fd_sc_hd__clkbuf_4 output300 (.A(net300),
    .X(data_o[20]));
 sky130_fd_sc_hd__clkbuf_4 output301 (.A(net301),
    .X(data_o[21]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(data_o[22]));
 sky130_fd_sc_hd__clkbuf_4 output303 (.A(net303),
    .X(data_o[23]));
 sky130_fd_sc_hd__clkbuf_4 output304 (.A(net304),
    .X(data_o[24]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(data_o[25]));
 sky130_fd_sc_hd__clkbuf_4 output306 (.A(net306),
    .X(data_o[26]));
 sky130_fd_sc_hd__clkbuf_4 output307 (.A(net307),
    .X(data_o[27]));
 sky130_fd_sc_hd__clkbuf_4 output308 (.A(net308),
    .X(data_o[28]));
 sky130_fd_sc_hd__clkbuf_4 output309 (.A(net309),
    .X(data_o[29]));
 sky130_fd_sc_hd__clkbuf_4 output310 (.A(net310),
    .X(data_o[2]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net311),
    .X(data_o[30]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .X(data_o[31]));
 sky130_fd_sc_hd__clkbuf_4 output313 (.A(net313),
    .X(data_o[32]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net314),
    .X(data_o[33]));
 sky130_fd_sc_hd__clkbuf_4 output315 (.A(net315),
    .X(data_o[34]));
 sky130_fd_sc_hd__clkbuf_4 output316 (.A(net316),
    .X(data_o[35]));
 sky130_fd_sc_hd__clkbuf_4 output317 (.A(net317),
    .X(data_o[36]));
 sky130_fd_sc_hd__clkbuf_4 output318 (.A(net318),
    .X(data_o[37]));
 sky130_fd_sc_hd__clkbuf_4 output319 (.A(net319),
    .X(data_o[38]));
 sky130_fd_sc_hd__clkbuf_4 output320 (.A(net320),
    .X(data_o[39]));
 sky130_fd_sc_hd__clkbuf_4 output321 (.A(net321),
    .X(data_o[3]));
 sky130_fd_sc_hd__clkbuf_4 output322 (.A(net322),
    .X(data_o[40]));
 sky130_fd_sc_hd__clkbuf_4 output323 (.A(net323),
    .X(data_o[41]));
 sky130_fd_sc_hd__clkbuf_4 output324 (.A(net324),
    .X(data_o[42]));
 sky130_fd_sc_hd__clkbuf_4 output325 (.A(net325),
    .X(data_o[43]));
 sky130_fd_sc_hd__clkbuf_4 output326 (.A(net326),
    .X(data_o[44]));
 sky130_fd_sc_hd__clkbuf_4 output327 (.A(net327),
    .X(data_o[45]));
 sky130_fd_sc_hd__clkbuf_4 output328 (.A(net328),
    .X(data_o[46]));
 sky130_fd_sc_hd__clkbuf_4 output329 (.A(net329),
    .X(data_o[47]));
 sky130_fd_sc_hd__clkbuf_4 output330 (.A(net330),
    .X(data_o[48]));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(data_o[49]));
 sky130_fd_sc_hd__clkbuf_4 output332 (.A(net332),
    .X(data_o[4]));
 sky130_fd_sc_hd__clkbuf_4 output333 (.A(net333),
    .X(data_o[50]));
 sky130_fd_sc_hd__clkbuf_4 output334 (.A(net334),
    .X(data_o[51]));
 sky130_fd_sc_hd__clkbuf_4 output335 (.A(net335),
    .X(data_o[52]));
 sky130_fd_sc_hd__clkbuf_4 output336 (.A(net336),
    .X(data_o[53]));
 sky130_fd_sc_hd__clkbuf_4 output337 (.A(net337),
    .X(data_o[54]));
 sky130_fd_sc_hd__clkbuf_4 output338 (.A(net338),
    .X(data_o[55]));
 sky130_fd_sc_hd__clkbuf_4 output339 (.A(net339),
    .X(data_o[56]));
 sky130_fd_sc_hd__clkbuf_4 output340 (.A(net340),
    .X(data_o[57]));
 sky130_fd_sc_hd__clkbuf_4 output341 (.A(net341),
    .X(data_o[58]));
 sky130_fd_sc_hd__clkbuf_4 output342 (.A(net342),
    .X(data_o[59]));
 sky130_fd_sc_hd__clkbuf_4 output343 (.A(net343),
    .X(data_o[5]));
 sky130_fd_sc_hd__clkbuf_4 output344 (.A(net344),
    .X(data_o[60]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net345),
    .X(data_o[61]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(data_o[62]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .X(data_o[63]));
 sky130_fd_sc_hd__clkbuf_4 output348 (.A(net348),
    .X(data_o[64]));
 sky130_fd_sc_hd__clkbuf_4 output349 (.A(net349),
    .X(data_o[65]));
 sky130_fd_sc_hd__clkbuf_4 output350 (.A(net350),
    .X(data_o[66]));
 sky130_fd_sc_hd__clkbuf_4 output351 (.A(net351),
    .X(data_o[67]));
 sky130_fd_sc_hd__clkbuf_4 output352 (.A(net352),
    .X(data_o[68]));
 sky130_fd_sc_hd__clkbuf_4 output353 (.A(net353),
    .X(data_o[69]));
 sky130_fd_sc_hd__clkbuf_4 output354 (.A(net354),
    .X(data_o[6]));
 sky130_fd_sc_hd__clkbuf_4 output355 (.A(net355),
    .X(data_o[70]));
 sky130_fd_sc_hd__clkbuf_4 output356 (.A(net356),
    .X(data_o[71]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(data_o[72]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(data_o[73]));
 sky130_fd_sc_hd__clkbuf_4 output359 (.A(net359),
    .X(data_o[74]));
 sky130_fd_sc_hd__clkbuf_4 output360 (.A(net360),
    .X(data_o[75]));
 sky130_fd_sc_hd__clkbuf_4 output361 (.A(net361),
    .X(data_o[76]));
 sky130_fd_sc_hd__clkbuf_4 output362 (.A(net362),
    .X(data_o[77]));
 sky130_fd_sc_hd__clkbuf_4 output363 (.A(net363),
    .X(data_o[78]));
 sky130_fd_sc_hd__clkbuf_4 output364 (.A(net364),
    .X(data_o[79]));
 sky130_fd_sc_hd__clkbuf_4 output365 (.A(net365),
    .X(data_o[7]));
 sky130_fd_sc_hd__clkbuf_4 output366 (.A(net366),
    .X(data_o[80]));
 sky130_fd_sc_hd__buf_2 output367 (.A(net367),
    .X(data_o[81]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .X(data_o[82]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(data_o[83]));
 sky130_fd_sc_hd__clkbuf_4 output370 (.A(net370),
    .X(data_o[84]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(data_o[85]));
 sky130_fd_sc_hd__clkbuf_4 output372 (.A(net372),
    .X(data_o[86]));
 sky130_fd_sc_hd__clkbuf_4 output373 (.A(net373),
    .X(data_o[87]));
 sky130_fd_sc_hd__clkbuf_4 output374 (.A(net374),
    .X(data_o[88]));
 sky130_fd_sc_hd__clkbuf_4 output375 (.A(net375),
    .X(data_o[89]));
 sky130_fd_sc_hd__clkbuf_4 output376 (.A(net376),
    .X(data_o[8]));
 sky130_fd_sc_hd__clkbuf_4 output377 (.A(net377),
    .X(data_o[90]));
 sky130_fd_sc_hd__clkbuf_4 output378 (.A(net378),
    .X(data_o[91]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(data_o[92]));
 sky130_fd_sc_hd__clkbuf_4 output380 (.A(net380),
    .X(data_o[93]));
 sky130_fd_sc_hd__clkbuf_4 output381 (.A(net381),
    .X(data_o[94]));
 sky130_fd_sc_hd__clkbuf_4 output382 (.A(net382),
    .X(data_o[95]));
 sky130_fd_sc_hd__clkbuf_4 output383 (.A(net383),
    .X(data_o[96]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .X(data_o[97]));
 sky130_fd_sc_hd__clkbuf_4 output385 (.A(net385),
    .X(data_o[98]));
 sky130_fd_sc_hd__clkbuf_4 output386 (.A(net386),
    .X(data_o[99]));
 sky130_fd_sc_hd__clkbuf_4 output387 (.A(net387),
    .X(data_o[9]));
 sky130_fd_sc_hd__clkbuf_4 output388 (.A(net388),
    .X(ready_o));
endmodule

