* NGSPICE file created from aes_Trojan.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt aes_Trojan clk data_i[0] data_i[100] data_i[101] data_i[102] data_i[103] data_i[104]
+ data_i[105] data_i[106] data_i[107] data_i[108] data_i[109] data_i[10] data_i[110]
+ data_i[111] data_i[112] data_i[113] data_i[114] data_i[115] data_i[116] data_i[117]
+ data_i[118] data_i[119] data_i[11] data_i[120] data_i[121] data_i[122] data_i[123]
+ data_i[124] data_i[125] data_i[126] data_i[127] data_i[12] data_i[13] data_i[14]
+ data_i[15] data_i[16] data_i[17] data_i[18] data_i[19] data_i[1] data_i[20] data_i[21]
+ data_i[22] data_i[23] data_i[24] data_i[25] data_i[26] data_i[27] data_i[28] data_i[29]
+ data_i[2] data_i[30] data_i[31] data_i[32] data_i[33] data_i[34] data_i[35] data_i[36]
+ data_i[37] data_i[38] data_i[39] data_i[3] data_i[40] data_i[41] data_i[42] data_i[43]
+ data_i[44] data_i[45] data_i[46] data_i[47] data_i[48] data_i[49] data_i[4] data_i[50]
+ data_i[51] data_i[52] data_i[53] data_i[54] data_i[55] data_i[56] data_i[57] data_i[58]
+ data_i[59] data_i[5] data_i[60] data_i[61] data_i[62] data_i[63] data_i[64] data_i[65]
+ data_i[66] data_i[67] data_i[68] data_i[69] data_i[6] data_i[70] data_i[71] data_i[72]
+ data_i[73] data_i[74] data_i[75] data_i[76] data_i[77] data_i[78] data_i[79] data_i[7]
+ data_i[80] data_i[81] data_i[82] data_i[83] data_i[84] data_i[85] data_i[86] data_i[87]
+ data_i[88] data_i[89] data_i[8] data_i[90] data_i[91] data_i[92] data_i[93] data_i[94]
+ data_i[95] data_i[96] data_i[97] data_i[98] data_i[99] data_i[9] data_o[0] data_o[100]
+ data_o[101] data_o[102] data_o[103] data_o[104] data_o[105] data_o[106] data_o[107]
+ data_o[108] data_o[109] data_o[10] data_o[110] data_o[111] data_o[112] data_o[113]
+ data_o[114] data_o[115] data_o[116] data_o[117] data_o[118] data_o[119] data_o[11]
+ data_o[120] data_o[121] data_o[122] data_o[123] data_o[124] data_o[125] data_o[126]
+ data_o[127] data_o[12] data_o[13] data_o[14] data_o[15] data_o[16] data_o[17] data_o[18]
+ data_o[19] data_o[1] data_o[20] data_o[21] data_o[22] data_o[23] data_o[24] data_o[25]
+ data_o[26] data_o[27] data_o[28] data_o[29] data_o[2] data_o[30] data_o[31] data_o[32]
+ data_o[33] data_o[34] data_o[35] data_o[36] data_o[37] data_o[38] data_o[39] data_o[3]
+ data_o[40] data_o[41] data_o[42] data_o[43] data_o[44] data_o[45] data_o[46] data_o[47]
+ data_o[48] data_o[49] data_o[4] data_o[50] data_o[51] data_o[52] data_o[53] data_o[54]
+ data_o[55] data_o[56] data_o[57] data_o[58] data_o[59] data_o[5] data_o[60] data_o[61]
+ data_o[62] data_o[63] data_o[64] data_o[65] data_o[66] data_o[67] data_o[68] data_o[69]
+ data_o[6] data_o[70] data_o[71] data_o[72] data_o[73] data_o[74] data_o[75] data_o[76]
+ data_o[77] data_o[78] data_o[79] data_o[7] data_o[80] data_o[81] data_o[82] data_o[83]
+ data_o[84] data_o[85] data_o[86] data_o[87] data_o[88] data_o[89] data_o[8] data_o[90]
+ data_o[91] data_o[92] data_o[93] data_o[94] data_o[95] data_o[96] data_o[97] data_o[98]
+ data_o[99] data_o[9] decrypt_i key_i[0] key_i[100] key_i[101] key_i[102] key_i[103]
+ key_i[104] key_i[105] key_i[106] key_i[107] key_i[108] key_i[109] key_i[10] key_i[110]
+ key_i[111] key_i[112] key_i[113] key_i[114] key_i[115] key_i[116] key_i[117] key_i[118]
+ key_i[119] key_i[11] key_i[120] key_i[121] key_i[122] key_i[123] key_i[124] key_i[125]
+ key_i[126] key_i[127] key_i[12] key_i[13] key_i[14] key_i[15] key_i[16] key_i[17]
+ key_i[18] key_i[19] key_i[1] key_i[20] key_i[21] key_i[22] key_i[23] key_i[24] key_i[25]
+ key_i[26] key_i[27] key_i[28] key_i[29] key_i[2] key_i[30] key_i[31] key_i[32] key_i[33]
+ key_i[34] key_i[35] key_i[36] key_i[37] key_i[38] key_i[39] key_i[3] key_i[40] key_i[41]
+ key_i[42] key_i[43] key_i[44] key_i[45] key_i[46] key_i[47] key_i[48] key_i[49]
+ key_i[4] key_i[50] key_i[51] key_i[52] key_i[53] key_i[54] key_i[55] key_i[56] key_i[57]
+ key_i[58] key_i[59] key_i[5] key_i[60] key_i[61] key_i[62] key_i[63] key_i[64] key_i[65]
+ key_i[66] key_i[67] key_i[68] key_i[69] key_i[6] key_i[70] key_i[71] key_i[72] key_i[73]
+ key_i[74] key_i[75] key_i[76] key_i[77] key_i[78] key_i[79] key_i[7] key_i[80] key_i[81]
+ key_i[82] key_i[83] key_i[84] key_i[85] key_i[86] key_i[87] key_i[88] key_i[89]
+ key_i[8] key_i[90] key_i[91] key_i[92] key_i[93] key_i[94] key_i[95] key_i[96] key_i[97]
+ key_i[98] key_i[99] key_i[9] load_i ready_o reset vccd1 vssd1
XFILLER_0_20_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09671_ _04644_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08622_ ks1.state\[2\] _04370_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08553_ _04595_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_210_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08484_ _04559_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09105_ sbox1.inversion_to_invert_var\[1\] _05105_ vssd1 vssd1 vccd1 vccd1 _05116_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ _05013_ _05057_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_143_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09938_ _05575_ _05777_ _05778_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__a21o_1
XFILLER_0_217_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09869_ _05712_ _05714_ _05715_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11900_ fifo_bank_register.bank\[5\]\[22\] _05317_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07225_ sky130_fd_sc_hd__mux2_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ fifo_bank_register.bank\[2\]\[101\] _05483_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07742_ sky130_fd_sc_hd__mux2_1
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_202 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11831_ _07187_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__clkbuf_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_224 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_235 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_257 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14550_ _02140_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__clkbuf_4
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11762_ _07151_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 addroundkey_data_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13501_ _08077_ vssd1 vssd1 vccd1 vccd1 _08078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10713_ _05602_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__buf_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _02815_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11693_ _07115_ vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__clkbuf_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16220_ _04165_ _04166_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__xor2_2
XFILLER_0_107_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ _05493_ fifo_bank_register.bank\[0\]\[106\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08033_ sky130_fd_sc_hd__mux2_1
X_10644_ _06415_ vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16151_ net208 ks1.key_reg\[55\] _03982_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__mux2_1
X_10575_ sub1.data_o\[82\] _06351_ _06113_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13363_ _05424_ fifo_bank_register.bank\[0\]\[73\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _07997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15102_ _03257_ _03273_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ _05459_ fifo_bank_register.bank\[4\]\[90\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07443_ sky130_fd_sc_hd__mux2_1
X_16082_ ks1.key_reg\[15\] _04041_ _03958_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13294_ _05354_ fifo_bank_register.bank\[0\]\[40\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15033_ _03168_ _03305_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__xnor2_2
X_12245_ _07406_ vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12176_ _07370_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11127_ _06816_ vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__clkbuf_1
X_16984_ net503 _00427_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11058_ _06779_ vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__clkbuf_1
X_15935_ _03907_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__buf_4
XFILLER_0_218_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10009_ _05841_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__xor2_1
XFILLER_0_189_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15866_ net675 _03593_ _03865_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14817_ sub1.data_o\[77\] _03063_ _03092_ sub1.data_o\[45\] vssd1 vssd1 vccd1 vccd1
+ _03093_ sky130_fd_sc_hd__a22o_1
X_17605_ net440 _01048_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18585_ clknet_leaf_81_clk _02014_ net588 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15797_ _03741_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__buf_4
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17536_ net556 _00979_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14748_ ks1.col\[26\] _05559_ _04911_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17467_ net435 _00910_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14679_ fifo_bank_register.bank\[7\]\[125\] _08077_ _08092_ fifo_bank_register.bank\[2\]\[125\]
+ _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16418_ net812 _03978_ _04281_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__mux2_1
X_17398_ net395 _00841_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16349_ net832 _03999_ _04240_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18019_ net482 _01462_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09723_ _05583_ vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__buf_2
XFILLER_0_226_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09654_ fifo_bank_register.bank\[9\]\[125\] _05532_ _05269_ vssd1 vssd1 vccd1 vccd1
+ _05533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08605_ net258 _04468_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__or2_1
XFILLER_0_210_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09585_ _05486_ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08536_ _04586_ vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08467_ _04550_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_1
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08398_ _04514_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10360_ _05609_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09019_ _04713_ _05039_ _05040_ _04716_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10291_ net205 ks1.key_reg\[52\] _06097_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12030_ fifo_bank_register.bank\[5\]\[84\] _05447_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold170 ks1.key_reg\[125\] vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout650 net670 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_2
Xfanout661 net663 vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_4
X_13981_ fifo_bank_register.bank\[0\]\[47\] _02369_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15720_ mix1.data_o\[62\] mix1.data_reg\[62\] _03786_ vssd1 vssd1 vccd1 vccd1 _03790_
+ sky130_fd_sc_hd__mux2_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ _07768_ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__clkbuf_1
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ mix1.data_o\[29\] _03529_ _03753_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__mux2_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12863_ fifo_bank_register.bank\[2\]\[93\] _05466_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07733_ sky130_fd_sc_hd__mux2_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ fifo_bank_register.bank\[0\]\[115\] _02922_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02923_ sky130_fd_sc_hd__mux2_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ clknet_leaf_36_clk _01800_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11814_ fifo_bank_register.bank\[6\]\[110\] _05501_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07179_ sky130_fd_sc_hd__mux2_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _03700_ _03709_ _05228_ _03716_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__a31o_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ fifo_bank_register.bank\[2\]\[60\] _05396_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17321_ net445 _00764_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ fifo_bank_register.bank\[6\]\[108\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[108\]
+ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a22o_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _07142_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ net418 _00695_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_14464_ _02148_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11676_ _07106_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _04112_ _04125_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__xor2_1
XFILLER_0_221_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13415_ _05476_ fifo_bank_register.bank\[0\]\[98\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10627_ sub1.data_o\[86\] _06341_ _06397_ _06399_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06400_ sky130_fd_sc_hd__a221o_1
X_17183_ net548 _00626_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
X_14395_ fifo_bank_register.bank\[9\]\[92\] _02712_ _02736_ _02737_ _02738_ vssd1
+ vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16134_ _04086_ _04087_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__xor2_2
X_13346_ _05407_ fifo_bank_register.bank\[0\]\[65\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07988_ sky130_fd_sc_hd__mux2_1
X_10558_ _06335_ _06336_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16065_ net695 ks1.next_ready_o _04025_ _04026_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__o22a_1
X_13277_ _05338_ fifo_bank_register.bank\[0\]\[32\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07952_ sky130_fd_sc_hd__mux2_1
X_10489_ mix1.data_o\[73\] _06217_ _06241_ _06242_ sub1.data_o\[73\] vssd1 vssd1 vccd1
+ vccd1 _06275_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15016_ _03287_ _03288_ _05198_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__a21oi_1
X_12228_ _07397_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12159_ _05305_ fifo_bank_register.bank\[4\]\[17\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16967_ net492 _00410_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15918_ sub1.data_o\[44\] _03576_ _03892_ sub1.data_o\[108\] vssd1 vssd1 vccd1 vccd1
+ _03897_ sky130_fd_sc_hd__a22o_1
X_16898_ net514 _00341_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15849_ mix1.data_o\[124\] net766 _03729_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__mux2_1
X_18637_ clknet_leaf_21_clk _02066_ net639 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[114\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09370_ fifo_bank_register.bank\[9\]\[33\] _05340_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05341_ sky130_fd_sc_hd__mux2_1
X_18568_ clknet_leaf_63_clk _01997_ net598 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08321_ _04473_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17519_ net398 _00962_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_18499_ clknet_leaf_57_clk _01928_ net618 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ net101 net100 net103 net102 vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__or4_1
XFILLER_0_172_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput264 net264 vssd1 vssd1 vccd1 vccd1 data_o[103] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput275 net275 vssd1 vssd1 vccd1 vccd1 data_o[113] sky130_fd_sc_hd__clkbuf_4
Xoutput286 net286 vssd1 vssd1 vccd1 vccd1 data_o[123] sky130_fd_sc_hd__clkbuf_4
Xoutput297 net297 vssd1 vssd1 vccd1 vccd1 data_o[18] sky130_fd_sc_hd__clkbuf_4
XTAP_5907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09706_ net258 _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09637_ _05521_ vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09568_ fifo_bank_register.bank\[9\]\[97\] _05474_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08519_ _04577_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_2
XFILLER_0_210_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09499_ net230 vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_182_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11530_ fifo_bank_register.bank\[7\]\[104\] _05489_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11461_ fifo_bank_register.bank\[7\]\[71\] _05420_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _06993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13200_ fifo_bank_register.bank\[1\]\[125\] _05532_ _07771_ vssd1 vssd1 vccd1 vccd1
+ _07910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10412_ addroundkey_data_o\[64\] _06206_ _06169_ vssd1 vssd1 vccd1 vccd1 _06207_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11392_ _06956_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__clkbuf_1
X_14180_ fifo_bank_register.bank\[9\]\[69\] _02469_ _02544_ _02545_ _02546_ vssd1
+ vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13131_ _07874_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__clkbuf_1
X_10343_ sub1.data_o\[57\] _06144_ _05991_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10274_ mix1.data_o\[51\] _05952_ _05916_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__o21a_1
X_13062_ fifo_bank_register.bank\[1\]\[59\] _05394_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12013_ fifo_bank_register.bank\[5\]\[76\] _05430_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17870_ net426 _01313_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16821_ clknet_leaf_81_clk _00265_ net586 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[112\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_206_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout480 net481 vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_219_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout491 net498 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_79_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16752_ clknet_leaf_70_clk _00196_ net609 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[43\]
+ sky130_fd_sc_hd__dfrtp_2
X_13964_ fifo_bank_register.bank\[9\]\[45\] _02307_ _02352_ _02353_ _02354_ vssd1
+ vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_191_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15703_ mix1.data_o\[54\] net710 _03775_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__mux2_1
X_12915_ fifo_bank_register.bank\[2\]\[118\] _05518_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16683_ net439 _00131_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13895_ fifo_bank_register.bank\[7\]\[38\] _02218_ _02227_ fifo_bank_register.bank\[2\]\[38\]
+ _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15634_ mix1.data_o\[21\] _03505_ _03742_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__mux2_1
X_18422_ clknet_leaf_83_clk _01852_ net582 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[107\]
+ sky130_fd_sc_hd__dfrtp_2
X_12846_ fifo_bank_register.bank\[2\]\[85\] _05449_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07724_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ clknet_leaf_15_clk _01783_ net629 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[38\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15565_ _03700_ _04935_ _05236_ _03706_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__a31o_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12777_ fifo_bank_register.bank\[2\]\[52\] _05380_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17304_ net539 _00747_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ fifo_bank_register.bank\[6\]\[106\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[106\]
+ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18284_ clknet_leaf_21_clk _01715_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[50\]
+ sky130_fd_sc_hd__dfrtp_4
X_11728_ _07133_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__clkbuf_1
X_15496_ _03652_ _04784_ _05236_ _03661_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17235_ net504 _00678_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _02784_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11659_ _07097_ vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17166_ net554 _00609_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14378_ fifo_bank_register.bank\[9\]\[90\] _02712_ _02717_ _02720_ _02723_ vssd1
+ vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16117_ _04796_ _04072_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13329_ _05390_ fifo_bank_register.bank\[0\]\[57\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07979_ sky130_fd_sc_hd__mux2_1
X_17097_ net473 _00540_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16048_ net139 ks1.key_reg\[108\] _04742_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08870_ addroundkey_data_o\[0\] mix1.data_o\[0\] _04702_ vssd1 vssd1 vccd1 vccd1
+ _04894_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17999_ net440 _01442_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[1\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_58_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09422_ _05312_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ net178 vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08304_ net173 net175 net174 net172 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__or4b_1
XFILLER_0_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09284_ net224 vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08235_ _04388_ _04389_ _04390_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__or4_1
XFILLER_0_160_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08999_ addroundkey_data_o\[50\] mix1.data_o\[50\] _04662_ vssd1 vssd1 vccd1 vccd1
+ _05021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10961_ _06630_ sub1.ready_o sub1.data_o\[119\] _05675_ vssd1 vssd1 vccd1 vccd1 _06701_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12700_ fifo_bank_register.bank\[2\]\[16\] _05303_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13680_ fifo_bank_register.bank\[6\]\[15\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a22o_1
XFILLER_0_195_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10892_ _06638_ vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12631_ _07610_ vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15350_ net798 _03521_ _03560_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ fifo_bank_register.bank\[3\]\[79\] _05436_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ fifo_bank_register.bank\[7\]\[82\] _02623_ _02632_ fifo_bank_register.bank\[2\]\[82\]
+ _02654_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__a221o_1
XFILLER_0_124_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11513_ fifo_bank_register.bank\[7\]\[96\] _05472_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15281_ _03528_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12493_ fifo_bank_register.bank\[3\]\[46\] _05367_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17020_ net556 _00463_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
X_14232_ _02593_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__clkbuf_1
X_11444_ fifo_bank_register.bank\[7\]\[63\] _05403_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14163_ fifo_bank_register.bank\[0\]\[67\] _02531_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11375_ fifo_bank_register.bank\[7\]\[30\] _05333_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13114_ _07865_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__clkbuf_1
X_10326_ mix1.data_o\[55\] _06129_ _06093_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__o21a_1
X_14094_ _02138_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__clkbuf_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ net513 _01365_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_13045_ _07829_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__clkbuf_1
X_10257_ net74 mix1.data_o\[50\] _05934_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__mux2_1
X_10188_ _04609_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__clkbuf_4
X_17853_ net469 _01296_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16804_ clknet_leaf_79_clk _00248_ net578 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[95\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_195_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14996_ addroundkey_data_o\[82\] _03064_ _03084_ addroundkey_data_o\[50\] vssd1 vssd1
+ vccd1 vccd1 _03270_ sky130_fd_sc_hd__a22o_1
X_17784_ net557 _01227_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16735_ clknet_leaf_52_clk _00179_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_13947_ fifo_bank_register.bank\[1\]\[43\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[43\]
+ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16666_ net465 _00114_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13878_ fifo_bank_register.bank\[7\]\[36\] _02218_ _02227_ fifo_bank_register.bank\[2\]\[36\]
+ _02277_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18405_ clknet_leaf_25_clk _01835_ net648 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[90\]
+ sky130_fd_sc_hd__dfrtp_4
X_15617_ _03735_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12829_ fifo_bank_register.bank\[2\]\[77\] _05432_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07715_ sky130_fd_sc_hd__mux2_1
X_16597_ net417 _00045_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18336_ clknet_leaf_37_clk _01766_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15548_ sub1.data_o\[65\] _03691_ _03694_ _03673_ vssd1 vssd1 vccd1 vccd1 _03695_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18267_ clknet_leaf_32_clk _01698_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[33\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ _03651_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ net495 _00661_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18198_ clknet_leaf_25_clk _01629_ net648 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17149_ net574 _00592_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09971_ addroundkey_data_o\[21\] _05808_ _05793_ vssd1 vssd1 vccd1 vccd1 _05809_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08922_ _04706_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08853_ _04649_ _04752_ _04875_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__a22o_4
XFILLER_0_225_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08784_ addroundkey_data_o\[107\] mix1.data_o\[107\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _04808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09405_ _05364_ vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09336_ fifo_bank_register.bank\[9\]\[22\] _05317_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09267_ fifo_bank_register.bank\[9\]\[0\] _05248_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08218_ _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__buf_4
XFILLER_0_16_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09198_ sbox1.alph\[0\] _05119_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11160_ _06833_ vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10111_ _05602_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11091_ _06797_ vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10042_ _05792_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__buf_4
XTAP_5534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold30 mix1.data_reg\[36\] vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold41 mix1.data_reg\[110\] vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14850_ sub1.data_o\[5\] _03100_ _03058_ _03125_ vssd1 vssd1 vccd1 vccd1 _03126_
+ sky130_fd_sc_hd__a211o_1
Xhold52 mix1.data_reg\[98\] vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold63 mix1.data_reg\[65\] vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold74 mix1.data_reg\[120\] vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 mix1.data_reg\[81\] vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold96 mix1.data_reg\[124\] vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13801_ _02208_ fifo_bank_register.data_out\[27\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14781_ _03056_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__buf_6
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11993_ _07273_ vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__clkbuf_1
X_16520_ _04344_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__clkbuf_1
X_13732_ _08106_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__buf_6
X_10944_ net149 ks1.key_reg\[117\] _04639_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16451_ net681 _03914_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13663_ fifo_bank_register.bank\[7\]\[13\] _08182_ _08191_ fifo_bank_register.bank\[2\]\[13\]
+ _02085_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__a221o_1
X_10875_ mix1.data_o\[111\] _06463_ _06575_ _06576_ sub1.data_o\[111\] vssd1 vssd1
+ vccd1 vccd1 _06623_ sky130_fd_sc_hd__a32o_1
XFILLER_0_128_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15402_ _03019_ _03593_ _05219_ _03601_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__a31o_1
XFILLER_0_186_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12614_ _07601_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__clkbuf_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16382_ net848 _04267_ _04264_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__mux2_1
X_13594_ fifo_bank_register.bank\[5\]\[6\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18121_ net428 _01564_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[123\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ mix1.data_reg\[50\] _03493_ _03549_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12545_ _07565_ vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18052_ net555 _01495_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[54\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_227_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15264_ _03515_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12476_ fifo_bank_register.bank\[3\]\[38\] _05350_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07529_ sky130_fd_sc_hd__mux2_1
X_17003_ net414 _00446_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_14215_ _02578_ fifo_bank_register.data_out\[72\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_5 _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ fifo_bank_register.bank\[7\]\[55\] _05386_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15195_ _03264_ _03273_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14146_ fifo_bank_register.bank\[9\]\[65\] _02469_ _02514_ _02515_ _02516_ vssd1
+ vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ fifo_bank_register.bank\[7\]\[22\] _05317_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06939_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10309_ sub1.data_o\[54\] _06112_ _06113_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__mux2_1
X_14077_ fifo_bank_register.bank\[7\]\[58\] _02380_ _02389_ fifo_bank_register.bank\[2\]\[58\]
+ _02454_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11289_ _05520_ fifo_bank_register.bank\[8\]\[119\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17905_ net393 _01348_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_13028_ _07820_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17836_ net465 _01279_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17767_ net423 _01210_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14979_ sub1.data_o\[106\] _03056_ _03252_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16718_ clknet_leaf_43_clk _00162_ net658 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17698_ net410 _01141_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16649_ net547 _00097_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ sbox1.inversion_to_invert_var\[1\] _05105_ sbox1.inversion_to_invert_var\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__or3b_1
XFILLER_0_57_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18319_ clknet_leaf_8_clk _01749_ net633 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09052_ _05068_ _05069_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ addroundkey_data_o\[19\] _05791_ _05793_ vssd1 vssd1 vccd1 vccd1 _05794_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08905_ addroundkey_data_o\[53\] mix1.data_o\[53\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04929_ sky130_fd_sc_hd__mux2_1
X_09885_ _05712_ _05729_ _05730_ _05716_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__a22o_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _04653_ _04834_ _04847_ _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__a211o_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _04776_ _04783_ _04787_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__or4_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ addroundkey_round\[1\] addroundkey_round\[2\] addroundkey_round\[3\] vssd1
+ vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__nor3_1
XFILLER_0_211_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ _06428_ _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09319_ fifo_bank_register.bank\[9\]\[17\] _05305_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10591_ _06076_ _06362_ _06366_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ _05476_ fifo_bank_register.bank\[4\]\[98\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12261_ _05407_ fifo_bank_register.bank\[4\]\[65\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14000_ _02386_ fifo_bank_register.data_out\[49\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11212_ _05443_ fifo_bank_register.bank\[8\]\[82\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06861_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12192_ _05338_ fifo_bank_register.bank\[4\]\[32\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11143_ _06824_ vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__clkbuf_1
XTAP_6021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11074_ _05305_ fifo_bank_register.bank\[8\]\[17\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06788_ sky130_fd_sc_hd__mux2_1
X_15951_ net703 ks1.next_ready_o _03923_ _03924_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__o22a_1
XTAP_6076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput120 data_i[92] vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_4
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput131 key_i[100] vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_4
XTAP_5342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10025_ _05855_ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__xor2_1
X_14902_ addroundkey_data_o\[30\] _04377_ _05606_ _03176_ vssd1 vssd1 vccd1 vccd1
+ _03177_ sky130_fd_sc_hd__a211o_1
Xinput142 key_i[110] vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_4
Xinput153 key_i[120] vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__buf_4
XTAP_5364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15882_ _03873_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__clkbuf_1
XTAP_5375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput164 key_i[15] vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_4
XTAP_5386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput175 key_i[25] vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_204_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput186 key_i[35] vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_4
XFILLER_0_215_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17621_ net534 _01064_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14833_ sub1.data_o\[85\] _03108_ _03066_ sub1.data_o\[53\] vssd1 vssd1 vccd1 vccd1
+ _03109_ sky130_fd_sc_hd__a22o_1
Xinput197 key_i[45] vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_4
XTAP_4674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ net547 _00995_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
X_14764_ ks1.col\[18\] _05559_ _00007_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11976_ _07264_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _04335_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13715_ fifo_bank_register.bank\[1\]\[19\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__a22o_1
X_10927_ sub1.data_o\[116\] _06669_ _05608_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__mux2_1
X_17483_ net476 _00926_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14695_ fifo_bank_register.bank\[7\]\[127\] _08077_ _08092_ fifo_bank_register.bank\[2\]\[127\]
+ _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13646_ fifo_bank_register.bank\[5\]\[11\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__a22o_1
X_16434_ _04297_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__clkbuf_1
X_10858_ mix1.data_o\[109\] _06463_ _06575_ _06576_ sub1.data_o\[109\] vssd1 vssd1
+ vccd1 vccd1 _06608_ sky130_fd_sc_hd__a32o_1
XFILLER_0_6_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _04258_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13577_ _08144_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_229_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10789_ _06395_ _06514_ sub1.data_o\[102\] _06384_ vssd1 vssd1 vccd1 vccd1 _06546_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15316_ _03550_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18104_ net466 _01547_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[106\]
+ sky130_fd_sc_hd__dfxtp_1
X_12528_ _07556_ vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16296_ _03957_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__buf_4
XFILLER_0_26_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15247_ net783 _03502_ _03498_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18035_ net415 _01478_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[37\]
+ sky130_fd_sc_hd__dfxtp_4
X_12459_ _07508_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__buf_4
XFILLER_0_112_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15178_ _03410_ _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__xor2_1
XFILLER_0_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14129_ fifo_bank_register.bank\[1\]\[63\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[63\]
+ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09670_ addroundkey_round\[3\] _05540_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08621_ _04642_ _04644_ ks1.state\[1\] ks1.state\[0\] ks1.state\[2\] vssd1 vssd1
+ vccd1 vccd1 _04645_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17819_ net566 _01262_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08552_ addroundkey_data_o\[114\] fifo_bank_register.data_out\[114\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08483_ addroundkey_data_o\[81\] fifo_bank_register.data_out\[81\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__mux2_2
XFILLER_0_159_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09104_ sbox1.inversion_to_invert_var\[3\] sbox1.inversion_to_invert_var\[0\] vssd1
+ vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09035_ _04966_ _05056_ _04874_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__mux2_4
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09937_ _05201_ _05754_ sub1.data_o\[18\] _05585_ vssd1 vssd1 vccd1 vccd1 _05778_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_99_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09868_ _05567_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__clkbuf_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _04677_ _04841_ _04842_ _04682_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ mix1.data_o\[4\] _05586_ _05618_ _05621_ sub1.data_o\[4\] vssd1 vssd1 vccd1
+ vccd1 _05654_ sky130_fd_sc_hd__a32o_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ fifo_bank_register.bank\[6\]\[118\] _05518_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07187_ sky130_fd_sc_hd__mux2_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_214 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_225 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_258 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11761_ fifo_bank_register.bank\[6\]\[85\] _05449_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07151_ sky130_fd_sc_hd__mux2_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 _05757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _08076_ vssd1 vssd1 vccd1 vccd1 _08077_ sky130_fd_sc_hd__clkbuf_4
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712_ _06475_ vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _02814_ fifo_bank_register.data_out\[101\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11692_ fifo_bank_register.bank\[6\]\[52\] _05380_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _08032_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__clkbuf_1
X_10643_ addroundkey_data_o\[87\] _06414_ _06327_ vssd1 vssd1 vccd1 vccd1 _06415_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16150_ _04100_ _04101_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__xor2_2
X_13362_ _07996_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__clkbuf_1
X_10574_ net109 mix1.data_o\[82\] _06111_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15101_ _03336_ _03371_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_140_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12313_ _07364_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16081_ _05005_ _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_210_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13293_ _07937_ vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__buf_4
XFILLER_0_146_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15032_ _03264_ _03304_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12244_ _05390_ fifo_bank_register.bank\[4\]\[57\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12175_ _05321_ fifo_bank_register.bank\[4\]\[24\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11126_ _05357_ fifo_bank_register.bank\[8\]\[41\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16983_ net497 _00426_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11057_ _05288_ fifo_bank_register.bank\[8\]\[9\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06779_ sky130_fd_sc_hd__mux2_1
X_15934_ _03904_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__xor2_1
XTAP_5161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10008_ net175 ks1.key_reg\[25\] _05825_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__mux2_1
XTAP_5194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15865_ net675 _03593_ _03861_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_204_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17604_ net494 _01047_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
X_14816_ _03091_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__clkbuf_4
X_18584_ clknet_leaf_81_clk _02013_ net578 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[111\]
+ sky130_fd_sc_hd__dfrtp_1
X_15796_ _03829_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__clkbuf_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17535_ net550 _00978_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14747_ _03037_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11959_ fifo_bank_register.bank\[5\]\[50\] _05375_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14678_ fifo_bank_register.bank\[5\]\[125\] _08096_ _08099_ fifo_bank_register.bank\[3\]\[125\]
+ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__a22o_1
X_17466_ net411 _00909_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13629_ _08089_ vssd1 vssd1 vccd1 vccd1 _08190_ sky130_fd_sc_hd__clkbuf_4
X_16417_ _04288_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17397_ net395 _00840_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348_ _04249_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16279_ ks1.next_ready_o _03992_ _04212_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18018_ net516 _01461_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[20\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09722_ _04617_ mix1.ready_o vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__and2_1
XFILLER_0_198_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09653_ net158 vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__clkbuf_4
X_08604_ _04611_ net671 _04619_ _04630_ vssd1 vssd1 vccd1 vccd1 next_addroundkey_start_i
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09584_ fifo_bank_register.bank\[9\]\[102\] _05485_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08535_ addroundkey_data_o\[106\] fifo_bank_register.data_out\[106\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ addroundkey_data_o\[73\] fifo_bank_register.data_out\[73\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__mux2_2
XFILLER_0_33_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08397_ addroundkey_data_o\[40\] fifo_bank_register.data_out\[40\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09018_ addroundkey_data_o\[90\] mix1.data_o\[90\] _04805_ vssd1 vssd1 vccd1 vccd1
+ _05040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10290_ _05707_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold160 ks1.key_reg\[47\] vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold171 ks1.key_reg\[46\] vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout640 net670 vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
Xfanout651 net652 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__clkbuf_4
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__buf_2
X_13980_ fifo_bank_register.bank\[9\]\[47\] _02307_ _02366_ _02367_ _02368_ vssd1
+ vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__a2111o_1
X_12931_ fifo_bank_register.bank\[2\]\[126\] _05534_ _07628_ vssd1 vssd1 vccd1 vccd1
+ _07768_ sky130_fd_sc_hd__mux2_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15650_ _03741_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__buf_4
X_12862_ _07732_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__clkbuf_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11813_ _07078_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__buf_4
X_14601_ fifo_bank_register.bank\[9\]\[115\] _02874_ _02919_ _02920_ _02921_ vssd1
+ vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__a2111o_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15581_ sub1.data_o\[13\] _03660_ _03710_ sub1.data_o\[77\] vssd1 vssd1 vccd1 vccd1
+ _03716_ sky130_fd_sc_hd__a22o_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _07651_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ net445 _00763_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14532_ fifo_bank_register.bank\[7\]\[108\] _02785_ _02794_ fifo_bank_register.bank\[2\]\[108\]
+ _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a221o_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ fifo_bank_register.bank\[6\]\[77\] _05432_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17251_ net499 _00694_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_14463_ _02146_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11675_ fifo_bank_register.bank\[6\]\[44\] _05363_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13414_ _08023_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__clkbuf_1
X_16202_ _03901_ _04149_ _04150_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__o21ai_1
X_10626_ mix1.data_o\[86\] _06129_ _06398_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__o21a_1
X_17182_ net565 _00625_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14394_ fifo_bank_register.bank\[1\]\[92\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[92\]
+ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16133_ net206 ks1.key_reg\[53\] _03910_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13345_ _07987_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10557_ net236 ks1.key_reg\[80\] _06097_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__mux2_8
XFILLER_0_180_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _04959_ _04024_ _04371_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__a21o_1
X_13276_ _07951_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10488_ sub1.data_o\[73\] _06273_ _06239_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__mux2_1
X_15015_ _03152_ _03247_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__xnor2_4
X_12227_ _05373_ fifo_bank_register.bank\[4\]\[49\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ _07360_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11109_ _05340_ fifo_bank_register.bank\[8\]\[33\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06807_ sky130_fd_sc_hd__mux2_1
X_16966_ net475 _00409_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_12089_ fifo_bank_register.bank\[5\]\[112\] _05506_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15917_ _03717_ _04943_ _05196_ _03896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__a31o_1
XFILLER_0_223_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16897_ net572 _00340_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18636_ clknet_leaf_21_clk _02065_ net639 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[113\]
+ sky130_fd_sc_hd__dfrtp_4
X_15848_ _03856_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__clkbuf_1
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18567_ clknet_leaf_66_clk _01996_ net604 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_15779_ mix1.data_o\[90\] net752 _03819_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ addroundkey_data_o\[4\] fifo_bank_register.data_out\[4\] _04468_ vssd1 vssd1
+ vccd1 vccd1 _04473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17518_ net392 _00961_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18498_ clknet_leaf_58_clk _01927_ net602 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08251_ _04404_ _04405_ _04406_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__or4_1
X_17449_ net445 _00892_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput265 net265 vssd1 vssd1 vccd1 vccd1 data_o[104] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput276 net276 vssd1 vssd1 vccd1 vccd1 data_o[114] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput287 net287 vssd1 vssd1 vccd1 vccd1 data_o[124] sky130_fd_sc_hd__buf_2
XFILLER_0_199_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput298 net298 vssd1 vssd1 vccd1 vccd1 data_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_226_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ addroundkey_ready_o _05568_ _04618_ net388 vssd1 vssd1 vccd1 vccd1 _05569_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09636_ fifo_bank_register.bank\[9\]\[119\] _05520_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09567_ net254 vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__buf_2
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08518_ addroundkey_data_o\[98\] fifo_bank_register.data_out\[98\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__mux2_4
X_09498_ _05427_ vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08449_ addroundkey_data_o\[65\] fifo_bank_register.data_out\[65\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__mux2_4
XFILLER_0_135_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11460_ _06992_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10411_ _06204_ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__xor2_1
X_11391_ fifo_bank_register.bank\[7\]\[38\] _05350_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13130_ fifo_bank_register.bank\[1\]\[91\] _05462_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07874_ sky130_fd_sc_hd__mux2_1
X_10342_ net81 mix1.data_o\[57\] _05989_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ _07837_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__clkbuf_1
X_10273_ _05949_ _06078_ _06080_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12012_ _07283_ vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16820_ clknet_leaf_4_clk _00264_ net584 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[111\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_219_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout470 net471 vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_2
Xfanout481 net530 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_2
X_16751_ clknet_leaf_70_clk _00195_ net608 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[42\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout492 net498 vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__buf_2
XFILLER_0_219_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13963_ fifo_bank_register.bank\[1\]\[45\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[45\]
+ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_221_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15702_ _03780_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__clkbuf_1
X_12914_ _07759_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__clkbuf_1
X_13894_ fifo_bank_register.bank\[5\]\[38\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[38\]
+ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a22o_1
X_16682_ net493 _00130_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18421_ clknet_leaf_84_clk _01851_ net582 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[106\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15633_ _03744_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__clkbuf_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ _07723_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ clknet_leaf_15_clk _01782_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ sub1.data_o\[70\] _03691_ _03705_ _03594_ vssd1 vssd1 vccd1 vccd1 _03706_
+ sky130_fd_sc_hd__a22o_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _07687_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ net540 _00746_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ fifo_bank_register.bank\[6\]\[69\] _05415_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07133_ sky130_fd_sc_hd__mux2_1
X_14515_ fifo_bank_register.bank\[7\]\[106\] _02785_ _02794_ fifo_bank_register.bank\[2\]\[106\]
+ _02844_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__a221o_1
X_18283_ clknet_leaf_22_clk _01714_ net643 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[49\]
+ sky130_fd_sc_hd__dfrtp_4
X_15495_ sub1.data_o\[110\] _03660_ _03653_ sub1.data_o\[46\] vssd1 vssd1 vccd1 vccd1
+ _03661_ sky130_fd_sc_hd__a22o_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234_ net500 _00677_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11658_ fifo_bank_register.bank\[6\]\[36\] _05346_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07097_ sky130_fd_sc_hd__mux2_1
X_14446_ _02783_ fifo_bank_register.data_out\[98\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10609_ sub1.data_o\[85\] _06382_ _06113_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14377_ fifo_bank_register.bank\[1\]\[90\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[90\]
+ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a22o_1
X_17165_ net527 _00608_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
X_11589_ _07060_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13328_ _07978_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16116_ _04070_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__xor2_2
X_17096_ net474 _00539_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13259_ _07942_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__clkbuf_1
X_16047_ net707 _03901_ _04009_ _04010_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_161_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17998_ net421 _01441_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16949_ net411 _00392_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_76_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09421_ net203 vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__buf_2
X_18619_ clknet_leaf_15_clk _02048_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[112\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09352_ _05328_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08303_ net177 net176 net179 net178 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_158_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09283_ _05281_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ net127 net126 net3 net2 vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__or4_2
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ _04661_ _05018_ _05019_ _04668_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_227_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_67_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10960_ sub1.data_o\[119\] _06699_ _05608_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _05509_ vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10891_ addroundkey_data_o\[112\] _06637_ _06612_ vssd1 vssd1 vccd1 vccd1 _06638_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12630_ fifo_bank_register.bank\[3\]\[111\] _05504_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12561_ _07573_ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ _07019_ vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__clkbuf_1
X_14300_ fifo_bank_register.bank\[5\]\[82\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[82\]
+ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__a22o_1
X_15280_ net782 _03527_ _03498_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__mux2_1
X_12492_ _07537_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _02592_ fifo_bank_register.data_out\[74\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02593_ sky130_fd_sc_hd__mux2_1
X_11443_ _06983_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14162_ fifo_bank_register.bank\[9\]\[67\] _02469_ _02528_ _02529_ _02530_ vssd1
+ vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_81_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11374_ _06935_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13113_ fifo_bank_register.bank\[1\]\[83\] _05445_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07865_ sky130_fd_sc_hd__mux2_1
X_10325_ _04626_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14093_ _02136_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ fifo_bank_register.bank\[1\]\[50\] _05375_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07829_ sky130_fd_sc_hd__mux2_1
X_17921_ net573 _01364_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_10256_ _06065_ vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17852_ net470 _01295_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
X_10187_ mix1.data_o\[42\] _05876_ _05993_ _05994_ sub1.data_o\[42\] vssd1 vssd1 vccd1
+ vccd1 _06004_ sky130_fd_sc_hd__a32o_1
XFILLER_0_205_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16803_ clknet_leaf_73_clk _00247_ net593 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[94\]
+ sky130_fd_sc_hd__dfrtp_2
X_17783_ net407 _01226_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14995_ sub1.data_o\[114\] _03079_ _03268_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_58_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16734_ clknet_leaf_50_clk _00178_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_13946_ fifo_bank_register.bank\[6\]\[43\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[43\]
+ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16665_ net468 _00113_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13877_ fifo_bank_register.bank\[5\]\[36\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[36\]
+ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18404_ clknet_leaf_25_clk _01834_ net648 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[89\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15616_ mix1.data_o\[13\] _03467_ _03730_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12828_ _07714_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__clkbuf_1
X_16596_ net423 _00044_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18335_ clknet_leaf_37_clk _01765_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_15547_ sub1.data_o\[97\] sub1.data_o\[33\] _03671_ vssd1 vssd1 vccd1 vccd1 _03694_
+ sky130_fd_sc_hd__mux2_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12759_ _07678_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18266_ clknet_leaf_34_clk _01697_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[32\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15478_ sub1.data_o\[39\] _03650_ _03636_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17217_ net439 _00660_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14429_ _02768_ fifo_bank_register.data_out\[96\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02769_ sky130_fd_sc_hd__mux2_1
X_18197_ clknet_leaf_25_clk _01628_ net648 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17148_ net556 _00591_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09970_ _05806_ _05807_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__xor2_1
X_17079_ net428 _00522_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
X_08921_ mix1.data_o\[101\] _04900_ _04943_ _04944_ vssd1 vssd1 vccd1 vccd1 _04945_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ _04794_ _04873_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_209_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08783_ _04668_ _04804_ _04806_ _04716_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_49_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ fifo_bank_register.bank\[9\]\[44\] _05363_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ net172 vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__buf_2
XFILLER_0_118_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09266_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08217_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09197_ sbox1.alph\[1\] _05111_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10110_ _05933_ vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11090_ _05321_ fifo_bank_register.bank\[8\]\[24\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10041_ _05869_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__xor2_1
XTAP_5524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold20 ks1.key_reg\[59\] vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold31 ks1.key_reg\[16\] vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold42 ks1.key_reg\[25\] vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold53 mix1.data_reg\[43\] vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold64 mix1.data_reg\[55\] vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold75 mix1.data_reg\[111\] vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 mix1.data_reg\[56\] vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13800_ _08068_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__buf_4
Xhold97 mix1.data_reg\[44\] vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14780_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__clkbuf_8
X_11992_ fifo_bank_register.bank\[5\]\[66\] _05409_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07273_ sky130_fd_sc_hd__mux2_1
XTAP_4889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10943_ _05623_ _06680_ _06684_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__o21ai_4
X_13731_ _02146_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16450_ _04305_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10874_ sub1.data_o\[111\] _06621_ _06573_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13662_ fifo_bank_register.bank\[5\]\[13\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ sub1.data_o\[76\] _03600_ _03595_ sub1.data_o\[12\] vssd1 vssd1 vccd1 vccd1
+ _03601_ sky130_fd_sc_hd__a22o_1
X_12613_ fifo_bank_register.bank\[3\]\[103\] _05487_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _08158_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16381_ _04132_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__inv_2
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ net428 _01563_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15332_ _03558_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12544_ fifo_bank_register.bank\[3\]\[70\] _05417_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07565_ sky130_fd_sc_hd__mux2_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18051_ net568 _01494_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[53\]
+ sky130_fd_sc_hd__dfxtp_2
X_15263_ net761 _03514_ _03498_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__mux2_1
X_12475_ _07528_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17002_ net422 _00445_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14214_ fifo_bank_register.bank\[0\]\[72\] _02577_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02578_ sky130_fd_sc_hd__mux2_1
X_11426_ _06974_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__clkbuf_1
X_15194_ _03457_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _02208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14145_ fifo_bank_register.bank\[1\]\[65\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[65\]
+ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__a22o_1
X_11357_ _06938_ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _05608_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__buf_4
X_14076_ fifo_bank_register.bank\[5\]\[58\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[58\]
+ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
X_11288_ _06900_ vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13027_ fifo_bank_register.bank\[1\]\[42\] _05359_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07820_ sky130_fd_sc_hd__mux2_1
X_17904_ net399 _01347_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_10239_ sub1.data_o\[48\] _05971_ _06048_ _06049_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _06050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_219_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17835_ net450 _01278_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17766_ net417 _01209_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14978_ sub1.data_o\[10\] _04377_ _03081_ _03251_ vssd1 vssd1 vccd1 vccd1 _03252_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16717_ clknet_leaf_51_clk _00161_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13929_ fifo_bank_register.bank\[7\]\[41\] _02299_ _02308_ fifo_bank_register.bank\[2\]\[41\]
+ _02323_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17697_ net401 _01140_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16648_ net565 _00096_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16579_ net505 _00027_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_09120_ _05113_ _05114_ _05117_ _05129_ _05130_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_57_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18318_ clknet_leaf_8_clk _01748_ net632 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09051_ _05016_ sbox1.ah\[2\] vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18249_ clknet_leaf_1_clk _01680_ net623 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_199_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09953_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08904_ _04879_ _04925_ _04926_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__a22o_1
X_09884_ mix1.data_o\[13\] _05677_ _05703_ _05704_ sub1.data_o\[13\] vssd1 vssd1 vccd1
+ vccd1 _05730_ sky130_fd_sc_hd__a32o_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08835_ _04850_ _04852_ _04855_ _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__or4_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08766_ _04710_ _04788_ _04684_ _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__a22o_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ ks1.state\[1\] ks1.state\[0\] _04720_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__nand3_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09318_ net166 vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10590_ sub1.data_o\[83\] _06341_ _06364_ _06365_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06366_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09249_ fifo_bank_register.write_ptr\[0\] fifo_bank_register.write_ptr\[1\] vssd1
+ vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12260_ _07414_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11211_ _06860_ vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__clkbuf_1
X_12191_ _07378_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11142_ _05373_ fifo_bank_register.bank\[8\]\[49\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11073_ _06787_ vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__clkbuf_1
X_15950_ _04759_ _03922_ _04373_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__o21ai_1
XTAP_5321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput110 data_i[83] vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput121 data_i[93] vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
XTAP_6088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14901_ addroundkey_data_o\[94\] _03063_ _03092_ addroundkey_data_o\[62\] vssd1 vssd1
+ vccd1 vccd1 _03176_ sky130_fd_sc_hd__a22o_1
Xinput132 key_i[101] vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__buf_4
X_10024_ net177 ks1.key_reg\[27\] _05825_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__mux2_1
XTAP_6099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput143 key_i[111] vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_4
Xinput154 key_i[121] vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__clkbuf_4
XTAP_5365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15881_ sub1.data_o\[95\] _05244_ _04888_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput165 key_i[16] vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__buf_2
XFILLER_0_76_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput176 key_i[26] vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__buf_4
X_17620_ net506 _01063_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14832_ _03061_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__buf_4
Xinput187 key_i[36] vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__buf_4
XFILLER_0_204_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput198 key_i[46] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XFILLER_0_208_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17551_ net543 _00994_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14763_ _03045_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11975_ fifo_bank_register.bank\[5\]\[58\] _05392_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07264_ sky130_fd_sc_hd__mux2_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ net758 _03456_ _04332_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13714_ fifo_bank_register.bank\[6\]\[19\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10926_ net19 mix1.data_o\[116\] _05602_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__mux2_1
X_17482_ net474 _00925_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14694_ fifo_bank_register.bank\[5\]\[127\] _08096_ _08099_ fifo_bank_register.bank\[3\]\[127\]
+ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_224_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16433_ ks1.key_reg\[111\] _04038_ _04295_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10857_ sub1.data_o\[109\] _06606_ _06573_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__mux2_1
X_13645_ _02070_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ ks1.key_reg\[81\] _04054_ _04252_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__mux2_1
X_10788_ sub1.data_o\[102\] _06544_ _06478_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__mux2_1
X_13576_ _08143_ fifo_bank_register.data_out\[3\] _08064_ vssd1 vssd1 vccd1 vccd1
+ _08144_ sky130_fd_sc_hd__mux2_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18103_ net468 _01546_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15315_ net754 _03424_ _03549_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12527_ fifo_bank_register.bank\[3\]\[62\] _05401_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16295_ _04221_ vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18034_ net425 _01477_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_15246_ _03385_ _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_169_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12458_ _07519_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11409_ _06965_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__clkbuf_1
X_15177_ _03257_ _03304_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12389_ _07481_ vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14128_ fifo_bank_register.bank\[6\]\[63\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[63\]
+ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14059_ fifo_bank_register.bank\[5\]\[56\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[56\]
+ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_207_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08620_ _04643_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__clkbuf_4
X_17818_ net547 _01261_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08551_ _04594_ vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_1
X_17749_ net517 _01192_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08482_ _04558_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09103_ sbox1.inversion_to_invert_var\[1\] sbox1.inversion_to_invert_var\[2\] vssd1
+ vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09034_ _04752_ _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09936_ sub1.data_o\[18\] _05776_ _05751_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09867_ mix1.data_o\[11\] _05677_ _05703_ _05704_ sub1.data_o\[11\] vssd1 vssd1 vccd1
+ vccd1 _05715_ sky130_fd_sc_hd__a32o_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ addroundkey_data_o\[118\] mix1.data_o\[118\] _04665_ vssd1 vssd1 vccd1 vccd1
+ _04842_ sky130_fd_sc_hd__mux2_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09798_ sub1.data_o\[4\] _05652_ _05610_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__mux2_1
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_204 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08749_ addroundkey_data_o\[17\] mix1.data_o\[17\] _04655_ vssd1 vssd1 vccd1 vccd1
+ _04773_ sky130_fd_sc_hd__mux2_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 net186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_226 net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_237 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _07150_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_248 net251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_259 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ addroundkey_data_o\[95\] _06474_ _06431_ vssd1 vssd1 vccd1 vccd1 _06475_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _07114_ vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10642_ _06412_ _06413_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13430_ _05491_ fifo_bank_register.bank\[0\]\[105\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13361_ _05422_ fifo_bank_register.bank\[0\]\[72\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _07996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10573_ _06350_ vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15100_ _03367_ _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nor2_8
X_12312_ _07441_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13292_ _07959_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__clkbuf_1
X_16080_ _04035_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15031_ _03300_ _03303_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nor2_8
X_12243_ _07405_ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12174_ _07369_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ _06815_ vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16982_ net496 _00425_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11056_ _06778_ vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__clkbuf_1
X_15933_ net218 ks1.key_reg\[64\] _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__mux2_1
XTAP_5151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10007_ _05829_ _05839_ _05840_ _05833_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a22o_1
XTAP_5184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15864_ _03864_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__clkbuf_1
XTAP_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17603_ net490 _01046_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14815_ _03065_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__buf_4
XTAP_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18583_ clknet_leaf_78_clk _02012_ net580 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15795_ mix1.data_o\[98\] net722 _03819_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__mux2_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17534_ net570 _00977_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ ks1.col\[25\] _05553_ _04911_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11958_ _07221_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__buf_4
XFILLER_0_171_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10909_ sub1.data_o\[114\] _06513_ _06652_ _06653_ _04610_ vssd1 vssd1 vccd1 vccd1
+ _06654_ sky130_fd_sc_hd__a221o_1
X_17465_ net470 _00908_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14677_ _02988_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11889_ _07218_ vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__clkbuf_1
X_16416_ net826 _03969_ _04281_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13628_ _08189_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17396_ net390 _00839_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16347_ ks1.key_reg\[73\] _03990_ _04240_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13559_ fifo_bank_register.bank\[0\]\[1\] _08128_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16278_ net683 _04373_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18017_ net502 _01460_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_15229_ _03488_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09721_ _04619_ _05580_ _05581_ _05582_ vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09652_ _05531_ vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08603_ _04623_ _04628_ _04629_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09583_ net133 vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__buf_2
XFILLER_0_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08534_ _04585_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_4
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08465_ _04549_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_1
XFILLER_0_147_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08396_ _04513_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09017_ addroundkey_data_o\[66\] mix1.data_o\[66\] _04665_ vssd1 vssd1 vccd1 vccd1
+ _05039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold150 ks1.key_reg\[34\] vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold161 ks1.key_reg\[87\] vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 ks1.key_reg\[116\] vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout630 net634 vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_4
Xfanout641 net650 vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_4
Xfanout652 net653 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__buf_4
X_09919_ _05707_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__buf_4
Xfanout663 net669 vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12930_ _07767_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__clkbuf_1
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12861_ fifo_bank_register.bank\[2\]\[92\] _05464_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07732_ sky130_fd_sc_hd__mux2_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ fifo_bank_register.bank\[1\]\[115\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[115\]
+ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__a22o_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _07177_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__clkbuf_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15580_ _03700_ _03709_ _05219_ _03715_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__a31o_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _07695_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__clkbuf_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ fifo_bank_register.bank\[5\]\[108\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[108\]
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a22o_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11743_ _07141_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__clkbuf_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17250_ net488 _00693_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14462_ fifo_bank_register.bank\[7\]\[100\] _02785_ _02794_ fifo_bank_register.bank\[2\]\[100\]
+ _02797_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11674_ _07105_ vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16201_ net714 _04136_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__nand2_1
X_13413_ _05474_ fifo_bank_register.bank\[0\]\[97\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08023_ sky130_fd_sc_hd__mux2_1
X_10625_ _05757_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17181_ net560 _00624_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14393_ fifo_bank_register.bank\[6\]\[92\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[92\]
+ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16132_ _04084_ _04085_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__xor2_2
X_10556_ _06076_ _06330_ _06334_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__o21ai_1
X_13344_ _05405_ fifo_bank_register.bank\[0\]\[64\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16063_ _04959_ _04024_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__nor2_1
X_10487_ net99 mix1.data_o\[73\] _06237_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ _05336_ fifo_bank_register.bank\[0\]\[31\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07951_ sky130_fd_sc_hd__mux2_1
X_15014_ _03141_ _03286_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_161_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12226_ _07396_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12157_ _05303_ fifo_bank_register.bank\[4\]\[16\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11108_ _06806_ vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12088_ _07323_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__clkbuf_1
X_16965_ net471 _00408_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15916_ sub1.data_o\[43\] _03576_ _03892_ sub1.data_o\[107\] vssd1 vssd1 vccd1 vccd1
+ _03896_ sky130_fd_sc_hd__a22o_1
X_11039_ _05248_ fifo_bank_register.bank\[8\]\[0\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06770_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16896_ net558 _00339_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18635_ clknet_leaf_21_clk _02064_ net639 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[112\]
+ sky130_fd_sc_hd__dfrtp_4
X_15847_ mix1.data_o\[123\] net774 _03729_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18566_ clknet_leaf_62_clk _01995_ net598 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[93\]
+ sky130_fd_sc_hd__dfrtp_1
X_15778_ _03820_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__clkbuf_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17517_ net414 _00960_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14729_ _03028_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__clkbuf_1
X_18497_ clknet_leaf_59_clk _01926_ net606 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08250_ net92 net91 net94 net93 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17448_ net447 _00891_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ net500 _00822_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput266 net266 vssd1 vssd1 vccd1 vccd1 data_o[105] sky130_fd_sc_hd__buf_2
XFILLER_0_26_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput277 net277 vssd1 vssd1 vccd1 vccd1 data_o[115] sky130_fd_sc_hd__buf_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput288 net288 vssd1 vssd1 vccd1 vccd1 data_o[125] sky130_fd_sc_hd__buf_2
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput299 net299 vssd1 vssd1 vccd1 vccd1 data_o[1] sky130_fd_sc_hd__clkbuf_4
XTAP_5909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09704_ _05567_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09635_ net151 vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09566_ _05473_ vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08517_ _04576_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09497_ fifo_bank_register.bank\[9\]\[74\] _05426_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08448_ _04540_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__buf_1
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _04504_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10410_ net218 ks1.key_reg\[64\] _06166_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ _06955_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10341_ _06143_ vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ fifo_bank_register.bank\[1\]\[58\] _05392_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07837_ sky130_fd_sc_hd__mux2_1
X_10272_ _05913_ _05972_ sub1.data_o\[51\] _06079_ vssd1 vssd1 vccd1 vccd1 _06080_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12011_ fifo_bank_register.bank\[5\]\[75\] _05428_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout460 net461 vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_205_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16750_ clknet_leaf_70_clk _00194_ net609 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[41\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout482 net484 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__buf_2
X_13962_ fifo_bank_register.bank\[6\]\[45\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[45\]
+ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__a22o_1
Xfanout493 net498 vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_219_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15701_ mix1.data_o\[53\] net740 _03775_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__mux2_1
X_12913_ fifo_bank_register.bank\[2\]\[117\] _05516_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16681_ net490 _00129_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13893_ _02291_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18420_ clknet_leaf_11_clk _01850_ net622 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[105\]
+ sky130_fd_sc_hd__dfrtp_4
X_15632_ mix1.data_o\[20\] _03502_ _03742_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12844_ fifo_bank_register.bank\[2\]\[84\] _05447_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07723_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18351_ clknet_leaf_15_clk _01781_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[36\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ sub1.data_o\[102\] sub1.data_o\[38\] _03574_ vssd1 vssd1 vccd1 vccd1 _03705_
+ sky130_fd_sc_hd__mux2_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12775_ fifo_bank_register.bank\[2\]\[51\] _05378_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07687_ sky130_fd_sc_hd__mux2_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17302_ net541 _00745_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ fifo_bank_register.bank\[5\]\[106\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[106\]
+ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__a22o_1
X_18282_ clknet_leaf_22_clk _01713_ net643 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[48\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _07132_ vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__clkbuf_1
X_15494_ _04369_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17233_ net504 _00676_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_14445_ fifo_bank_register.bank\[0\]\[98\] _02782_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02783_ sky130_fd_sc_hd__mux2_1
X_11657_ _07096_ vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__clkbuf_1
X_10608_ net112 mix1.data_o\[85\] _06111_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17164_ net518 _00607_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14376_ _02153_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__clkbuf_4
X_11588_ fifo_bank_register.bank\[6\]\[3\] _05276_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07060_ sky130_fd_sc_hd__mux2_1
X_16115_ net204 ks1.key_reg\[51\] _03937_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__mux2_1
X_13327_ _05388_ fifo_bank_register.bank\[0\]\[56\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10539_ sub1.data_o\[79\] _06317_ _06318_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17095_ net490 _00538_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16046_ _04798_ _04008_ _03914_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__a21oi_1
X_13258_ _05319_ fifo_bank_register.bank\[0\]\[23\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12209_ _05354_ fifo_bank_register.bank\[4\]\[40\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _07904_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17997_ net434 _01440_ net596 vssd1 vssd1 vccd1 vccd1 fifo_bank_register.write_ptr\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_208_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16948_ net432 _00391_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16879_ net398 _00322_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09420_ _05374_ vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18618_ clknet_leaf_0_clk _02047_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[111\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09351_ fifo_bank_register.bank\[9\]\[27\] _05327_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18549_ clknet_leaf_78_clk _01978_ net579 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[76\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08302_ _04455_ _04456_ _04457_ _04458_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09282_ fifo_bank_register.bank\[9\]\[5\] _05280_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08233_ net123 net122 net125 net124 vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__or4_1
XFILLER_0_144_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08997_ addroundkey_data_o\[74\] mix1.data_o\[74\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _05019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09618_ fifo_bank_register.bank\[9\]\[113\] _05508_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10890_ _06635_ _06636_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_211_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09549_ net248 vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__buf_2
XFILLER_0_183_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ fifo_bank_register.bank\[3\]\[78\] _05434_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11511_ fifo_bank_register.bank\[7\]\[95\] _05470_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12491_ fifo_bank_register.bank\[3\]\[45\] _05365_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14230_ fifo_bank_register.bank\[0\]\[74\] _02591_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02592_ sky130_fd_sc_hd__mux2_1
X_11442_ fifo_bank_register.bank\[7\]\[62\] _05401_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14161_ fifo_bank_register.bank\[1\]\[67\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[67\]
+ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a22o_1
X_11373_ _06946_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__clkbuf_1
X_10324_ _06126_ _06125_ _06127_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13112_ _07864_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14092_ _02468_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10255_ addroundkey_data_o\[49\] _06063_ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_
+ sky130_fd_sc_hd__mux2_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ net557 _01363_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_13043_ _07794_ vssd1 vssd1 vccd1 vccd1 _07828_ sky130_fd_sc_hd__buf_4
XFILLER_0_219_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17851_ net433 _01294_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
X_10186_ sub1.data_o\[42\] _06002_ _05991_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16802_ clknet_leaf_79_clk _00246_ net579 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[93\]
+ sky130_fd_sc_hd__dfrtp_4
X_17782_ net393 _01225_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14994_ sub1.data_o\[18\] _03208_ _03059_ _03267_ vssd1 vssd1 vccd1 vccd1 _03268_
+ sky130_fd_sc_hd__a211o_1
X_16733_ clknet_leaf_51_clk _00177_ net616 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_13945_ fifo_bank_register.bank\[7\]\[43\] _02299_ _02308_ fifo_bank_register.bank\[2\]\[43\]
+ _02337_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__a221o_1
XFILLER_0_205_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16664_ net463 _00112_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13876_ _02276_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18403_ clknet_leaf_25_clk _01833_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[88\]
+ sky130_fd_sc_hd__dfrtp_4
X_15615_ _03734_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12827_ fifo_bank_register.bank\[2\]\[76\] _05430_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07714_ sky130_fd_sc_hd__mux2_1
X_16595_ net428 _00043_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18334_ clknet_leaf_35_clk _01764_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_173_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15546_ _03668_ _04935_ _05548_ _03693_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__a31o_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12758_ fifo_bank_register.bank\[2\]\[43\] _05361_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18265_ clknet_leaf_43_clk _01696_ net655 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11709_ fifo_bank_register.bank\[6\]\[60\] _05396_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15477_ sub1.data_o\[71\] _05244_ _03633_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12689_ _07641_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17216_ net490 _00659_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14428_ fifo_bank_register.bank\[0\]\[96\] _02767_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18196_ clknet_leaf_25_clk _01627_ net648 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ net567 _00590_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14359_ fifo_bank_register.bank\[7\]\[89\] _02704_ _02632_ fifo_bank_register.bank\[2\]\[89\]
+ _02705_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17078_ net432 _00521_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08920_ addroundkey_data_o\[101\] _04657_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__or2_1
X_16029_ _03994_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08851_ _04794_ _04873_ _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08782_ addroundkey_data_o\[91\] mix1.data_o\[91\] _04805_ vssd1 vssd1 vccd1 vccd1
+ _04806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09403_ net196 vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__buf_2
XFILLER_0_172_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09334_ _05316_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09265_ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__buf_4
XFILLER_0_209_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08216_ mix1.state\[0\] mix1.state\[1\] vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09196_ sbox1.alph\[3\] _05134_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__nand2_2
XFILLER_0_105_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10040_ net179 ks1.key_reg\[29\] _05825_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__mux2_2
XTAP_5514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold10 ks1.key_reg\[58\] vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold21 ks1.key_reg\[2\] vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold32 ks1.key_reg\[6\] vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold43 ks1.key_reg\[7\] vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold54 mix1.data_reg\[61\] vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold65 mix1.data_reg\[35\] vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold76 mix1.data_reg\[107\] vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 mix1.data_reg\[121\] vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold98 mix1.data_reg\[47\] vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _07272_ vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ _08103_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__buf_6
XFILLER_0_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10942_ sub1.data_o\[117\] _05613_ _06682_ _06683_ _04610_ vssd1 vssd1 vccd1 vccd1
+ _06684_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ _02084_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10873_ net14 mix1.data_o\[111\] _06571_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15400_ _04369_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12612_ _07600_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16380_ _04266_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13592_ _08157_ fifo_bank_register.data_out\[5\] _08064_ vssd1 vssd1 vccd1 vccd1
+ _08158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15331_ mix1.data_reg\[49\] _03491_ _03549_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__mux2_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _07508_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18050_ net567 _01493_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[52\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15262_ _03407_ _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12474_ fifo_bank_register.bank\[3\]\[37\] _05348_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17001_ net416 _00444_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14213_ fifo_bank_register.bank\[9\]\[72\] _02550_ _02574_ _02575_ _02576_ vssd1
+ vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_152_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11425_ fifo_bank_register.bank\[7\]\[54\] _05384_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06974_ sky130_fd_sc_hd__mux2_1
X_15193_ net777 _03456_ _03425_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 _03143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14144_ fifo_bank_register.bank\[6\]\[65\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[65\]
+ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__a22o_1
X_11356_ fifo_bank_register.bank\[7\]\[21\] _05315_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10307_ net78 mix1.data_o\[54\] _06111_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14075_ _02453_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11287_ _05518_ fifo_bank_register.bank\[8\]\[118\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06900_ sky130_fd_sc_hd__mux2_1
X_13026_ _07819_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__clkbuf_1
X_17903_ net398 _01346_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10238_ mix1.data_o\[48\] _05952_ _05916_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10169_ addroundkey_data_o\[40\] _05987_ _05980_ vssd1 vssd1 vccd1 vccd1 _05988_
+ sky130_fd_sc_hd__mux2_1
X_17834_ net452 _01277_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14977_ sub1.data_o\[74\] _03209_ _03067_ sub1.data_o\[42\] vssd1 vssd1 vccd1 vccd1
+ _03251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17765_ net437 _01208_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16716_ clknet_leaf_49_clk _00160_ net616 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13928_ fifo_bank_register.bank\[5\]\[41\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[41\]
+ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17696_ net409 _01139_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16647_ net561 _00095_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
X_13859_ _02261_ fifo_bank_register.data_out\[33\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16578_ net533 _00026_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18317_ clknet_leaf_9_clk _01747_ net633 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_15529_ sub1.data_o\[57\] _05553_ _04884_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09050_ _05016_ sbox1.ah\[2\] vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18248_ clknet_leaf_10_clk _01679_ net623 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18179_ clknet_leaf_12_clk _01610_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09952_ _04640_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__buf_4
XFILLER_0_102_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08903_ _04668_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09883_ sub1.data_o\[13\] _05728_ _05701_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__mux2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _04713_ _04856_ _04857_ _04716_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__a22o_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ addroundkey_data_o\[57\] mix1.data_o\[57\] _04778_ vssd1 vssd1 vccd1 vccd1
+ _04789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ ks1.state\[2\] vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09317_ _05304_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09248_ _05249_ _05250_ fifo_bank_register.write_ptr\[2\] vssd1 vssd1 vccd1 vccd1
+ _05252_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09179_ sbox1.alph\[3\] _05127_ _05188_ _05189_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__o211a_1
XFILLER_0_181_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11210_ _05441_ fifo_bank_register.bank\[8\]\[81\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12190_ _05336_ fifo_bank_register.bank\[4\]\[31\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ _06823_ vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__clkbuf_1
XTAP_6001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11072_ _05303_ fifo_bank_register.bank\[8\]\[16\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06787_ sky130_fd_sc_hd__mux2_1
XTAP_6045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput100 data_i[74] vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_4
XTAP_6067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput111 data_i[84] vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_4
Xinput122 data_i[94] vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_4
XTAP_6078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10023_ _05829_ _05853_ _05854_ _05833_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__a22o_1
X_14900_ sub1.data_o\[126\] _03078_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__a21oi_2
XTAP_5344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput133 key_i[102] vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
XTAP_6089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15880_ _03872_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__clkbuf_1
XTAP_5355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput144 key_i[112] vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_204_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput155 key_i[122] vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_4
XTAP_5377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput166 key_i[17] vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_4
Xinput177 key_i[27] vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_4
XFILLER_0_208_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14831_ _03103_ _03106_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__nor2_8
XTAP_4654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput188 key_i[37] vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_4
Xinput199 key_i[47] vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_4
XFILLER_0_204_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ net544 _00993_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ ks1.col\[17\] _05553_ _00007_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11974_ _07263_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16501_ _04334_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__clkbuf_1
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ fifo_bank_register.bank\[7\]\[19\] _02128_ _08191_ fifo_bank_register.bank\[2\]\[19\]
+ _02129_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10925_ _06668_ vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__clkbuf_1
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17481_ net475 _00924_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14693_ _03002_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16432_ _04296_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__clkbuf_1
X_13644_ _02069_ fifo_bank_register.data_out\[10\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _02070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10856_ net11 mix1.data_o\[109\] _06571_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _04257_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__clkbuf_1
X_13575_ fifo_bank_register.bank\[0\]\[3\] _08142_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08143_ sky130_fd_sc_hd__mux2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10787_ net4 mix1.data_o\[102\] _06476_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18102_ net466 _01545_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[104\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_82_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _03145_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__buf_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _07555_ vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16294_ net811 _04048_ _04206_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18033_ net429 _01476_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[35\]
+ sky130_fd_sc_hd__dfxtp_4
X_15245_ _03372_ _03500_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__xnor2_2
X_12457_ fifo_bank_register.bank\[3\]\[29\] _05331_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11408_ fifo_bank_register.bank\[7\]\[46\] _05367_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15176_ _03415_ _03439_ _03440_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__o21ai_4
X_12388_ _05534_ fifo_bank_register.bank\[4\]\[126\] _07341_ vssd1 vssd1 vccd1 vccd1
+ _07481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14127_ fifo_bank_register.bank\[7\]\[63\] _02461_ _02470_ fifo_bank_register.bank\[2\]\[63\]
+ _02499_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11339_ _06928_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ _02438_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__clkbuf_1
X_13009_ _07810_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17817_ net561 _01260_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08550_ addroundkey_data_o\[113\] fifo_bank_register.data_out\[113\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__mux2_2
X_17748_ net534 _01191_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08481_ addroundkey_data_o\[80\] fifo_bank_register.data_out\[80\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__mux2_2
XFILLER_0_134_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17679_ net543 _01122_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09102_ sbox1.inversion_to_invert_var\[3\] vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09033_ _05009_ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09935_ net38 mix1.data_o\[18\] _05749_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09866_ sub1.data_o\[11\] _05713_ _05701_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__mux2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08817_ addroundkey_data_o\[86\] mix1.data_o\[86\] _04662_ vssd1 vssd1 vccd1 vccd1
+ _04841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09797_ net73 mix1.data_o\[4\] _05604_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__mux2_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _04677_ _04770_ _04706_ _04771_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__a22o_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_205 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_216 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_169_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_217_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08679_ addroundkey_data_o\[100\] _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__or2_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_249 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _06472_ _06473_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__xor2_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ fifo_bank_register.bank\[6\]\[51\] _05378_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07114_ sky130_fd_sc_hd__mux2_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ net243 ks1.key_reg\[87\] _06402_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__mux2_8
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ _07995_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__clkbuf_1
X_10572_ addroundkey_data_o\[81\] _06349_ _06327_ vssd1 vssd1 vccd1 vccd1 _06350_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12311_ _05457_ fifo_bank_register.bank\[4\]\[89\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13291_ _05352_ fifo_bank_register.bank\[0\]\[39\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15030_ addroundkey_data_o\[98\] _03077_ _03302_ vssd1 vssd1 vccd1 vccd1 _03303_
+ sky130_fd_sc_hd__a21oi_4
X_12242_ _05388_ fifo_bank_register.bank\[4\]\[56\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12173_ _05319_ fifo_bank_register.bank\[4\]\[23\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07369_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ _05354_ fifo_bank_register.bank\[8\]\[40\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06815_ sky130_fd_sc_hd__mux2_1
X_16981_ net505 _00424_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11055_ _05286_ fifo_bank_register.bank\[8\]\[8\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06778_ sky130_fd_sc_hd__mux2_1
X_15932_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__buf_4
XTAP_5141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10006_ mix1.data_o\[25\] _05797_ _05821_ _05822_ sub1.data_o\[25\] vssd1 vssd1 vccd1
+ vccd1 _05840_ sky130_fd_sc_hd__a32o_1
XTAP_5174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15863_ _03709_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__or2_1
XTAP_5185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14814_ _03076_ _03089_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__xnor2_4
XTAP_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17602_ net494 _01045_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15794_ _03828_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18582_ clknet_leaf_65_clk _02011_ net590 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _03036_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__clkbuf_1
X_17533_ net570 _00976_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _07254_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ mix1.data_o\[114\] _06494_ _05617_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__o21a_1
X_17464_ net456 _00907_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14676_ _02987_ fifo_bank_register.data_out\[124\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _02988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ fifo_bank_register.bank\[5\]\[17\] _05305_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16415_ _04287_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13627_ _08188_ fifo_bank_register.data_out\[9\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _08189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17395_ net406 _00838_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_10839_ _06591_ vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16346_ _04248_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__clkbuf_1
X_13558_ fifo_bank_register.bank\[9\]\[1\] _08090_ _08125_ _08126_ _08127_ vssd1 vssd1
+ vccd1 vccd1 _08128_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_229_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12509_ _07546_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16277_ _03901_ _03984_ _04211_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13489_ _08065_ _08066_ vssd1 vssd1 vccd1 vccd1 _08067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15228_ net778 _03487_ _03425_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__mux2_1
X_18016_ net533 _01459_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[18\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_160_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15159_ net770 _03424_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09720_ round\[1\] net258 vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__or2_1
X_09651_ fifo_bank_register.bank\[9\]\[124\] _05530_ _05269_ vssd1 vssd1 vccd1 vccd1
+ _05531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08602_ sub1.ready_o _04622_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__and2_2
XFILLER_0_175_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09582_ _05484_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08533_ addroundkey_data_o\[105\] fifo_bank_register.data_out\[105\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08464_ addroundkey_data_o\[72\] fifo_bank_register.data_out\[72\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08395_ addroundkey_data_o\[39\] fifo_bank_register.data_out\[39\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09016_ _04706_ _05036_ _05037_ _04710_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold140 ks1.key_reg\[53\] vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_143_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold151 ks1.key_reg\[54\] vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold162 ks1.key_reg\[74\] vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_218_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold173 ks1.key_reg\[82\] vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_218_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout620 net626 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
XFILLER_0_217_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout631 net633 vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__clkbuf_4
X_09918_ _05568_ _05752_ _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__o21ai_1
Xfanout642 net650 vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__clkbuf_4
Xfanout653 net660 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout664 net667 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
X_09849_ _05698_ vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _07731_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__clkbuf_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ fifo_bank_register.bank\[6\]\[109\] _05499_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07177_ sky130_fd_sc_hd__mux2_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ fifo_bank_register.bank\[2\]\[59\] _05394_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07695_ sky130_fd_sc_hd__mux2_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _02858_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__clkbuf_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ fifo_bank_register.bank\[6\]\[76\] _05430_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07141_ sky130_fd_sc_hd__mux2_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ fifo_bank_register.bank\[5\]\[100\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[100\]
+ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11673_ fifo_bank_register.bank\[6\]\[43\] _05361_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07105_ sky130_fd_sc_hd__mux2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16200_ _05046_ _04148_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13412_ _08022_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__clkbuf_1
X_10624_ _06126_ _06394_ _06396_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__a21o_1
X_17180_ net561 _00623_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14392_ fifo_bank_register.bank\[7\]\[92\] _02704_ _02713_ fifo_bank_register.bank\[2\]\[92\]
+ _02735_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__a221o_1
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16131_ net241 ks1.key_reg\[85\] _03918_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13343_ _07986_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10555_ sub1.data_o\[80\] _05971_ _06332_ _06333_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06334_ sky130_fd_sc_hd__a221o_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16062_ _04019_ _04023_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__xnor2_2
X_13274_ _07950_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10486_ _06272_ vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__clkbuf_1
X_15013_ _03218_ _03285_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__xnor2_1
X_12225_ _05371_ fifo_bank_register.bank\[4\]\[48\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12156_ _07359_ vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11107_ _05338_ fifo_bank_register.bank\[8\]\[32\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12087_ fifo_bank_register.bank\[5\]\[111\] _05504_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07323_ sky130_fd_sc_hd__mux2_1
X_16964_ net531 _00407_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
X_15915_ _03717_ _04943_ _05560_ _03895_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a31o_1
X_11038_ _06768_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16895_ net550 _00338_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_18634_ clknet_leaf_0_clk _02063_ net620 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[127\]
+ sky130_fd_sc_hd__dfrtp_1
X_15846_ _03855_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18565_ clknet_leaf_63_clk _01994_ net598 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[92\]
+ sky130_fd_sc_hd__dfrtp_1
X_15777_ mix1.data_o\[89\] net785 _03819_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ fifo_bank_register.bank\[1\]\[24\] _05321_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07800_ sky130_fd_sc_hd__mux2_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17516_ net416 _00959_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14728_ net806 _05547_ _04916_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18496_ clknet_leaf_58_clk _01925_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14659_ fifo_bank_register.bank\[0\]\[122\] _02972_ _08120_ vssd1 vssd1 vccd1 vccd1
+ _02973_ sky130_fd_sc_hd__mux2_1
X_17447_ net454 _00890_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17378_ net485 _00821_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16329_ _04239_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput267 net267 vssd1 vssd1 vccd1 vccd1 data_o[106] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput278 net278 vssd1 vssd1 vccd1 vccd1 data_o[116] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput289 net289 vssd1 vssd1 vccd1 vccd1 data_o[126] sky130_fd_sc_hd__buf_2
XFILLER_0_199_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09703_ _04609_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__buf_4
XFILLER_0_226_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09634_ _05519_ vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09565_ fifo_bank_register.bank\[9\]\[96\] _05472_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08516_ addroundkey_data_o\[97\] fifo_bank_register.data_out\[97\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ net229 vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__buf_2
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08447_ addroundkey_data_o\[64\] fifo_bank_register.data_out\[64\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__mux2_2
XFILLER_0_93_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08378_ addroundkey_data_o\[31\] fifo_bank_register.data_out\[31\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__mux2_2
XFILLER_0_191_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10340_ addroundkey_data_o\[56\] _06142_ _06064_ vssd1 vssd1 vccd1 vccd1 _06143_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10271_ _05584_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12010_ _07282_ vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout450 net451 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__buf_2
Xfanout461 net472 vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_217_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout472 fifo_bank_register.clk vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__buf_2
X_13961_ fifo_bank_register.bank\[7\]\[45\] _02299_ _02308_ fifo_bank_register.bank\[2\]\[45\]
+ _02351_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__a221o_1
XFILLER_0_205_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout483 net484 vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__buf_2
Xfanout494 net498 vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__buf_2
X_15700_ _03779_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__clkbuf_1
X_12912_ _07758_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__clkbuf_1
X_16680_ net441 _00128_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
X_13892_ _02289_ fifo_bank_register.data_out\[37\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_216_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15631_ _03743_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__clkbuf_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ _07722_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__clkbuf_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18350_ clknet_leaf_18_clk _01780_ net637 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[35\]
+ sky130_fd_sc_hd__dfrtp_4
X_15562_ _03700_ _04935_ _05228_ _03704_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _07686_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ net543 _00744_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
X_14513_ _02843_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ fifo_bank_register.bank\[6\]\[68\] _05413_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18281_ clknet_leaf_3_clk _01712_ net624 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[47\]
+ sky130_fd_sc_hd__dfrtp_4
X_15493_ _03652_ _04784_ _05228_ _03659_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17232_ net493 _00675_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14444_ fifo_bank_register.bank\[9\]\[98\] _02712_ _02779_ _02780_ _02781_ vssd1
+ vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_154_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11656_ fifo_bank_register.bank\[6\]\[35\] _05344_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _05567_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__buf_8
X_17163_ net514 _00606_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
X_14375_ _02151_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11587_ _07059_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16114_ _04068_ _04069_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__xor2_4
X_13326_ _07977_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ _05751_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__clkbuf_4
X_17094_ net481 _00537_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16045_ _04798_ _04008_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__or2_1
X_13257_ _07941_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10469_ addroundkey_data_o\[70\] _06257_ _06248_ vssd1 vssd1 vccd1 vccd1 _06258_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12208_ _07364_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13188_ fifo_bank_register.bank\[1\]\[119\] _05520_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12139_ _07350_ vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17996_ net442 _01439_ net596 vssd1 vssd1 vccd1 vccd1 fifo_bank_register.write_ptr\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16947_ net459 _00390_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_193_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16878_ net393 _00321_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18617_ clknet_leaf_83_clk _02046_ net583 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[110\]
+ sky130_fd_sc_hd__dfrtp_1
X_15829_ mix1.data_o\[114\] net749 _03841_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09350_ net177 vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18548_ clknet_leaf_64_clk _01977_ net599 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08301_ net203 net205 net206 net204 vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_34_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09281_ net213 vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__buf_2
XFILLER_0_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18479_ clknet_leaf_55_clk _01908_ net615 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08232_ net114 net113 net116 net115 vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ addroundkey_data_o\[18\] mix1.data_o\[18\] _04665_ vssd1 vssd1 vccd1 vccd1
+ _05018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09617_ net145 vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__buf_2
XFILLER_0_211_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09548_ _05461_ vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09479_ _05414_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11510_ _07018_ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12490_ _07536_ vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11441_ _06982_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14160_ fifo_bank_register.bank\[6\]\[67\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[67\]
+ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ fifo_bank_register.bank\[7\]\[29\] _05331_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13111_ fifo_bank_register.bank\[1\]\[82\] _05443_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07864_ sky130_fd_sc_hd__mux2_1
X_10323_ _06090_ _05972_ sub1.data_o\[55\] _06079_ vssd1 vssd1 vccd1 vccd1 _06127_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14091_ _02467_ fifo_bank_register.data_out\[59\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02468_ sky130_fd_sc_hd__mux2_1
X_13042_ _07827_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__clkbuf_1
X_10254_ _05792_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_219_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17850_ net456 _01293_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10185_ net65 mix1.data_o\[42\] _05989_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16801_ clknet_leaf_69_clk _00245_ net593 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[92\]
+ sky130_fd_sc_hd__dfrtp_2
X_17781_ net393 _01224_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14993_ sub1.data_o\[82\] _03064_ _03084_ sub1.data_o\[50\] vssd1 vssd1 vccd1 vccd1
+ _03267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16732_ clknet_leaf_43_clk _00176_ net658 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_13944_ fifo_bank_register.bank\[5\]\[43\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[43\]
+ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13875_ _02275_ fifo_bank_register.data_out\[35\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16663_ net458 _00111_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18402_ clknet_leaf_25_clk _01832_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_15614_ mix1.data_o\[12\] _03456_ _03730_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__mux2_1
X_12826_ _07713_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16594_ net430 _00042_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18333_ clknet_leaf_16_clk _01763_ net630 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15545_ sub1.data_o\[64\] _03691_ _03692_ _03673_ vssd1 vssd1 vccd1 vccd1 _03693_
+ sky130_fd_sc_hd__a22o_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _07677_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11708_ _07078_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__buf_4
X_15476_ _03649_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__clkbuf_1
X_18264_ clknet_leaf_52_clk _01695_ net655 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ fifo_bank_register.bank\[2\]\[10\] _05290_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17215_ net440 _00658_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14427_ fifo_bank_register.bank\[9\]\[96\] _02712_ _02764_ _02765_ _02766_ vssd1
+ vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_181_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11639_ fifo_bank_register.bank\[6\]\[27\] _05327_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07087_ sky130_fd_sc_hd__mux2_1
X_18195_ clknet_leaf_25_clk _01626_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17146_ net567 _00589_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14358_ fifo_bank_register.bank\[5\]\[89\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[89\]
+ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13309_ _07968_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17077_ net412 _00520_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
X_14289_ fifo_bank_register.bank\[0\]\[80\] _02643_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16028_ ks1.key_reg\[9\] _03993_ _03958_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08850_ _04624_ _04648_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__and2_2
XFILLER_0_23_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08781_ _04655_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__buf_4
XFILLER_0_137_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17979_ net435 _01422_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09402_ _05362_ vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09333_ fifo_bank_register.bank\[9\]\[21\] _05315_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09264_ fifo_bank_register.write_ptr\[2\] fifo_bank_register.write_ptr\[3\] _05266_
+ _05267_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__and4b_1
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08215_ _04373_ vssd1 vssd1 vccd1 vccd1 ks1.next_ready_o sky130_fd_sc_hd__buf_4
XFILLER_0_111_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ _05104_ _04946_ _05196_ _05205_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold11 ks1.key_reg\[120\] vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_220_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold22 ks1.key_reg\[75\] vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold33 ks1.key_reg\[1\] vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold44 ks1.key_reg\[26\] vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _05000_ _04741_ _04750_ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a2bb2o_1
XTAP_4825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold55 mix1.data_reg\[95\] vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold66 mix1.data_reg\[91\] vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold77 mix1.data_reg\[87\] vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold88 mix1.data_reg\[108\] vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ fifo_bank_register.bank\[5\]\[65\] _05407_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold99 mix1.data_reg\[72\] vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10941_ mix1.data_o\[117\] _04626_ _05617_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__o21a_1
XFILLER_0_168_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13660_ _02083_ fifo_bank_register.data_out\[12\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _02084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ _06620_ vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12611_ fifo_bank_register.bank\[3\]\[102\] _05485_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13591_ fifo_bank_register.bank\[0\]\[5\] _08156_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _03557_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _07563_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15261_ _03076_ _03512_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12473_ _07527_ vssd1 vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17000_ net417 _00443_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_14212_ fifo_bank_register.bank\[1\]\[72\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[72\]
+ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11424_ _06973_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__clkbuf_1
X_15192_ _03452_ _03455_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__xor2_4
XFILLER_0_151_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_8 _03143_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14143_ fifo_bank_register.bank\[7\]\[65\] _02461_ _02470_ fifo_bank_register.bank\[2\]\[65\]
+ _02513_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a221o_1
X_11355_ _06937_ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10306_ _05602_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14074_ _02451_ fifo_bank_register.data_out\[57\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11286_ _06899_ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17902_ net395 _01345_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13025_ fifo_bank_register.bank\[1\]\[41\] _05357_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07819_ sky130_fd_sc_hd__mux2_1
X_10237_ _05949_ _06046_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17833_ net448 _01276_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
X_10168_ _05985_ _05986_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__xor2_1
XFILLER_0_174_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17764_ net437 _01207_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1092 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14976_ _03198_ _03248_ _03249_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__a21oi_2
X_10099_ _05923_ vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16715_ clknet_leaf_51_clk _00159_ net651 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_13927_ _02322_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17695_ net536 _01138_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16646_ net560 _00094_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13858_ fifo_bank_register.bank\[0\]\[33\] _02260_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ _07704_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16577_ net532 _00025_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
X_13789_ fifo_bank_register.bank\[1\]\[26\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18316_ clknet_leaf_17_clk _01746_ net633 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15528_ _03683_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18247_ clknet_leaf_2_clk _01678_ net625 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_170_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15459_ sub1.data_o\[65\] _05553_ _03633_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18178_ clknet_leaf_12_clk _01609_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[72\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17129_ net429 _00572_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09951_ _05789_ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08902_ addroundkey_data_o\[77\] mix1.data_o\[77\] _04657_ vssd1 vssd1 vccd1 vccd1
+ _04926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09882_ net33 mix1.data_o\[13\] _05699_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__mux2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08833_ addroundkey_data_o\[94\] mix1.data_o\[94\] _04805_ vssd1 vssd1 vccd1 vccd1
+ _04857_ sky130_fd_sc_hd__mux2_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08764_ addroundkey_data_o\[9\] mix1.data_o\[9\] _04656_ vssd1 vssd1 vccd1 vccd1
+ _04788_ sky130_fd_sc_hd__mux2_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _04653_ _04659_ _04691_ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__a211o_1
XFILLER_0_178_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09316_ fifo_bank_register.bank\[9\]\[16\] _05303_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09247_ _05249_ _05250_ fifo_bank_register.write_ptr\[2\] vssd1 vssd1 vccd1 vccd1
+ _05251_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09178_ sbox1.alph\[3\] _05155_ _05177_ sbox1.alph\[0\] vssd1 vssd1 vccd1 vccd1 _05189_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_17_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11140_ _05371_ fifo_bank_register.bank\[8\]\[48\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11071_ _06786_ vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__clkbuf_1
XTAP_6046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput101 data_i[75] vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_2
XTAP_6057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput112 data_i[85] vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_2
X_10022_ mix1.data_o\[27\] _05797_ _05821_ _05822_ sub1.data_o\[27\] vssd1 vssd1 vccd1
+ vccd1 _05854_ sky130_fd_sc_hd__a32o_1
XTAP_6079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput123 data_i[95] vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_2
XTAP_5345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput134 key_i[103] vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_4
XTAP_5356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput145 key_i[113] vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_216_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput156 key_i[123] vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__buf_4
XFILLER_0_204_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14830_ addroundkey_data_o\[102\] _03077_ _03105_ vssd1 vssd1 vccd1 vccd1 _03106_
+ sky130_fd_sc_hd__a21oi_4
Xinput167 key_i[18] vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_4
XTAP_5389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput178 key_i[28] vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput189 key_i[38] vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_4
XTAP_4666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14761_ _03044_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__clkbuf_1
X_11973_ fifo_bank_register.bank\[5\]\[57\] _05390_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ net746 _03446_ _04332_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10924_ addroundkey_data_o\[115\] _06667_ _06612_ vssd1 vssd1 vccd1 vccd1 _06668_
+ sky130_fd_sc_hd__mux2_1
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ fifo_bank_register.bank\[5\]\[19\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[19\]
+ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17480_ net476 _00923_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_14692_ _03001_ fifo_bank_register.data_out\[126\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _03002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_224_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16431_ ks1.key_reg\[110\] _04028_ _04295_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13643_ fifo_bank_register.bank\[0\]\[10\] _02067_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02069_ sky130_fd_sc_hd__mux2_1
X_10855_ _06605_ vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ fifo_bank_register.bank\[9\]\[3\] _08090_ _08139_ _08140_ _08141_ vssd1 vssd1
+ vccd1 vccd1 _08142_ sky130_fd_sc_hd__a2111o_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ net837 _04046_ _04252_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__mux2_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _06543_ vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__clkbuf_1
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18101_ net459 _01544_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[103\]
+ sky130_fd_sc_hd__dfxtp_1
X_15313_ _03548_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__clkbuf_1
X_12525_ fifo_bank_register.bank\[3\]\[61\] _05399_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16293_ _04220_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18032_ net431 _01475_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_15244_ _03329_ _03361_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12456_ _07518_ vssd1 vssd1 vccd1 vccd1 _00949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11407_ _06964_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15175_ _03415_ _03439_ _05198_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12387_ _07480_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14126_ fifo_bank_register.bank\[5\]\[63\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[63\]
+ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__a22o_1
X_11338_ fifo_bank_register.bank\[7\]\[13\] _05297_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14057_ _02437_ fifo_bank_register.data_out\[55\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02438_ sky130_fd_sc_hd__mux2_1
X_11269_ _06890_ vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ fifo_bank_register.bank\[1\]\[33\] _05340_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17816_ net560 _01259_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17747_ net516 _01190_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_14959_ _03218_ _03233_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__xor2_1
XFILLER_0_222_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08480_ _04557_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_221_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17678_ net544 _01121_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16629_ net518 _00077_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09101_ sbox1.alph\[0\] _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09032_ _05044_ _05049_ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__and3_2
XFILLER_0_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09934_ _05775_ vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09865_ net23 mix1.data_o\[11\] _05699_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__mux2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _04670_ _04838_ _04839_ _04675_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_198_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09796_ _05651_ vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__clkbuf_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08747_ addroundkey_data_o\[105\] mix1.data_o\[105\] _04655_ vssd1 vssd1 vccd1 vccd1
+ _04771_ sky130_fd_sc_hd__mux2_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_206 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 net229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_239 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08678_ _04656_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__buf_4
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10640_ _06381_ _06407_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10571_ _06347_ _06348_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12310_ _07440_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13290_ _07958_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12241_ _07404_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12172_ _07368_ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11123_ _06791_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__buf_4
XFILLER_0_124_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16980_ net506 _00423_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11054_ _06777_ vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__clkbuf_1
X_15931_ _03905_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__buf_4
XTAP_5131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10005_ sub1.data_o\[25\] _05838_ _05819_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__mux2_1
XTAP_5164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15862_ _04365_ _04687_ _04364_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17601_ net438 _01044_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ _03083_ _03088_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__nor2_4
XTAP_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18581_ clknet_leaf_65_clk _02010_ net590 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ mix1.data_o\[97\] net759 _03819_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__mux2_1
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17532_ net556 _00975_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ ks1.col\[24\] _05547_ _04911_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ fifo_bank_register.bank\[5\]\[49\] _05373_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07254_ sky130_fd_sc_hd__mux2_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10907_ _06491_ _06650_ _06651_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17463_ net469 _00906_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
X_11887_ _07217_ vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__clkbuf_1
X_14675_ fifo_bank_register.bank\[0\]\[124\] _02986_ _08120_ vssd1 vssd1 vccd1 vccd1
+ _02987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16414_ net804 _03961_ _04281_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ fifo_bank_register.bank\[0\]\[9\] _08187_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08188_ sky130_fd_sc_hd__mux2_1
X_10838_ addroundkey_data_o\[106\] _06590_ _06522_ vssd1 vssd1 vccd1 vccd1 _06591_
+ sky130_fd_sc_hd__mux2_1
X_17394_ net389 _00837_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16345_ ks1.key_reg\[72\] _03981_ _04240_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10769_ mix1.data_o\[100\] _06494_ _06398_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__o21a_1
X_13557_ fifo_bank_register.bank\[1\]\[1\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12508_ fifo_bank_register.bank\[3\]\[53\] _05382_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07546_ sky130_fd_sc_hd__mux2_1
X_13488_ fifo_bank_register.read_ptr\[0\] fifo_bank_register.read_ptr\[1\] vssd1 vssd1
+ vccd1 vccd1 _08066_ sky130_fd_sc_hd__or2b_1
X_16276_ net677 _04136_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18015_ net531 _01458_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[17\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_180_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15227_ _03217_ _03486_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__xnor2_2
X_12439_ fifo_bank_register.bank\[3\]\[20\] _05311_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15158_ _03144_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14109_ _02484_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__clkbuf_1
X_15089_ _03357_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__nor2_8
XFILLER_0_227_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09650_ net157 vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__clkbuf_4
X_08601_ first_round_reg _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09581_ fifo_bank_register.bank\[9\]\[101\] _05483_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08532_ _04584_ vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_171_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08463_ _04548_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08394_ _04478_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__buf_8
XFILLER_0_174_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ addroundkey_data_o\[10\] mix1.data_o\[10\] _04805_ vssd1 vssd1 vccd1 vccd1
+ _05037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold130 ks1.key_reg\[85\] vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold141 ks1.key_reg\[48\] vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 ks1.key_reg\[88\] vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 ks1.key_reg\[50\] vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 ks1.key_reg\[91\] vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_217_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout610 net611 vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__clkbuf_4
Xfanout621 net626 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_4
X_09917_ sub1.data_o\[16\] _05753_ _05756_ _05759_ _04611_ vssd1 vssd1 vccd1 vccd1
+ _05760_ sky130_fd_sc_hd__a221o_1
Xfanout632 net633 vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_217_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout643 net646 vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__clkbuf_4
Xfanout654 net655 vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__clkbuf_4
Xfanout665 net666 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09848_ addroundkey_data_o\[9\] _05695_ _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__mux2_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09779_ addroundkey_data_o\[1\] _05636_ next_addroundkey_ready_o vssd1 vssd1 vccd1
+ vccd1 _05637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _07176_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__clkbuf_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _07694_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__clkbuf_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11741_ _07140_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__clkbuf_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _07104_ vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__clkbuf_1
X_14460_ _02142_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__clkbuf_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10623_ _06395_ _06342_ sub1.data_o\[86\] _06384_ vssd1 vssd1 vccd1 vccd1 _06396_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13411_ _05472_ fifo_bank_register.bank\[0\]\[96\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14391_ fifo_bank_register.bank\[5\]\[92\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[92\]
+ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_21_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13342_ _05403_ fifo_bank_register.bank\[0\]\[63\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07986_ sky130_fd_sc_hd__mux2_1
X_16130_ ks1.col\[21\] _04083_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__xor2_2
X_10554_ mix1.data_o\[80\] _06129_ _06093_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ _05333_ fifo_bank_register.bank\[0\]\[30\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07950_ sky130_fd_sc_hd__mux2_1
X_16061_ _04020_ _04022_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10485_ addroundkey_data_o\[72\] _06271_ _06248_ vssd1 vssd1 vccd1 vccd1 _06272_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15012_ _03232_ _03280_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_161_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12224_ _07395_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12155_ _05301_ fifo_bank_register.bank\[4\]\[15\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07359_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11106_ _06805_ vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__clkbuf_1
X_12086_ _07322_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__clkbuf_1
X_16963_ net495 _00406_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15914_ sub1.data_o\[42\] _03576_ _03892_ sub1.data_o\[106\] vssd1 vssd1 vccd1 vccd1
+ _03895_ sky130_fd_sc_hd__a22o_1
X_11037_ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16894_ net571 _00337_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18633_ clknet_leaf_1_clk _02062_ net622 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15845_ mix1.data_o\[122\] net684 _03729_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ clknet_leaf_63_clk _01993_ net598 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[91\]
+ sky130_fd_sc_hd__dfrtp_1
X_15776_ _03741_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__clkbuf_8
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _07799_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ net414 _00958_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_14727_ _03019_ _04927_ _05245_ _03027_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__a31o_1
X_11939_ _07245_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18495_ clknet_leaf_59_clk _01924_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17446_ net448 _00889_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
X_14658_ fifo_bank_register.bank\[9\]\[122\] _08089_ _02969_ _02970_ _02971_ vssd1
+ vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_156_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13609_ _08171_ fifo_bank_register.data_out\[7\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _08173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17377_ net499 _00820_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14589_ fifo_bank_register.bank\[5\]\[114\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[114\]
+ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_clk clknet_3_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16328_ net845 _03909_ _04222_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16259_ net824 _03912_ _04106_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput268 net268 vssd1 vssd1 vccd1 vccd1 data_o[107] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput279 net279 vssd1 vssd1 vccd1 vccd1 data_o[117] sky130_fd_sc_hd__buf_2
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_79_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09702_ _05566_ vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09633_ fifo_bank_register.bank\[9\]\[118\] _05518_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09564_ net253 vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ _04575_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09495_ _05425_ vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08446_ _04539_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08377_ _04503_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10270_ sub1.data_o\[51\] _06077_ _05936_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout440 net443 vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_1
Xfanout451 net461 vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_2
Xfanout462 net466 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__clkbuf_2
Xfanout473 net474 vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__buf_2
X_13960_ fifo_bank_register.bank\[5\]\[45\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[45\]
+ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__a22o_1
Xfanout484 net489 vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__clkbuf_2
Xfanout495 net498 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_2
X_12911_ fifo_bank_register.bank\[2\]\[116\] _05514_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13891_ _08068_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__buf_4
X_15630_ mix1.data_o\[19\] _03497_ _03742_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ fifo_bank_register.bank\[2\]\[83\] _05445_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15561_ sub1.data_o\[69\] _03691_ _03703_ _03594_ vssd1 vssd1 vccd1 vccd1 _03704_
+ sky130_fd_sc_hd__a22o_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ fifo_bank_register.bank\[2\]\[50\] _05375_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ net517 _00743_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _02842_ fifo_bank_register.data_out\[105\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02843_ sky130_fd_sc_hd__mux2_1
X_18280_ clknet_leaf_1_clk _01711_ net583 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[46\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _07131_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__clkbuf_1
X_15492_ sub1.data_o\[109\] _03600_ _03653_ sub1.data_o\[45\] vssd1 vssd1 vccd1 vccd1
+ _03659_ sky130_fd_sc_hd__a22o_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17231_ net479 _00674_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11655_ _07095_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__clkbuf_1
X_14443_ fifo_bank_register.bank\[1\]\[98\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[98\]
+ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17162_ net521 _00605_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
X_10606_ _06380_ vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11586_ fifo_bank_register.bank\[6\]\[2\] _05274_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07059_ sky130_fd_sc_hd__mux2_1
X_14374_ fifo_bank_register.bank\[6\]\[90\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[90\]
+ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16113_ net239 ks1.key_reg\[83\] _03906_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__mux2_2
X_10537_ net105 mix1.data_o\[79\] _06316_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__mux2_1
X_13325_ _05386_ fifo_bank_register.bank\[0\]\[55\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17093_ net441 _00536_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16044_ _04003_ _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__xnor2_2
X_13256_ _05317_ fifo_bank_register.bank\[0\]\[22\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07941_ sky130_fd_sc_hd__mux2_1
X_10468_ _06255_ _06256_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__xor2_1
XFILLER_0_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12207_ _07386_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13187_ _07903_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__clkbuf_1
X_10399_ sub1.data_o\[63\] _06194_ _06160_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12138_ _05284_ fifo_bank_register.bank\[4\]\[7\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17995_ net442 _01438_ net602 vssd1 vssd1 vccd1 vccd1 fifo_bank_register.write_ptr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_202_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16946_ net452 _00389_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
X_12069_ _07313_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16877_ net415 _00320_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18616_ clknet_leaf_83_clk _02045_ net584 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[109\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15828_ _03846_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__clkbuf_1
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18547_ clknet_leaf_77_clk _01976_ net589 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15759_ _03810_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08300_ net199 net201 net200 net198 vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__or4bb_1
X_09280_ _05279_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__clkbuf_1
X_18478_ clknet_leaf_57_clk _01907_ net602 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08231_ net119 net118 net121 net120 vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17429_ net553 _00872_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ addroundkey_data_o\[122\] mix1.data_o\[122\] _04657_ vssd1 vssd1 vccd1 vccd1
+ _05017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09616_ _05507_ vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09547_ fifo_bank_register.bank\[9\]\[90\] _05459_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ fifo_bank_register.bank\[9\]\[68\] _05413_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08429_ _04530_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_1
XFILLER_0_108_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11440_ fifo_bank_register.bank\[7\]\[61\] _05399_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11371_ _06945_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10322_ _05574_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__clkbuf_4
X_13110_ _07863_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__clkbuf_1
X_14090_ fifo_bank_register.bank\[0\]\[59\] _02466_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ fifo_bank_register.bank\[1\]\[49\] _05373_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07827_ sky130_fd_sc_hd__mux2_1
X_10253_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_219_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10184_ _05615_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__buf_2
XFILLER_0_219_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16800_ clknet_leaf_63_clk _00244_ net598 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[91\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_227_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17780_ net394 _01223_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14992_ _03250_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_156_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16731_ clknet_leaf_42_clk _00175_ net659 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_205_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13943_ _02336_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16662_ net465 _00110_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13874_ fifo_bank_register.bank\[0\]\[35\] _02274_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18401_ clknet_leaf_24_clk _01831_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[86\]
+ sky130_fd_sc_hd__dfrtp_2
X_15613_ _03733_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12825_ fifo_bank_register.bank\[2\]\[75\] _05428_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16593_ net423 _00041_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18332_ clknet_leaf_16_clk _01762_ net637 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_15544_ sub1.data_o\[96\] sub1.data_o\[32\] _03671_ vssd1 vssd1 vccd1 vccd1 _03692_
+ sky130_fd_sc_hd__mux2_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ fifo_bank_register.bank\[2\]\[42\] _05359_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18263_ clknet_leaf_52_clk _01694_ net655 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_127_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11707_ _07122_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__clkbuf_1
X_15475_ sub1.data_o\[38\] _03648_ _03636_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12687_ _07628_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17214_ net441 _00657_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14426_ fifo_bank_register.bank\[1\]\[96\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[96\]
+ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18194_ clknet_leaf_24_clk _01625_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11638_ _07086_ vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17145_ net575 _00588_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_14357_ _08181_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ fifo_bank_register.bank\[7\]\[123\] _05528_ _06912_ vssd1 vssd1 vccd1 vccd1
+ _07049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13308_ _05369_ fifo_bank_register.bank\[0\]\[47\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17076_ net434 _00519_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
X_14288_ _02157_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__buf_4
X_16027_ _04757_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13239_ _07931_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08780_ addroundkey_data_o\[75\] mix1.data_o\[75\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _04804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17978_ net456 _01421_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16929_ net401 _00372_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09401_ fifo_bank_register.bank\[9\]\[43\] _05361_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09332_ net171 vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_133_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _05250_ _05249_ net597 vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__and3b_1
XFILLER_0_168_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08214_ _04372_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__buf_4
X_09194_ sub1.data_o\[115\] _05197_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__a21o_1
XFILLER_0_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold12 ks1.key_reg\[123\] vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold23 mix1.data_reg\[34\] vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold34 ks1.key_reg\[0\] vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ ks1.key_reg\[31\] _04725_ _05001_ net182 vssd1 vssd1 vccd1 vccd1 _05002_
+ sky130_fd_sc_hd__a22o_1
Xhold45 mix1.data_reg\[57\] vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold56 mix1.data_reg\[40\] vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold67 mix1.data_reg\[78\] vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 mix1.data_reg\[82\] vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold89 mix1.data_reg\[97\] vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10940_ _05574_ _06680_ _06681_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__a21o_1
XFILLER_0_168_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_211_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10871_ addroundkey_data_o\[110\] _06619_ _06612_ vssd1 vssd1 vccd1 vccd1 _06620_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12610_ _07599_ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13590_ fifo_bank_register.bank\[9\]\[5\] _08090_ _08153_ _08154_ _08155_ vssd1 vssd1
+ vccd1 vccd1 _08156_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12541_ fifo_bank_register.bank\[3\]\[69\] _05415_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _03394_ _03413_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__xnor2_1
X_12472_ fifo_bank_register.bank\[3\]\[36\] _05346_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14211_ fifo_bank_register.bank\[6\]\[72\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[72\]
+ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11423_ fifo_bank_register.bank\[7\]\[53\] _05382_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06973_ sky130_fd_sc_hd__mux2_1
X_15191_ _03336_ _03454_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_9 _03926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11354_ fifo_bank_register.bank\[7\]\[20\] _05311_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14142_ fifo_bank_register.bank\[5\]\[65\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[65\]
+ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10305_ _06110_ vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14073_ _08068_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__clkbuf_8
X_11285_ _05516_ fifo_bank_register.bank\[8\]\[117\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10236_ _05913_ _05972_ sub1.data_o\[48\] _05902_ vssd1 vssd1 vccd1 vccd1 _06047_
+ sky130_fd_sc_hd__a31o_1
X_17901_ net415 _01344_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_13024_ _07818_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17832_ net448 _01275_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10167_ net192 ks1.key_reg\[40\] _05825_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17763_ net499 _01206_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14975_ _03198_ _03248_ _05201_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__o21ai_1
X_10098_ addroundkey_data_o\[34\] _05922_ _05872_ vssd1 vssd1 vccd1 vccd1 _05923_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16714_ clknet_leaf_41_clk _00158_ net658 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_13926_ _02321_ fifo_bank_register.data_out\[40\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17694_ net541 _01137_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16645_ net567 _00093_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ fifo_bank_register.bank\[9\]\[33\] _02226_ _02257_ _02258_ _02259_ vssd1
+ vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12808_ fifo_bank_register.bank\[2\]\[67\] _05411_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16576_ net496 _00024_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_13788_ fifo_bank_register.bank\[6\]\[26\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__a22o_1
X_18315_ clknet_leaf_9_clk _01745_ net633 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15527_ sub1.data_o\[56\] _05547_ _04884_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__mux2_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ fifo_bank_register.bank\[2\]\[34\] _05342_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18246_ clknet_leaf_10_clk _01677_ net625 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_199_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15458_ _03637_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14409_ fifo_bank_register.bank\[6\]\[94\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[94\]
+ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__a22o_1
X_18177_ clknet_leaf_13_clk _01608_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[71\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ _04689_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17128_ net431 _00571_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17059_ net400 _00502_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_09950_ net168 ks1.key_reg\[19\] _05708_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08901_ addroundkey_data_o\[21\] mix1.data_o\[21\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09881_ _05727_ vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__clkbuf_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ addroundkey_data_o\[70\] mix1.data_o\[70\] _04665_ vssd1 vssd1 vccd1 vccd1
+ _04856_ sky130_fd_sc_hd__mux2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08763_ _04784_ _04785_ _04786_ _04698_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _04699_ _04704_ _04711_ _04717_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09315_ net165 vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__buf_2
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09246_ fifo_bank_register.write_ptr\[1\] vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__buf_2
XFILLER_0_111_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09177_ sbox1.alph\[0\] _05177_ _05155_ sbox1.alph\[3\] vssd1 vssd1 vccd1 vccd1 _05188_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_1_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11070_ _05301_ fifo_bank_register.bank\[8\]\[15\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06786_ sky130_fd_sc_hd__mux2_1
XTAP_6025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput102 data_i[76] vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__buf_2
X_10021_ sub1.data_o\[27\] _05852_ _05819_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__mux2_1
XTAP_6069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput113 data_i[86] vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__buf_4
XTAP_5335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput124 data_i[96] vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_179_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput135 key_i[104] vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__clkbuf_4
Xinput146 key_i[114] vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_4
XTAP_5357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput157 key_i[124] vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_4
XTAP_5379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput168 key_i[19] vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_4
XTAP_4645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput179 key_i[29] vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_4
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ ks1.col\[16\] _05547_ _00007_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__mux2_1
XTAP_4689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11972_ _07262_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__clkbuf_1
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _08181_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__clkbuf_4
X_10923_ _06665_ _06666_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__xnor2_1
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ fifo_bank_register.bank\[0\]\[126\] _03000_ _08120_ vssd1 vssd1 vccd1 vccd1
+ _03001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16430_ _04372_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__buf_4
X_13642_ _08120_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__buf_4
XFILLER_0_224_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10854_ addroundkey_data_o\[108\] _06604_ _06522_ vssd1 vssd1 vccd1 vccd1 _06605_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ ks1.next_ready_o _04039_ _04256_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_184_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13573_ fifo_bank_register.bank\[1\]\[3\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ addroundkey_data_o\[101\] _06542_ _06522_ vssd1 vssd1 vccd1 vccd1 _06543_
+ sky130_fd_sc_hd__mux2_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18100_ net466 _01543_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15312_ net726 _03411_ _03539_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ _07554_ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__clkbuf_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ net830 _04040_ _04206_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18031_ net426 _01474_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_15243_ _03499_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12455_ fifo_bank_register.bank\[3\]\[28\] _05329_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11406_ fifo_bank_register.bank\[7\]\[45\] _05365_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06964_ sky130_fd_sc_hd__mux2_1
X_15174_ _03406_ _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ _05532_ fifo_bank_register.bank\[4\]\[125\] _07341_ vssd1 vssd1 vccd1 vccd1
+ _07480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ _02498_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11337_ _06927_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14056_ fifo_bank_register.bank\[0\]\[55\] _02436_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02437_ sky130_fd_sc_hd__mux2_1
X_11268_ _05499_ fifo_bank_register.bank\[8\]\[109\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13007_ _07809_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10219_ sub1.data_o\[46\] _06031_ _05991_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__mux2_1
X_11199_ _05430_ fifo_bank_register.bank\[8\]\[76\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17815_ net561 _01258_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17746_ net504 _01189_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_14958_ _03225_ _03232_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_168_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ _02305_ fifo_bank_register.data_out\[39\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17677_ net517 _01120_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
X_14889_ addroundkey_data_o\[31\] _04375_ _04900_ _03164_ vssd1 vssd1 vccd1 vccd1
+ _03165_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16628_ net511 _00076_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16559_ clknet_leaf_49_clk _00007_ net615 vssd1 vssd1 vccd1 vccd1 ks1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09100_ _05109_ _05110_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__nand2_2
XFILLER_0_169_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09031_ _04863_ _05050_ _05052_ _04741_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__o2bb2a_1
X_18229_ clknet_leaf_38_clk _01660_ net668 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09933_ addroundkey_data_o\[17\] _05774_ _05697_ vssd1 vssd1 vccd1 vccd1 _05775_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09864_ _05615_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__clkbuf_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ addroundkey_data_o\[30\] mix1.data_o\[30\] _04665_ vssd1 vssd1 vccd1 vccd1
+ _04839_ sky130_fd_sc_hd__mux2_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ addroundkey_data_o\[3\] _05650_ next_addroundkey_ready_o vssd1 vssd1 vccd1
+ vccd1 _05651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08746_ addroundkey_data_o\[81\] mix1.data_o\[81\] _04654_ vssd1 vssd1 vccd1 vccd1
+ _04770_ sky130_fd_sc_hd__mux2_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_207 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _04700_ _04681_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nor2_4
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_229 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ net237 ks1.key_reg\[81\] _06097_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__mux2_4
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09229_ sub1.data_o\[22\] _05200_ _05203_ sub1.data_o\[86\] vssd1 vssd1 vccd1 vccd1
+ _05237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12240_ _05386_ fifo_bank_register.bank\[4\]\[55\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ _05317_ fifo_bank_register.bank\[4\]\[22\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11122_ _06813_ vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11053_ _05284_ fifo_bank_register.bank\[8\]\[7\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15930_ _04742_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__buf_4
XTAP_5110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10004_ net46 mix1.data_o\[25\] _05817_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15861_ _04365_ _04700_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__xnor2_1
XTAP_5165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17600_ net492 _01043_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14812_ addroundkey_data_o\[120\] _03079_ _03087_ vssd1 vssd1 vccd1 vccd1 _03088_
+ sky130_fd_sc_hd__a21oi_1
XTAP_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18580_ clknet_leaf_75_clk _02009_ net588 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15792_ _03827_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__clkbuf_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17531_ net562 _00974_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14743_ _03035_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__clkbuf_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _07253_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_169_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10906_ _06630_ _06514_ sub1.data_o\[114\] _05675_ vssd1 vssd1 vccd1 vccd1 _06651_
+ sky130_fd_sc_hd__a31o_1
X_17462_ net411 _00905_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
X_14674_ fifo_bank_register.bank\[9\]\[124\] _08089_ _02983_ _02984_ _02985_ vssd1
+ vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11886_ fifo_bank_register.bank\[5\]\[16\] _05303_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16413_ _04286_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ fifo_bank_register.bank\[9\]\[9\] _08090_ _08184_ _08185_ _08186_ vssd1 vssd1
+ vccd1 vccd1 _08187_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17393_ net393 _00836_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_10837_ _06588_ _06589_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__xor2_1
XFILLER_0_184_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16344_ _04247_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_229_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ fifo_bank_register.bank\[6\]\[1\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10768_ _06491_ _06525_ _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12507_ _07545_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__clkbuf_1
X_16275_ _04210_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__clkbuf_1
X_13487_ fifo_bank_register.read_ptr\[1\] fifo_bank_register.read_ptr\[0\] vssd1 vssd1
+ vccd1 vccd1 _08065_ sky130_fd_sc_hd__or2b_1
X_10699_ mix1.data_o\[94\] _06463_ _06320_ _06321_ sub1.data_o\[94\] vssd1 vssd1 vccd1
+ vccd1 _06464_ sky130_fd_sc_hd__a32o_1
X_18014_ net471 _01457_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[16\]
+ sky130_fd_sc_hd__dfxtp_4
X_15226_ _03153_ _03246_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ _07508_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15157_ _03415_ _03423_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__xor2_4
XFILLER_0_160_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12369_ _07471_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14108_ _02483_ fifo_bank_register.data_out\[60\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15088_ addroundkey_data_o\[108\] _03057_ _03359_ vssd1 vssd1 vccd1 vccd1 _03360_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14039_ fifo_bank_register.bank\[9\]\[53\] _02388_ _02419_ _02420_ _02421_ vssd1
+ vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_219_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08600_ _04625_ _04626_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__nand2_2
X_09580_ net132 vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__buf_2
XFILLER_0_222_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08531_ addroundkey_data_o\[104\] fifo_bank_register.data_out\[104\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17729_ net439 _01172_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08462_ addroundkey_data_o\[71\] fifo_bank_register.data_out\[71\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08393_ _04511_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09014_ addroundkey_data_o\[106\] mix1.data_o\[106\] _04665_ vssd1 vssd1 vccd1 vccd1
+ _05036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold120 mix1.data_reg\[119\] vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold131 ks1.key_reg\[119\] vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 ks1.key_reg\[104\] vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 ks1.key_reg\[69\] vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 ks1.key_reg\[49\] vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 ks1.key_reg\[64\] vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout600 net601 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_217_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout611 net612 vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09916_ mix1.data_o\[16\] _05576_ _05758_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__o21a_1
Xfanout622 net626 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__buf_2
XFILLER_0_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout633 net634 vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout644 net646 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout655 net657 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout666 net667 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_4
X_09847_ _05696_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__buf_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09778_ _05634_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ ks1.key_reg\[17\] _04730_ _04732_ net166 vssd1 vssd1 vccd1 vccd1 _04753_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_217_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11740_ fifo_bank_register.bank\[6\]\[75\] _05428_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07140_ sky130_fd_sc_hd__mux2_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ fifo_bank_register.bank\[6\]\[42\] _05359_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13410_ _08021_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__clkbuf_1
X_10622_ _04624_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1086 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14390_ _02734_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13341_ _07985_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10553_ _06126_ _06330_ _06331_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16060_ _05227_ _04021_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13272_ _07937_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__buf_4
X_10484_ _06269_ _06270_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15011_ _03284_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12223_ _05369_ fifo_bank_register.bank\[4\]\[47\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12154_ _07358_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11105_ _05336_ fifo_bank_register.bank\[8\]\[31\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12085_ fifo_bank_register.bank\[5\]\[110\] _05501_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07322_ sky130_fd_sc_hd__mux2_1
X_16962_ net471 _00405_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15913_ _03717_ _04943_ _05554_ _03894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__a31o_1
X_11036_ fifo_bank_register.write_ptr\[2\] _05254_ _06765_ _06766_ vssd1 vssd1 vccd1
+ vccd1 _06767_ sky130_fd_sc_hd__or4_2
X_16893_ net571 _00336_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15844_ _03854_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__clkbuf_1
X_18632_ clknet_leaf_36_clk _02061_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ _03818_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__clkbuf_1
X_18563_ clknet_leaf_63_clk _01992_ net598 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ fifo_bank_register.bank\[1\]\[23\] _05319_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07799_ sky130_fd_sc_hd__mux2_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ sub1.data_o\[87\] _03010_ _03026_ sub1.next_ready_o vssd1 vssd1 vccd1 vccd1
+ _03027_ sky130_fd_sc_hd__a22o_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17514_ net422 _00957_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11938_ fifo_bank_register.bank\[5\]\[40\] _05354_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18494_ clknet_leaf_56_clk _01923_ net614 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17445_ net402 _00888_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14657_ fifo_bank_register.bank\[1\]\[122\] _08111_ _08114_ fifo_bank_register.bank\[8\]\[122\]
+ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__a22o_1
X_11869_ fifo_bank_register.bank\[5\]\[8\] _05286_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13608_ _08068_ vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17376_ net483 _00819_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14588_ _02910_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16327_ _04215_ _04199_ _04238_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__o21ai_1
X_13539_ _08056_ _08087_ vssd1 vssd1 vccd1 vccd1 _08110_ sky130_fd_sc_hd__and2b_1
XFILLER_0_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16258_ _04201_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15209_ _03361_ _03394_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__xor2_2
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16189_ _04112_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput269 net269 vssd1 vssd1 vccd1 vccd1 data_o[108] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09701_ sub1.data_o\[127\] _05245_ _04891_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09632_ net150 vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_156_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09563_ _05471_ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08514_ addroundkey_data_o\[96\] fifo_bank_register.data_out\[96\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__mux2_2
XFILLER_0_136_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09494_ fifo_bank_register.bank\[9\]\[73\] _05424_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08445_ addroundkey_data_o\[63\] fifo_bank_register.data_out\[63\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08376_ addroundkey_data_o\[30\] fifo_bank_register.data_out\[30\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__mux2_2
XFILLER_0_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout430 net431 vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__buf_2
Xfanout441 net442 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_2
Xfanout452 net461 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__buf_2
Xfanout463 net466 vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_217_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout474 net481 vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__buf_2
Xfanout485 net489 vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_2
XFILLER_0_226_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12910_ _07757_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__clkbuf_1
Xfanout496 net498 vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_2
X_13890_ fifo_bank_register.bank\[0\]\[37\] _02288_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12841_ _07721_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__clkbuf_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15560_ sub1.data_o\[101\] sub1.data_o\[37\] _03574_ vssd1 vssd1 vccd1 vccd1 _03703_
+ sky130_fd_sc_hd__mux2_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _07651_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__buf_4
XFILLER_0_154_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ fifo_bank_register.bank\[0\]\[105\] _02841_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ fifo_bank_register.bank\[6\]\[67\] _05411_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07131_ sky130_fd_sc_hd__mux2_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _03652_ _04784_ _05219_ _03658_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a31o_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ net492 _00673_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14442_ fifo_bank_register.bank\[6\]\[98\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[98\]
+ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a22o_1
X_11654_ fifo_bank_register.bank\[6\]\[34\] _05342_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17161_ net514 _00604_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_10605_ addroundkey_data_o\[84\] _06379_ _06327_ vssd1 vssd1 vccd1 vccd1 _06380_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14373_ _02148_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__clkbuf_4
X_11585_ _07058_ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16112_ ks1.col\[19\] _04067_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__xor2_4
X_13324_ _07976_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _05749_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__buf_4
X_17092_ net494 _00535_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16043_ _04004_ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__xnor2_2
X_13255_ _07940_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__clkbuf_1
X_10467_ net225 ks1.key_reg\[70\] _06245_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12206_ _05352_ fifo_bank_register.bank\[4\]\[39\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07386_ sky130_fd_sc_hd__mux2_1
X_13186_ fifo_bank_register.bank\[1\]\[118\] _05518_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ net88 mix1.data_o\[63\] _06158_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12137_ _07349_ vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17994_ net442 _01437_ net597 vssd1 vssd1 vccd1 vccd1 fifo_bank_register.write_ptr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16945_ net451 _00388_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
X_12068_ fifo_bank_register.bank\[5\]\[102\] _05485_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11019_ sub1.data_o\[126\] _06751_ _05609_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__mux2_1
X_16876_ net416 _00319_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18615_ clknet_leaf_83_clk _02044_ net582 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[108\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15827_ mix1.data_o\[113\] net738 _03841_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__mux2_1
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15758_ mix1.data_o\[80\] net778 _03808_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__mux2_1
X_18546_ clknet_leaf_63_clk _01975_ net599 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[73\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14709_ sub1.data_o\[50\] sub1.data_o\[114\] _05598_ vssd1 vssd1 vccd1 vccd1 _03015_
+ sky130_fd_sc_hd__mux2_1
X_15689_ _03773_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18477_ clknet_leaf_58_clk _01906_ net602 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ _04383_ _04384_ _04385_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17428_ net525 _00871_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17359_ net478 _00802_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08994_ _04971_ _05016_ vssd1 vssd1 vccd1 vccd1 sbox1.ah\[1\] sky130_fd_sc_hd__xnor2_4
XFILLER_0_228_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09615_ fifo_bank_register.bank\[9\]\[112\] _05506_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09546_ _05312_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ net222 vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__buf_2
XFILLER_0_210_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08428_ addroundkey_data_o\[55\] fifo_bank_register.data_out\[55\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08359_ addroundkey_data_o\[22\] fifo_bank_register.data_out\[22\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11370_ fifo_bank_register.bank\[7\]\[28\] _05329_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10321_ sub1.data_o\[55\] _06124_ _06113_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13040_ _07826_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__clkbuf_1
X_10252_ net201 ks1.key_reg\[49\] _05920_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__mux2_4
XFILLER_0_218_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10183_ _06000_ vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_218_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14991_ _03257_ _03264_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_227_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16730_ clknet_leaf_41_clk _00174_ net659 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_13942_ _02335_ fifo_bank_register.data_out\[42\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16661_ net450 _00109_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13873_ fifo_bank_register.bank\[9\]\[35\] _02226_ _02271_ _02272_ _02273_ vssd1
+ vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18400_ clknet_leaf_24_clk _01830_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[85\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_199_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15612_ mix1.data_o\[11\] _03446_ _03730_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__mux2_1
X_12824_ _07712_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__clkbuf_1
X_16592_ net423 _00040_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15543_ _04368_ _04935_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__nor2_2
X_18331_ clknet_leaf_16_clk _01761_ net630 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _07676_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__clkbuf_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18262_ clknet_leaf_43_clk _01693_ net658 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ fifo_bank_register.bank\[6\]\[59\] _05394_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07122_ sky130_fd_sc_hd__mux2_1
X_15474_ sub1.data_o\[70\] _05235_ _03633_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__mux2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _07639_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17213_ net435 _00656_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14425_ fifo_bank_register.bank\[6\]\[96\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[96\]
+ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__a22o_1
X_18193_ clknet_leaf_24_clk _01624_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_11637_ fifo_bank_register.bank\[6\]\[26\] _05325_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17144_ net572 _00587_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_14356_ _02703_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__clkbuf_1
X_11568_ _07048_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13307_ _07967_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17075_ net455 _00518_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
X_10519_ _06301_ vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14287_ fifo_bank_register.bank\[9\]\[80\] _02631_ _02636_ _02639_ _02642_ vssd1
+ vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_208_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11499_ _07012_ vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16026_ _03990_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__xnor2_2
X_13238_ _05299_ fifo_bank_register.bank\[0\]\[14\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13169_ _07794_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17977_ net470 _01420_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16928_ net409 _00371_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16859_ net484 _00302_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09400_ net195 vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__buf_2
XFILLER_0_215_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09331_ _05314_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__clkbuf_1
X_18529_ clknet_leaf_66_clk _01958_ net606 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _05257_ _05259_ _05261_ _05265_ net258 vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__o41a_4
XFILLER_0_34_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08213_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09193_ sub1.data_o\[19\] _05200_ _05203_ sub1.data_o\[83\] vssd1 vssd1 vccd1 vccd1
+ _05204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold13 ks1.key_reg\[41\] vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold24 mix1.data_reg\[32\] vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ ks1.key_reg\[31\] _04729_ _04731_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__or3_1
XTAP_4805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold35 mix1.state\[0\] vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_216_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold46 mix1.data_reg\[94\] vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold57 mix1.data_reg\[74\] vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold68 mix1.data_reg\[113\] vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold79 mix1.data_reg\[114\] vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_199_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10870_ _06617_ _06618_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _05448_ vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _07562_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_213_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12471_ _07526_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ fifo_bank_register.bank\[7\]\[72\] _02542_ _02551_ fifo_bank_register.bank\[2\]\[72\]
+ _02573_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a221o_1
X_11422_ _06972_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15190_ _03410_ _03453_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14141_ _02512_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11353_ _06935_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10304_ addroundkey_data_o\[53\] _06109_ _06064_ vssd1 vssd1 vccd1 vccd1 _06110_
+ sky130_fd_sc_hd__mux2_1
X_14072_ fifo_bank_register.bank\[0\]\[57\] _02450_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11284_ _06898_ vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13023_ fifo_bank_register.bank\[1\]\[40\] _05354_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07818_ sky130_fd_sc_hd__mux2_1
X_17900_ net428 _01343_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
X_10235_ sub1.data_o\[48\] _06045_ _05936_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17831_ net454 _01274_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
X_10166_ _05829_ _05983_ _05984_ _05833_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17762_ net486 _01205_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14974_ _03238_ _03247_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__xnor2_1
X_10097_ _05919_ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__xnor2_1
X_16713_ clknet_leaf_51_clk _00157_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_13925_ fifo_bank_register.bank\[0\]\[40\] _02319_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17693_ net538 _01136_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13856_ fifo_bank_register.bank\[1\]\[33\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[33\]
+ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__a22o_1
X_16644_ net550 _00092_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12807_ _07703_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13787_ fifo_bank_register.bank\[7\]\[26\] _02128_ _02139_ fifo_bank_register.bank\[2\]\[26\]
+ _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__a221o_1
X_16575_ net534 _00023_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10999_ _06733_ _06734_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18314_ clknet_leaf_21_clk sub1.next_ready_o net643 vssd1 vssd1 vccd1 vccd1 sub1.ready_o
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15526_ _03668_ _04777_ _05245_ _03682_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _07667_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__clkbuf_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15457_ sub1.data_o\[32\] _03634_ _03636_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__mux2_1
X_18245_ clknet_leaf_2_clk _01676_ net625 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_12669_ fifo_bank_register.bank\[2\]\[1\] _05272_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14408_ fifo_bank_register.bank\[7\]\[94\] _02704_ _02713_ fifo_bank_register.bank\[2\]\[94\]
+ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15388_ _03592_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18176_ clknet_leaf_13_clk _01607_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[70\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17127_ net423 _00570_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_14339_ _02688_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ net410 _00501_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08900_ addroundkey_data_o\[125\] mix1.data_o\[125\] _04658_ vssd1 vssd1 vccd1 vccd1
+ _04924_ sky130_fd_sc_hd__mux2_1
X_16009_ _04742_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09880_ addroundkey_data_o\[12\] _05726_ _05697_ vssd1 vssd1 vccd1 vccd1 _05727_
+ sky130_fd_sc_hd__mux2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08831_ _04706_ _04853_ _04854_ _04710_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__a22o_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ addroundkey_data_o\[25\] _04675_ _04670_ addroundkey_data_o\[49\] vssd1 vssd1
+ vccd1 vccd1 _04786_ sky130_fd_sc_hd__a22o_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08693_ _04713_ _04714_ _04715_ _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09314_ _05302_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09245_ fifo_bank_register.write_ptr\[0\] vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__buf_2
XFILLER_0_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09176_ _05185_ _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10020_ net48 mix1.data_o\[27\] _05817_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__mux2_1
XTAP_6059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput103 data_i[77] vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_4
XTAP_5325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput114 data_i[87] vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__buf_4
XTAP_5336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput125 data_i[97] vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_8
Xinput136 key_i[105] vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_4
XTAP_5347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput147 key_i[115] vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_4
XFILLER_0_76_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput158 key_i[125] vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_4
XTAP_5369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput169 key_i[1] vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_4
XTAP_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ fifo_bank_register.bank\[5\]\[56\] _05388_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13710_ _02127_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__clkbuf_1
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10922_ net147 ks1.key_reg\[115\] _04639_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__mux2_2
XFILLER_0_169_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14690_ fifo_bank_register.bank\[9\]\[126\] _08089_ _02997_ _02998_ _02999_ vssd1
+ vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__a2111o_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ fifo_bank_register.bank\[9\]\[10\] _08190_ _08195_ _08198_ _08201_ vssd1
+ vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_211_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10853_ _06602_ _06603_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ net685 _04373_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13572_ fifo_bank_register.bank\[6\]\[3\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _06540_ _06541_ vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _03547_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12523_ fifo_bank_register.bank\[3\]\[60\] _05396_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07554_ sky130_fd_sc_hd__mux2_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16291_ _04219_ vssd1 vssd1 vccd1 vccd1 _01948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ net786 _03497_ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__mux2_1
X_18030_ net416 _01473_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_12454_ _07517_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11405_ _06963_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__clkbuf_1
X_15173_ _03394_ _03437_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__xnor2_4
X_12385_ _07479_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14124_ _02497_ fifo_bank_register.data_out\[62\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11336_ fifo_bank_register.bank\[7\]\[12\] _05295_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14055_ fifo_bank_register.bank\[9\]\[55\] _02388_ _02433_ _02434_ _02435_ vssd1
+ vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__a2111o_1
X_11267_ _06889_ vssd1 vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13006_ fifo_bank_register.bank\[1\]\[32\] _05338_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10218_ net69 mix1.data_o\[46\] _05989_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11198_ _06853_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17814_ net566 _01257_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
X_10149_ net61 mix1.data_o\[39\] _05934_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17745_ net533 _01188_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14957_ _03228_ _03231_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__nor2_4
XFILLER_0_222_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13908_ fifo_bank_register.bank\[0\]\[39\] _02304_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02305_ sky130_fd_sc_hd__mux2_1
X_17676_ net519 _01119_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14888_ addroundkey_data_o\[95\] _03061_ _03065_ addroundkey_data_o\[63\] vssd1 vssd1
+ vccd1 vccd1 _03164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16627_ net521 _00075_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13839_ fifo_bank_register.bank\[6\]\[31\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16558_ clknet_leaf_54_clk _00006_ net615 vssd1 vssd1 vccd1 vccd1 ks1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15509_ _03668_ _04777_ _05560_ _03670_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16489_ net717 _03392_ _04321_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09030_ ks1.key_reg\[18\] _04735_ _05051_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__a21oi_1
X_18228_ clknet_leaf_37_clk _01659_ net666 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18159_ clknet_leaf_48_clk _01590_ net610 vssd1 vssd1 vccd1 vccd1 ks1.col\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09932_ _05772_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09863_ _05711_ vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__clkbuf_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ addroundkey_data_o\[54\] mix1.data_o\[54\] _04662_ vssd1 vssd1 vccd1 vccd1
+ _04838_ sky130_fd_sc_hd__mux2_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _05648_ _05649_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__xor2_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08745_ _04682_ _04767_ _04701_ _04768_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08676_ _04362_ _04363_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_219 net205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09228_ _05235_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09159_ _05164_ _05169_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_82_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12170_ _07367_ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11121_ _05352_ fifo_bank_register.bank\[8\]\[39\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11052_ _06776_ vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__clkbuf_1
XTAP_5111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10003_ _05837_ vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__clkbuf_1
XTAP_5144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15860_ _04705_ _04680_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14811_ addroundkey_data_o\[88\] _03072_ _03085_ _03086_ vssd1 vssd1 vccd1 vccd1
+ _03087_ sky130_fd_sc_hd__a211o_1
XTAP_5199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ mix1.data_o\[96\] net739 _03819_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__mux2_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17530_ net562 _00973_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11954_ fifo_bank_register.bank\[5\]\[48\] _05371_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07253_ sky130_fd_sc_hd__mux2_1
X_14742_ ks1.col\[7\] _05244_ _04916_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10905_ sub1.data_o\[114\] _06649_ _05608_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__mux2_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17461_ net411 _00904_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
X_14673_ fifo_bank_register.bank\[1\]\[124\] _08111_ _08114_ fifo_bank_register.bank\[8\]\[124\]
+ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__a22o_1
XFILLER_0_212_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ _07216_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13624_ fifo_bank_register.bank\[1\]\[9\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__a22o_1
X_16412_ ks1.key_reg\[101\] _03951_ _04281_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10836_ net137 ks1.key_reg\[106\] _06579_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17392_ net398 _00835_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13555_ fifo_bank_register.bank\[7\]\[1\] _08078_ _08093_ fifo_bank_register.bank\[2\]\[1\]
+ _08124_ vssd1 vssd1 vccd1 vccd1 _08125_ sky130_fd_sc_hd__a221o_1
X_16343_ net829 _03971_ _04240_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ _06395_ _06514_ sub1.data_o\[100\] _06384_ vssd1 vssd1 vccd1 vccd1 _06526_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ fifo_bank_register.bank\[3\]\[52\] _05380_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07545_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16274_ ks1.key_reg\[39\] _03973_ _04206_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13486_ fifo_bank_register.read_ptr\[0\] _08064_ vssd1 vssd1 vccd1 vccd1 _01433_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10698_ _05585_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15225_ _03485_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__clkbuf_1
X_18013_ net535 _01456_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_12437_ _07484_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__buf_6
XFILLER_0_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15156_ _03285_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__xor2_4
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12368_ _05514_ fifo_bank_register.bank\[4\]\[116\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14107_ fifo_bank_register.bank\[0\]\[60\] _02481_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02483_ sky130_fd_sc_hd__mux2_1
X_11319_ fifo_bank_register.bank\[7\]\[4\] _05278_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15087_ addroundkey_data_o\[12\] _04378_ _05607_ _03358_ vssd1 vssd1 vccd1 vccd1
+ _03359_ sky130_fd_sc_hd__a211o_1
X_12299_ _05445_ fifo_bank_register.bank\[4\]\[83\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14038_ fifo_bank_register.bank\[1\]\[53\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[53\]
+ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15989_ ks1.key_reg\[5\] _03956_ _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__mux2_1
X_08530_ _04583_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17728_ net493 _01171_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08461_ _04547_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__dlymetal6s2s_1
X_17659_ net562 _01102_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08392_ addroundkey_data_o\[38\] fifo_bank_register.data_out\[38\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__mux2_2
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ mix1.data_o\[98\] _04698_ _04701_ _05034_ vssd1 vssd1 vccd1 vccd1 _05035_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold110 mix1.data_reg\[77\] vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 mix1.data_reg\[39\] vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold132 ks1.key_reg\[70\] vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold143 ks1.key_reg\[33\] vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 ks1.key_reg\[32\] vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 ks1.key_reg\[118\] vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 ks1.key_reg\[117\] vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout601 net602 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_229_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout612 net617 vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_2
X_09915_ _05757_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__buf_4
XFILLER_0_217_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout623 net625 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_4
Xfanout634 net635 vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_2
XFILLER_0_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout645 net646 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout667 net669 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__buf_2
X_09846_ _04640_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ net169 ks1.key_reg\[1\] _05625_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__mux2_2
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08728_ _04648_ _04719_ _04739_ _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a211o_2
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08659_ _04677_ _04678_ _04679_ _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a22o_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _07103_ vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__clkbuf_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10621_ sub1.data_o\[86\] _06393_ _06113_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13340_ _05401_ fifo_bank_register.bank\[0\]\[62\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10552_ _06090_ _05972_ sub1.data_o\[80\] _06079_ vssd1 vssd1 vccd1 vccd1 _06331_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13271_ _07948_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10483_ net227 ks1.key_reg\[72\] _06245_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15010_ mix1.data_reg\[66\] _03283_ _03171_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12222_ _07394_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _05299_ fifo_bank_register.bank\[4\]\[14\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ _06804_ vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__clkbuf_1
X_16961_ net437 _00404_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
X_12084_ _07221_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__buf_4
XFILLER_0_159_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15912_ sub1.data_o\[41\] _03576_ _03892_ sub1.data_o\[105\] vssd1 vssd1 vccd1 vccd1
+ _03894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11035_ _05249_ _05250_ net597 vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__or3b_1
XFILLER_0_95_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16892_ net570 _00335_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18631_ clknet_leaf_36_clk _02060_ net666 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_200_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15843_ mix1.data_o\[121\] net757 _03729_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__mux2_1
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18562_ clknet_leaf_63_clk _01991_ net598 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[89\]
+ sky130_fd_sc_hd__dfrtp_1
X_15774_ mix1.data_o\[88\] net761 _03808_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__mux2_1
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _07798_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17513_ net416 _00956_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_14725_ sub1.data_o\[55\] sub1.data_o\[119\] _05598_ vssd1 vssd1 vccd1 vccd1 _03026_
+ sky130_fd_sc_hd__mux2_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _07221_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__buf_4
X_18493_ clknet_leaf_54_clk _01922_ net615 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_185_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ net455 _00887_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11868_ _07207_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14656_ fifo_bank_register.bank\[6\]\[122\] _08104_ _08107_ fifo_bank_register.bank\[4\]\[122\]
+ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10819_ _05751_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__buf_4
X_13607_ fifo_bank_register.bank\[0\]\[7\] _08170_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17375_ net509 _00818_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14587_ _02909_ fifo_bank_register.data_out\[113\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02910_ sky130_fd_sc_hd__mux2_1
X_11799_ fifo_bank_register.bank\[6\]\[103\] _05487_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16326_ net674 _04136_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13538_ fifo_bank_register.bank\[6\]\[0\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13469_ _05530_ fifo_bank_register.bank\[0\]\[124\] _07914_ vssd1 vssd1 vccd1 vccd1
+ _08052_ sky130_fd_sc_hd__mux2_1
X_16257_ ks1.key_reg\[31\] _04200_ _04106_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15208_ _03297_ _03314_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16188_ _03901_ _04135_ _04137_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15139_ _05201_ _03406_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__nand2_4
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09700_ _05565_ vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ _05517_ vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09562_ fifo_bank_register.bank\[9\]\[95\] _05470_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08513_ _04574_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_195_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09493_ net228 vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08444_ _04538_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08375_ _04502_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout420 net427 vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__buf_2
Xfanout431 net436 vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_217_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__buf_2
XFILLER_0_100_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout453 net461 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout464 net466 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__clkbuf_2
Xfanout475 net476 vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_2
XFILLER_0_214_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout486 net489 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_2
X_09829_ _05679_ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__xor2_1
Xfanout497 net498 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12840_ fifo_bank_register.bank\[2\]\[82\] _05443_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07721_ sky130_fd_sc_hd__mux2_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _07684_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__clkbuf_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _07130_ vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__clkbuf_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ fifo_bank_register.bank\[9\]\[105\] _02793_ _02838_ _02839_ _02840_ vssd1
+ vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a2111o_1
X_15490_ sub1.data_o\[108\] _03600_ _03653_ sub1.data_o\[44\] vssd1 vssd1 vccd1 vccd1
+ _03658_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11653_ _07094_ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__clkbuf_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ fifo_bank_register.bank\[7\]\[98\] _02704_ _02713_ fifo_bank_register.bank\[2\]\[98\]
+ _02778_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__a221o_1
XFILLER_0_193_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10604_ _06377_ _06378_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17160_ net523 _00603_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
X_14372_ _02146_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ fifo_bank_register.bank\[6\]\[1\] _05272_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13323_ _05384_ fifo_bank_register.bank\[0\]\[54\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07976_ sky130_fd_sc_hd__mux2_1
X_16111_ net147 ks1.key_reg\[115\] _03976_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__mux2_2
XFILLER_0_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10535_ _06315_ vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17091_ net496 _00534_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13254_ _05315_ fifo_bank_register.bank\[0\]\[21\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16042_ _05195_ _04005_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__xor2_4
X_10466_ _06250_ _06252_ _06253_ _06254_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12205_ _07385_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13185_ _07902_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10397_ _06193_ vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__clkbuf_1
X_12136_ _05282_ fifo_bank_register.bank\[4\]\[6\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ net442 _01436_ net597 vssd1 vssd1 vccd1 vccd1 fifo_bank_register.read_ptr\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12067_ _07312_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__clkbuf_1
X_16944_ net463 _00387_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11018_ net30 mix1.data_o\[126\] _05603_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16875_ net417 _00318_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18614_ clknet_leaf_83_clk _02043_ net582 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[107\]
+ sky130_fd_sc_hd__dfrtp_1
X_15826_ _03845_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__clkbuf_1
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18545_ clknet_leaf_65_clk _01974_ net603 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[72\]
+ sky130_fd_sc_hd__dfrtp_1
X_15757_ _03809_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__clkbuf_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ fifo_bank_register.bank\[1\]\[15\] _05301_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14708_ _05104_ _04927_ _05554_ _03014_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a31o_1
XFILLER_0_158_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18476_ clknet_leaf_54_clk _01905_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_15688_ mix1.data_o\[47\] net768 _03764_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17427_ net552 _00870_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
X_14639_ fifo_bank_register.bank\[7\]\[120\] _08077_ _08092_ fifo_bank_register.bank\[2\]\[120\]
+ _02954_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17358_ net478 _00801_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16309_ net809 _04104_ _04222_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17289_ net522 _00732_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08993_ _05013_ _05015_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__xor2_4
XFILLER_0_167_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09614_ net144 vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__buf_2
XFILLER_0_218_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09545_ net247 vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09476_ _05412_ vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08427_ _04529_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_176_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08358_ _04493_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_149_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ net208 net210 net209 net207 vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__or4b_1
XFILLER_0_190_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10320_ net79 mix1.data_o\[55\] _06111_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10251_ _05899_ _06056_ _06060_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10182_ addroundkey_data_o\[41\] _05999_ _05980_ vssd1 vssd1 vccd1 vccd1 _06000_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14990_ _03260_ _03263_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__nor2_4
XFILLER_0_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13941_ fifo_bank_register.bank\[0\]\[42\] _02334_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16660_ net452 _00108_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13872_ fifo_bank_register.bank\[1\]\[35\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[35\]
+ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15611_ _03732_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12823_ fifo_bank_register.bank\[2\]\[74\] _05426_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07712_ sky130_fd_sc_hd__mux2_1
X_16591_ net437 _00039_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18330_ clknet_leaf_11_clk _01760_ net628 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15542_ _03690_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__clkbuf_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ fifo_bank_register.bank\[2\]\[41\] _05357_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07676_ sky130_fd_sc_hd__mux2_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ clknet_leaf_42_clk _01692_ net655 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _07121_ vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15473_ _03647_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__clkbuf_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ fifo_bank_register.bank\[2\]\[9\] _05288_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07639_ sky130_fd_sc_hd__mux2_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17212_ net469 _00655_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
X_11636_ _07085_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__clkbuf_1
X_14424_ fifo_bank_register.bank\[7\]\[96\] _02704_ _02713_ fifo_bank_register.bank\[2\]\[96\]
+ _02763_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__a221o_1
X_18192_ clknet_leaf_24_clk _01623_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17143_ net407 _00586_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14355_ _02702_ fifo_bank_register.data_out\[88\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02703_ sky130_fd_sc_hd__mux2_1
X_11567_ fifo_bank_register.bank\[7\]\[122\] _05526_ _06912_ vssd1 vssd1 vccd1 vccd1
+ _07048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13306_ _05367_ fifo_bank_register.bank\[0\]\[46\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07967_ sky130_fd_sc_hd__mux2_1
X_10518_ addroundkey_data_o\[76\] _06300_ _06248_ vssd1 vssd1 vccd1 vccd1 _06301_
+ sky130_fd_sc_hd__mux2_1
X_14286_ fifo_bank_register.bank\[1\]\[80\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[80\]
+ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a22o_1
X_17074_ net452 _00517_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ fifo_bank_register.bank\[7\]\[89\] _05457_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13237_ _07930_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__clkbuf_1
X_16025_ net193 ks1.key_reg\[41\] _03982_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__mux2_1
X_10449_ _05751_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__buf_4
XFILLER_0_62_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13168_ _07893_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12119_ fifo_bank_register.bank\[5\]\[127\] _05536_ _07198_ vssd1 vssd1 vccd1 vccd1
+ _07339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13099_ _07857_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__clkbuf_1
X_17976_ net457 _01419_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16927_ net548 _00370_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16858_ net501 _00301_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15809_ _03836_ vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16789_ clknet_leaf_36_clk _00233_ net649 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[80\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_172_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ fifo_bank_register.bank\[9\]\[20\] _05311_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18528_ clknet_leaf_60_clk _01957_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09261_ _05262_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18459_ clknet_leaf_27_clk _01889_ net642 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[99\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_145_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08212_ ks1.state\[2\] _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__nand2_4
XFILLER_0_44_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09192_ _05202_ _04367_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold14 mix1.data_reg\[122\] vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08976_ ks1.key_reg\[23\] _04735_ _04999_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a21oi_1
XTAP_4806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 ks1.key_reg\[13\] vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold36 mix1.data_reg\[127\] vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 mix1.data_reg\[102\] vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold58 mix1.data_reg\[103\] vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold69 mix1.data_reg\[96\] vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_224_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09528_ fifo_bank_register.bank\[9\]\[84\] _05447_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09459_ net216 vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__buf_2
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12470_ fifo_bank_register.bank\[3\]\[35\] _05344_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11421_ fifo_bank_register.bank\[7\]\[52\] _05380_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14140_ _02511_ fifo_bank_register.data_out\[64\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02512_ sky130_fd_sc_hd__mux2_1
X_11352_ _06911_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__buf_6
XFILLER_0_50_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10303_ _06107_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14071_ fifo_bank_register.bank\[9\]\[57\] _02388_ _02447_ _02448_ _02449_ vssd1
+ vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11283_ _05514_ fifo_bank_register.bank\[8\]\[116\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06898_ sky130_fd_sc_hd__mux2_1
X_13022_ _07794_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__buf_4
X_10234_ net71 mix1.data_o\[48\] _05934_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17830_ net445 _01273_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10165_ mix1.data_o\[40\] _05876_ _05821_ _05822_ sub1.data_o\[40\] vssd1 vssd1 vccd1
+ vccd1 _05984_ sky130_fd_sc_hd__a32o_1
XFILLER_0_218_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17761_ net486 _01204_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14973_ _03076_ _03246_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__xor2_4
X_10096_ net185 ks1.key_reg\[34\] _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__mux2_4
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16712_ clknet_leaf_51_clk _00156_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13924_ _02157_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__buf_4
X_17692_ net538 _01135_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16643_ net561 _00091_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
X_13855_ fifo_bank_register.bank\[6\]\[33\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[33\]
+ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ fifo_bank_register.bank\[2\]\[66\] _05409_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07703_ sky130_fd_sc_hd__mux2_1
X_16574_ net534 _00022_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_13786_ fifo_bank_register.bank\[5\]\[26\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[26\]
+ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a22o_1
X_10998_ net156 ks1.key_reg\[123\] _05762_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18313_ clknet_leaf_1_clk _01744_ net624 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[79\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15525_ sub1.data_o\[55\] _03663_ _03681_ _03673_ vssd1 vssd1 vccd1 vccd1 _03682_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ fifo_bank_register.bank\[2\]\[33\] _05340_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ clknet_leaf_10_clk _01675_ net625 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_15456_ _03635_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12668_ _07630_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14407_ fifo_bank_register.bank\[5\]\[94\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[94\]
+ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__a22o_1
X_18175_ clknet_leaf_12_clk _01606_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ fifo_bank_register.bank\[6\]\[18\] _05307_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07076_ sky130_fd_sc_hd__mux2_1
X_15387_ sub1.data_o\[7\] _03591_ _03581_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12599_ _07593_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17126_ net422 _00569_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14338_ _02687_ fifo_bank_register.data_out\[86\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17057_ net401 _00500_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14269_ fifo_bank_register.bank\[6\]\[79\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[79\]
+ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16008_ net713 _03901_ _03974_ _03975_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08830_ addroundkey_data_o\[14\] mix1.data_o\[14\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _04854_ sky130_fd_sc_hd__mux2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ addroundkey_data_o\[33\] mix1.data_o\[33\] _04656_ vssd1 vssd1 vccd1 vccd1
+ _04785_ sky130_fd_sc_hd__mux2_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ net455 _01402_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08692_ _04362_ _04363_ _04364_ _04365_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__nor4b_4
XFILLER_0_212_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ fifo_bank_register.bank\[9\]\[15\] _05301_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ net130 vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09175_ sbox1.alph\[1\] _05134_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_173_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput104 data_i[78] vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__buf_4
XTAP_5326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput115 data_i[88] vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_4
Xinput126 data_i[98] vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__clkbuf_4
XTAP_5337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput137 key_i[106] vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
XTAP_5359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput148 key_i[116] vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_4
Xinput159 key_i[126] vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_196_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08959_ addroundkey_data_o\[7\] mix1.data_o\[7\] _04663_ vssd1 vssd1 vccd1 vccd1
+ _04983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _07261_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__clkbuf_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10921_ _05623_ _06660_ _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__o21ai_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13640_ fifo_bank_register.bank\[1\]\[10\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _08201_ sky130_fd_sc_hd__a22o_1
X_10852_ net139 ks1.key_reg\[108\] _06579_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ fifo_bank_register.bank\[7\]\[3\] _08078_ _08093_ fifo_bank_register.bank\[2\]\[3\]
+ _08138_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__a221o_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ net132 ks1.key_reg\[101\] _06402_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__mux2_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clknet_3_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15310_ net791 _03402_ _03539_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12522_ _07508_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ net841 _04032_ _04206_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15241_ _03144_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_192_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12453_ fifo_bank_register.bank\[3\]\[27\] _05327_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11404_ fifo_bank_register.bank\[7\]\[44\] _05363_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15172_ _03090_ _03225_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__xor2_2
X_12384_ _05530_ fifo_bank_register.bank\[4\]\[124\] _07341_ vssd1 vssd1 vccd1 vccd1
+ _07479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14123_ fifo_bank_register.bank\[0\]\[62\] _02496_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11335_ _06926_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11266_ _05497_ fifo_bank_register.bank\[8\]\[108\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06889_ sky130_fd_sc_hd__mux2_1
X_14054_ fifo_bank_register.bank\[1\]\[55\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[55\]
+ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_197_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13005_ _07808_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__clkbuf_1
X_10217_ _06030_ vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11197_ _05428_ fifo_bank_register.bank\[8\]\[75\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17813_ net546 _01256_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10148_ _05968_ vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__clkbuf_1
XTAP_5860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ net503 _01187_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10079_ mix1.data_o\[33\] _05576_ _05758_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__o21a_1
X_14956_ addroundkey_data_o\[113\] _03056_ _03230_ vssd1 vssd1 vccd1 vccd1 _03231_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_221_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13907_ fifo_bank_register.bank\[9\]\[39\] _02226_ _02301_ _02302_ _02303_ vssd1
+ vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__a2111o_1
X_17675_ net516 _01118_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14887_ sub1.data_o\[127\] _03054_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16626_ net527 _00074_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13838_ fifo_bank_register.bank\[7\]\[31\] _02218_ _02227_ fifo_bank_register.bank\[2\]\[31\]
+ _02242_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a221o_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16557_ clknet_leaf_54_clk _00005_ net615 vssd1 vssd1 vccd1 vccd1 ks1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13769_ _02181_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_clk clknet_3_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15508_ sub1.data_o\[50\] _03663_ _03669_ _03611_ vssd1 vssd1 vccd1 vccd1 _03670_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16488_ _04327_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18227_ clknet_leaf_36_clk _01658_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15439_ sub1.data_o\[25\] _05553_ _04879_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18158_ clknet_leaf_49_clk _01589_ net616 vssd1 vssd1 vccd1 vccd1 ks1.col\[28\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17109_ net534 _00552_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18089_ net472 _01532_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09931_ net166 ks1.key_reg\[17\] _05762_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__mux2_2
XFILLER_0_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09862_ addroundkey_data_o\[10\] _05710_ _05697_ vssd1 vssd1 vccd1 vccd1 _05711_
+ sky130_fd_sc_hd__mux2_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08813_ _04661_ _04835_ _04836_ _04668_ vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__a22o_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ net191 ks1.key_reg\[3\] _05625_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ addroundkey_data_o\[97\] mix1.data_o\[97\] _04655_ vssd1 vssd1 vccd1 vccd1
+ _04768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ _04696_ _04697_ _04698_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__mux2_1
XANTENNA_209 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_193_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_187_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09227_ _05231_ _05232_ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_84_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09158_ _05165_ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_228_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09089_ sbox1.ah\[0\] _05074_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11120_ _06812_ vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11051_ _05282_ fifo_bank_register.bank\[8\]\[6\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10002_ addroundkey_data_o\[24\] _05836_ _05793_ vssd1 vssd1 vccd1 vccd1 _05837_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14810_ _05606_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__clkbuf_4
XTAP_5189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _03826_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__clkbuf_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _03034_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11953_ _07252_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10904_ net17 mix1.data_o\[114\] _05602_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__mux2_1
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17460_ net434 _00903_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ fifo_bank_register.bank\[6\]\[124\] _08104_ _08107_ fifo_bank_register.bank\[4\]\[124\]
+ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ fifo_bank_register.bank\[5\]\[15\] _05301_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16411_ _04285_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__clkbuf_1
X_13623_ fifo_bank_register.bank\[6\]\[9\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10835_ _06583_ _06585_ _06586_ _06587_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__a22o_1
X_17391_ net398 _00834_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_24_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16342_ _04246_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__clkbuf_1
X_13554_ fifo_bank_register.bank\[5\]\[1\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[1\]
+ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ sub1.data_o\[100\] _06524_ _06478_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12505_ _07544_ vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__clkbuf_1
X_16273_ _04209_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10697_ sub1.data_o\[94\] _06461_ _06318_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__mux2_1
X_13485_ _08063_ vssd1 vssd1 vccd1 vccd1 _08064_ sky130_fd_sc_hd__buf_4
X_18012_ net534 _01455_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15224_ net731 _03484_ _03425_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12436_ _07507_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15155_ _05201_ _03421_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__nand2_2
X_12367_ _07470_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14106_ _02157_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__buf_4
XFILLER_0_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _06917_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__clkbuf_1
X_15086_ addroundkey_data_o\[76\] _03072_ _03068_ addroundkey_data_o\[44\] vssd1 vssd1
+ vccd1 vccd1 _03358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12298_ _07434_ vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14037_ fifo_bank_register.bank\[6\]\[53\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[53\]
+ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a22o_1
X_11249_ _06791_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15988_ _03957_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__buf_4
XFILLER_0_222_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17727_ net491 _01170_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
X_14939_ addroundkey_data_o\[0\] _03208_ _03086_ _03213_ vssd1 vssd1 vccd1 vccd1 _03214_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08460_ addroundkey_data_o\[70\] fifo_bank_register.data_out\[70\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__mux2_1
X_17658_ net563 _01101_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16609_ net407 _00057_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_08391_ _04510_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_148_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17589_ net409 _01032_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ addroundkey_data_o\[98\] _04778_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 mix1.data_reg\[73\] vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold111 mix1.data_reg\[104\] vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 mix1.data_reg\[86\] vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold133 ks1.key_reg\[84\] vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 ks1.key_reg\[113\] vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 ks1.key_reg\[36\] vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 ks1.key_reg\[67\] vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 ks1.key_reg\[68\] vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09914_ _05616_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__buf_8
XFILLER_0_10_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout602 net618 vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__buf_4
Xfanout613 net614 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__buf_4
Xfanout624 net626 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__clkbuf_4
Xfanout635 net670 vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout646 net650 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_2
XFILLER_0_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09845_ _05693_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__xor2_1
Xfanout657 net660 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__clkbuf_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout668 net669 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09776_ _05629_ _05631_ _05632_ _05633_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__a22o_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _04741_ _04744_ _04748_ _04750_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_217_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _04680_ _04681_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__nor2_2
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08589_ net129 vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__inv_4
XFILLER_0_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10620_ net113 mix1.data_o\[86\] _06111_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10551_ sub1.data_o\[80\] _06329_ _06113_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10482_ _06250_ _06267_ _06268_ _06254_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__a22o_1
X_13270_ _05331_ fifo_bank_register.bank\[0\]\[29\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ _05367_ fifo_bank_register.bank\[4\]\[46\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12152_ _07357_ vssd1 vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11103_ _05333_ fifo_bank_register.bank\[8\]\[30\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16960_ net491 _00403_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
X_12083_ _07320_ vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15911_ _03717_ _04943_ _05548_ _03893_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__a31o_1
X_11034_ _05266_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__inv_2
XFILLER_0_198_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16891_ net563 _00334_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18630_ clknet_leaf_36_clk _02059_ net666 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_194_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15842_ _03853_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__clkbuf_1
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18561_ clknet_leaf_65_clk _01990_ net604 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[88\]
+ sky130_fd_sc_hd__dfrtp_1
X_15773_ _03817_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__clkbuf_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ fifo_bank_register.bank\[1\]\[22\] _05317_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07798_ sky130_fd_sc_hd__mux2_1
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ net418 _00955_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14724_ _03019_ _04927_ _05236_ _03025_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__a31o_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11936_ _07243_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__clkbuf_1
X_18492_ clknet_leaf_54_clk _01921_ net614 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_169_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17443_ net400 _00886_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14655_ fifo_bank_register.bank\[7\]\[122\] _08077_ _08092_ fifo_bank_register.bank\[2\]\[122\]
+ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__a221o_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11867_ fifo_bank_register.bank\[5\]\[7\] _05284_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ fifo_bank_register.bank\[9\]\[7\] _08090_ _08167_ _08168_ _08169_ vssd1 vssd1
+ vccd1 vccd1 _08170_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10818_ net7 mix1.data_o\[105\] _06571_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__mux2_1
X_17374_ net485 _00817_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14586_ fifo_bank_register.bank\[0\]\[113\] _02908_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11798_ _07170_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16325_ _04237_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13537_ _08107_ vssd1 vssd1 vccd1 vccd1 _08108_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_171_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10749_ addroundkey_data_o\[98\] _06509_ _06431_ vssd1 vssd1 vccd1 vccd1 _06510_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16256_ _05002_ _04199_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13468_ _08051_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15207_ _03107_ _03404_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__xor2_4
XFILLER_0_140_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12419_ fifo_bank_register.bank\[3\]\[11\] _05293_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07499_ sky130_fd_sc_hd__mux2_1
X_16187_ net712 _04136_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13399_ _05459_ fifo_bank_register.bank\[0\]\[90\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15138_ _03390_ _03405_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15069_ addroundkey_data_o\[20\] _04379_ _05607_ _03340_ vssd1 vssd1 vccd1 vccd1
+ _03341_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_4_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09630_ fifo_bank_register.bank\[9\]\[117\] _05516_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09561_ net252 vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08512_ addroundkey_data_o\[95\] fifo_bank_register.data_out\[95\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09492_ _05423_ vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08443_ addroundkey_data_o\[62\] fifo_bank_register.data_out\[62\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08374_ addroundkey_data_o\[29\] fifo_bank_register.data_out\[29\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout410 net413 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout421 net422 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__buf_1
Xfanout432 net436 vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_2
Xfanout443 net444 vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__buf_2
XFILLER_0_217_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout454 net460 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_2
XFILLER_0_219_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout465 net466 vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_2
Xfanout476 net481 vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_2
Xfanout487 net489 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__buf_2
X_09828_ net235 ks1.key_reg\[7\] _05625_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__mux2_1
Xfanout498 net530 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__buf_2
XFILLER_0_119_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09759_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__clkbuf_4
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ fifo_bank_register.bank\[2\]\[49\] _05373_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ fifo_bank_register.bank\[6\]\[66\] _05409_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14440_ fifo_bank_register.bank\[5\]\[98\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[98\]
+ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__a22o_1
X_11652_ fifo_bank_register.bank\[6\]\[33\] _05340_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07094_ sky130_fd_sc_hd__mux2_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ net240 ks1.key_reg\[84\] _06097_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14371_ fifo_bank_register.bank\[7\]\[90\] _02704_ _02713_ fifo_bank_register.bank\[2\]\[90\]
+ _02716_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11583_ _07057_ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16110_ _04066_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__clkbuf_1
X_13322_ _07975_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17090_ net494 _00533_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
X_10534_ addroundkey_data_o\[78\] _06314_ _06248_ vssd1 vssd1 vccd1 vccd1 _06315_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16041_ net138 ks1.key_reg\[107\] _03902_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__mux2_2
XFILLER_0_161_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10465_ _04609_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__clkbuf_4
X_13253_ _07939_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ _05350_ fifo_bank_register.bank\[4\]\[38\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10396_ addroundkey_data_o\[62\] _06192_ _06169_ vssd1 vssd1 vccd1 vccd1 _06193_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13184_ fifo_bank_register.bank\[1\]\[117\] _05516_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12135_ _07348_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17992_ net437 _01435_ net597 vssd1 vssd1 vccd1 vccd1 fifo_bank_register.read_ptr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16943_ net468 _00386_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
X_12066_ fifo_bank_register.bank\[5\]\[101\] _05483_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11017_ _06750_ vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__clkbuf_1
X_16874_ net423 _00317_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_159_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15825_ mix1.data_o\[112\] net771 _03841_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__mux2_1
X_18613_ clknet_leaf_84_clk _02042_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15756_ mix1.data_o\[79\] net731 _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__mux2_1
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18544_ clknet_leaf_63_clk _01973_ net599 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[71\]
+ sky130_fd_sc_hd__dfrtp_1
X_12968_ _07788_ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ sub1.data_o\[81\] _03010_ _03013_ sub1.next_ready_o vssd1 vssd1 vccd1 vccd1
+ _03014_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11919_ fifo_bank_register.bank\[5\]\[31\] _05336_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18475_ clknet_leaf_58_clk _01904_ net602 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15687_ _03772_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12899_ fifo_bank_register.bank\[2\]\[110\] _05501_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07752_ sky130_fd_sc_hd__mux2_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ net545 _00869_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14638_ fifo_bank_register.bank\[5\]\[120\] _08096_ _08099_ fifo_bank_register.bank\[3\]\[120\]
+ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a22o_1
XFILLER_0_185_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ net477 _00800_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14569_ fifo_bank_register.bank\[9\]\[111\] _02874_ _02891_ _02892_ _02893_ vssd1
+ vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16308_ _04228_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__clkbuf_1
X_17288_ net522 _00731_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16239_ net159 ks1.key_reg\[126\] _03976_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__mux2_2
XFILLER_0_207_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08992_ _04794_ _05014_ _04874_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__mux2_4
XFILLER_0_103_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09613_ _05505_ vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09544_ _05458_ vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09475_ fifo_bank_register.bank\[9\]\[67\] _05411_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08426_ addroundkey_data_o\[54\] fifo_bank_register.data_out\[54\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__mux2_4
XFILLER_0_136_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08357_ addroundkey_data_o\[21\] fifo_bank_register.data_out\[21\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08288_ net212 net211 net215 net214 vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_85_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10250_ sub1.data_o\[49\] _05971_ _06058_ _06059_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _06060_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10181_ _05996_ _05998_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13940_ fifo_bank_register.bank\[9\]\[42\] _02307_ _02331_ _02332_ _02333_ vssd1
+ vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_227_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13871_ fifo_bank_register.bank\[6\]\[35\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[35\]
+ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15610_ mix1.data_o\[10\] _03435_ _03730_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12822_ _07711_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16590_ net437 _00038_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15541_ sub1.data_o\[63\] _05244_ _04884_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__mux2_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12753_ _07675_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18260_ clknet_leaf_51_clk _01691_ net655 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ fifo_bank_register.bank\[6\]\[58\] _05392_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15472_ sub1.data_o\[37\] _03646_ _03636_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _07638_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ net435 _00654_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14423_ fifo_bank_register.bank\[5\]\[96\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[96\]
+ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a22o_1
X_18191_ clknet_leaf_24_clk _01622_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11635_ fifo_bank_register.bank\[6\]\[25\] _05323_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17142_ net395 _00585_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_14354_ fifo_bank_register.bank\[0\]\[88\] _02701_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02702_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11566_ _07047_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13305_ _07966_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10517_ _06298_ _06299_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__xor2_1
X_17073_ net462 _00516_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14285_ _02153_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11497_ _07011_ vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__clkbuf_1
X_16024_ _03987_ _03989_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__xnor2_2
X_13236_ _05297_ fifo_bank_register.bank\[0\]\[13\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10448_ net94 mix1.data_o\[69\] _06237_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ fifo_bank_register.bank\[1\]\[109\] _05499_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07893_ sky130_fd_sc_hd__mux2_1
X_10379_ _06176_ _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ _07338_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__clkbuf_1
X_13098_ fifo_bank_register.bank\[1\]\[76\] _05430_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07857_ sky130_fd_sc_hd__mux2_1
X_17975_ net469 _01418_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16926_ net566 _00369_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
X_12049_ fifo_bank_register.bank\[5\]\[93\] _05466_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16857_ net505 _00300_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15808_ mix1.data_o\[104\] net781 _03830_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16788_ clknet_3_1__leaf_clk _00232_ net594 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[79\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_220_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15739_ mix1.data_o\[71\] net720 _03797_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18527_ clknet_leaf_60_clk _01956_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09260_ _05263_ fifo_bank_register.write_ptr\[3\] _05251_ vssd1 vssd1 vccd1 vccd1
+ _05264_ sky130_fd_sc_hd__mux2_1
X_18458_ clknet_leaf_32_clk _01888_ net653 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[98\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08211_ ks1.state\[1\] ks1.state\[0\] vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__nor2_1
X_09191_ _05201_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__buf_4
XFILLER_0_172_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17409_ net573 _00852_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_18389_ clknet_leaf_0_clk _01819_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[74\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08975_ ks1.key_reg\[23\] _04745_ _04746_ net173 vssd1 vssd1 vccd1 vccd1 _04999_
+ sky130_fd_sc_hd__o31a_1
Xhold15 ks1.key_reg\[79\] vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_228_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold26 mix1.data_reg\[115\] vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold37 ks1.key_reg\[11\] vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold48 mix1.data_reg\[45\] vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 mix1.data_reg\[125\] vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09527_ net240 vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_196_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _05400_ vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__clkbuf_1
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ addroundkey_data_o\[46\] fifo_bank_register.data_out\[46\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__mux2_2
XFILLER_0_164_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09389_ _05353_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11420_ _06971_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ _06934_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10302_ net206 ks1.key_reg\[53\] _06097_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__mux2_4
X_14070_ fifo_bank_register.bank\[1\]\[57\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[57\]
+ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11282_ _06897_ vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__clkbuf_1
X_13021_ _07816_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10233_ _06044_ vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10164_ sub1.data_o\[40\] _05982_ _05819_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14972_ _03187_ _03245_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__xnor2_4
X_17760_ net483 _01203_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_10095_ _05707_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__buf_4
XFILLER_0_195_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16711_ clknet_leaf_51_clk _00155_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_13923_ fifo_bank_register.bank\[9\]\[40\] _02307_ _02312_ _02315_ _02318_ vssd1
+ vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__a2111o_1
X_17691_ net540 _01134_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16642_ net560 _00090_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13854_ fifo_bank_register.bank\[7\]\[33\] _02218_ _02227_ fifo_bank_register.bank\[2\]\[33\]
+ _02256_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__a221o_1
XFILLER_0_202_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12805_ _07702_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16573_ net505 _00021_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13785_ _02195_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__clkbuf_1
X_10997_ _06583_ _06731_ _06732_ _06587_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15524_ sub1.data_o\[23\] sub1.data_o\[87\] _03671_ vssd1 vssd1 vccd1 vccd1 _03681_
+ sky130_fd_sc_hd__mux2_1
X_18312_ clknet_leaf_1_clk _01743_ net624 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[78\]
+ sky130_fd_sc_hd__dfrtp_4
X_12736_ _07666_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__clkbuf_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ clknet_leaf_2_clk _01674_ net623 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15455_ _04368_ _04675_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12667_ fifo_bank_register.bank\[2\]\[0\] _05248_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14406_ _02748_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18174_ clknet_leaf_20_clk _01605_ net640 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ _07075_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__clkbuf_1
X_15386_ sub1.data_o\[39\] sub1.data_o\[103\] _05202_ vssd1 vssd1 vccd1 vccd1 _03591_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ fifo_bank_register.bank\[3\]\[96\] _05472_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17125_ net437 _00568_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14337_ fifo_bank_register.bank\[0\]\[86\] _02686_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11549_ fifo_bank_register.bank\[7\]\[113\] _05508_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17056_ net409 _00499_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
X_14268_ fifo_bank_register.bank\[7\]\[79\] _02623_ _02551_ fifo_bank_register.bank\[2\]\[79\]
+ _02624_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16007_ _05007_ _03973_ _03914_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ _05280_ fifo_bank_register.bank\[0\]\[5\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07921_ sky130_fd_sc_hd__mux2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14199_ _02564_ fifo_bank_register.data_out\[70\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02565_ sky130_fd_sc_hd__mux2_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08760_ _04695_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__clkbuf_4
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ net403 _01401_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16909_ net525 _00352_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08691_ addroundkey_data_o\[92\] mix1.data_o\[92\] _04666_ vssd1 vssd1 vccd1 vccd1
+ _04715_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17889_ net480 _01332_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09312_ net164 vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09243_ _04741_ _04755_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09174_ _05120_ _05121_ sbox1.alph\[2\] vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput105 data_i[79] vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_2
XTAP_5316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput116 data_i[89] vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput127 data_i[99] vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_4
XFILLER_0_216_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput138 key_i[107] vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__buf_4
X_08958_ addroundkey_data_o\[63\] mix1.data_o\[63\] _04778_ vssd1 vssd1 vccd1 vccd1
+ _04982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput149 key_i[117] vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_4
XTAP_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ ks1.key_reg\[8\] _04726_ _04912_ net246 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10920_ sub1.data_o\[115\] _06513_ _06662_ _06663_ _04610_ vssd1 vssd1 vccd1 vccd1
+ _06664_ sky130_fd_sc_hd__a221o_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _06583_ _06600_ _06601_ _06587_ vssd1 vssd1 vccd1 vccd1 _06602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ fifo_bank_register.bank\[5\]\[3\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[3\]
+ vssd1 vssd1 vccd1 vccd1 _08138_ sky130_fd_sc_hd__a22o_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _06381_ _06535_ _06539_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__o21ai_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _07552_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _03495_ _03496_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12452_ _07516_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11403_ _06962_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__clkbuf_1
X_15171_ _03436_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__clkbuf_1
X_12383_ _07478_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14122_ fifo_bank_register.bank\[9\]\[62\] _02469_ _02493_ _02494_ _02495_ vssd1
+ vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__a2111o_1
X_11334_ fifo_bank_register.bank\[7\]\[11\] _05293_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14053_ fifo_bank_register.bank\[6\]\[55\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[55\]
+ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a22o_1
X_11265_ _06888_ vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13004_ fifo_bank_register.bank\[1\]\[31\] _05336_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07808_ sky130_fd_sc_hd__mux2_1
X_10216_ addroundkey_data_o\[45\] _06029_ _05980_ vssd1 vssd1 vccd1 vccd1 _06030_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11196_ _06852_ vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17812_ net525 _01255_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10147_ addroundkey_data_o\[38\] _05967_ _05872_ vssd1 vssd1 vccd1 vccd1 _05968_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14955_ addroundkey_data_o\[17\] _04377_ _03086_ _03229_ vssd1 vssd1 vccd1 vccd1
+ _03230_ sky130_fd_sc_hd__a211o_1
X_17743_ net478 _01186_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_10078_ _05575_ _05901_ _05903_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__a21o_1
XTAP_5894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13906_ fifo_bank_register.bank\[1\]\[39\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[39\]
+ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14886_ sub1.data_o\[31\] _04374_ _04658_ _03161_ vssd1 vssd1 vccd1 vccd1 _03162_
+ sky130_fd_sc_hd__a211o_1
X_17674_ net521 _01117_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13837_ fifo_bank_register.bank\[5\]\[31\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__a22o_1
X_16625_ net526 _00073_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16556_ clknet_leaf_28_clk _00004_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[119\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13768_ _02180_ fifo_bank_register.data_out\[23\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15507_ sub1.data_o\[18\] sub1.data_o\[82\] _03609_ vssd1 vssd1 vccd1 vccd1 _03669_
+ sky130_fd_sc_hd__mux2_1
X_12719_ _07657_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__clkbuf_1
X_16487_ net784 _03382_ _04321_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13699_ fifo_bank_register.bank\[0\]\[17\] _02117_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_216_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18226_ clknet_leaf_37_clk _01657_ net666 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[56\]
+ sky130_fd_sc_hd__dfrtp_1
X_15438_ _03625_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15369_ _03579_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18157_ clknet_leaf_67_clk _01588_ net606 vssd1 vssd1 vccd1 vccd1 ks1.col\[27\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_142_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17108_ net534 _00551_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_18088_ net405 _01531_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[90\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09930_ _05568_ _05767_ _05771_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17039_ net545 _00482_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09861_ _05706_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__xor2_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08812_ addroundkey_data_o\[78\] mix1.data_o\[78\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _04836_ sky130_fd_sc_hd__mux2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _05629_ _05646_ _05647_ _05633_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a22o_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08743_ addroundkey_data_o\[113\] mix1.data_o\[113\] _04655_ vssd1 vssd1 vccd1 vccd1
+ _04767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _04650_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__clkbuf_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_191_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09226_ _04649_ _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09157_ _05166_ _05167_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _05094_ _05099_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__xnor2_1
X_11050_ _06775_ vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10001_ _05834_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__xor2_1
XTAP_5124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ ks1.col\[6\] _05235_ _04916_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__mux2_1
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ fifo_bank_register.bank\[5\]\[47\] _05369_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ _06648_ vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__clkbuf_1
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ fifo_bank_register.bank\[7\]\[124\] _08077_ _08092_ fifo_bank_register.bank\[2\]\[124\]
+ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a221o_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _07215_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16410_ ks1.key_reg\[100\] _03943_ _04281_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13622_ fifo_bank_register.bank\[7\]\[9\] _08182_ _08093_ fifo_bank_register.bank\[2\]\[9\]
+ _08183_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10834_ _04609_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__clkbuf_4
X_17390_ net395 _00833_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16341_ net802 _03963_ _04240_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__mux2_1
X_13553_ _08123_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__clkbuf_1
X_10765_ net2 mix1.data_o\[100\] _06476_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12504_ fifo_bank_register.bank\[3\]\[51\] _05378_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16272_ ks1.key_reg\[38\] _03965_ _04206_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13484_ _05258_ _08062_ _04466_ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__o21ai_4
X_10696_ net122 mix1.data_o\[94\] _06316_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15223_ _03482_ _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18011_ net506 _01454_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[13\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_202_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ fifo_bank_register.bank\[3\]\[19\] _05309_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15154_ _03406_ _03420_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__xor2_2
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12366_ _05512_ fifo_bank_register.bank\[4\]\[115\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14105_ fifo_bank_register.bank\[9\]\[60\] _02469_ _02474_ _02477_ _02480_ vssd1
+ vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__a2111o_1
X_11317_ fifo_bank_register.bank\[7\]\[3\] _05276_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15085_ sub1.data_o\[108\] _03057_ _03356_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12297_ _05443_ fifo_bank_register.bank\[4\]\[82\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14036_ fifo_bank_register.bank\[7\]\[53\] _02380_ _02389_ fifo_bank_register.bank\[2\]\[53\]
+ _02418_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__a221o_1
XFILLER_0_226_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11248_ _06879_ vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11179_ _06843_ vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15987_ _04372_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__buf_4
XTAP_5691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17726_ net441 _01169_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
X_14938_ addroundkey_data_o\[64\] _03209_ _03067_ addroundkey_data_o\[32\] vssd1 vssd1
+ vccd1 vccd1 _03213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17657_ net573 _01100_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_14869_ _03068_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__buf_6
XFILLER_0_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16608_ net395 _00056_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08390_ addroundkey_data_o\[37\] fifo_bank_register.data_out\[37\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__mux2_2
XFILLER_0_147_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17588_ net432 _01031_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16539_ net765 _03533_ _03143_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09011_ _05031_ _05032_ _04650_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18209_ clknet_leaf_15_clk _01640_ net629 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 mix1.data_reg\[112\] vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 mix1.data_reg\[92\] vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 ks1.key_reg\[115\] vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 ks1.key_reg\[102\] vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold145 ks1.key_reg\[122\] vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 ks1.key_reg\[103\] vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 ks1.key_reg\[80\] vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_229_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09913_ _05575_ _05752_ _05755_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__a21o_1
Xhold178 ks1.key_reg\[89\] vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 net607 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout614 net617 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_2
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout636 net638 vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__clkbuf_4
Xfanout647 net648 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__clkbuf_4
X_09844_ net257 ks1.key_reg\[9\] _05625_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__mux2_2
XFILLER_0_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__buf_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout669 net670 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_4
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _05567_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08726_ _04723_ _04749_ _04720_ _04370_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__o211a_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08657_ sub1.state\[3\] sub1.state\[2\] vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__or2_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _04613_ round\[2\] round\[3\] round\[1\] vssd1 vssd1 vccd1 vccd1 _04616_
+ sky130_fd_sc_hd__and4bb_2
XFILLER_0_165_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10550_ net107 mix1.data_o\[80\] _06111_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09209_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10481_ mix1.data_o\[72\] _06217_ _06241_ _06242_ sub1.data_o\[72\] vssd1 vssd1 vccd1
+ vccd1 _06268_ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12220_ _07393_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ _05297_ fifo_bank_register.bank\[4\]\[13\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11102_ _06791_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__buf_4
XFILLER_0_208_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12082_ fifo_bank_register.bank\[5\]\[109\] _05499_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15910_ sub1.data_o\[40\] _03576_ _03892_ sub1.data_o\[104\] vssd1 vssd1 vccd1 vccd1
+ _03893_ sky130_fd_sc_hd__a22o_1
X_11033_ _06764_ vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16890_ net562 _00333_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15841_ mix1.data_o\[120\] net744 _03729_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__mux2_1
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18560_ clknet_leaf_64_clk _01989_ net603 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[87\]
+ sky130_fd_sc_hd__dfrtp_1
X_15772_ mix1.data_o\[87\] net747 _03808_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__mux2_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _07797_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__clkbuf_1
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ net424 _00954_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_14723_ sub1.data_o\[86\] _03010_ _03024_ sub1.next_ready_o vssd1 vssd1 vccd1 vccd1
+ _03025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11935_ fifo_bank_register.bank\[5\]\[39\] _05352_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ clknet_leaf_55_clk _01920_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14654_ fifo_bank_register.bank\[5\]\[122\] _08096_ _08099_ fifo_bank_register.bank\[3\]\[122\]
+ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__a22o_1
X_17442_ net410 _00885_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11866_ _07206_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__clkbuf_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13605_ fifo_bank_register.bank\[1\]\[7\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10817_ _05749_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17373_ net484 _00816_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14585_ fifo_bank_register.bank\[9\]\[113\] _02874_ _02905_ _02906_ _02907_ vssd1
+ vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11797_ fifo_bank_register.bank\[6\]\[102\] _05485_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13536_ _08106_ vssd1 vssd1 vccd1 vccd1 _08107_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16324_ ks1.key_reg\[62\] _04236_ _04222_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__mux2_1
X_10748_ _06507_ _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16255_ _04197_ _04198_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__xor2_2
X_13467_ _05528_ fifo_bank_register.bank\[0\]\[123\] _07914_ vssd1 vssd1 vccd1 vccd1
+ _08051_ sky130_fd_sc_hd__mux2_1
X_10679_ _06446_ vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15206_ _03468_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12418_ _07498_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__clkbuf_1
X_16186_ _04371_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13398_ _07937_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__buf_4
X_15137_ _03380_ _03404_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__xor2_4
XFILLER_0_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12349_ _05495_ fifo_bank_register.bank\[4\]\[107\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07461_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ addroundkey_data_o\[84\] _03072_ _03068_ addroundkey_data_o\[52\] vssd1 vssd1
+ vccd1 vccd1 _03340_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14019_ fifo_bank_register.bank\[5\]\[51\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[51\]
+ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09560_ _05469_ vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08511_ _04573_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17709_ net453 _01152_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
X_09491_ fifo_bank_register.bank\[9\]\[72\] _05422_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08442_ _04537_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08373_ _04478_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__buf_8
XFILLER_0_163_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout400 net404 vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__buf_2
XFILLER_0_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout422 net427 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__buf_2
XFILLER_0_10_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout433 net436 vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__buf_1
Xfanout444 fifo_bank_register.clk vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 net460 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout466 net472 vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__buf_2
X_09827_ _05629_ _05674_ _05678_ _05633_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__a22o_1
Xfanout477 net481 vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__buf_2
XFILLER_0_214_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_225_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout499 net507 vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_2
XFILLER_0_216_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09758_ _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__buf_4
XFILLER_0_198_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ ks1.key_reg\[4\] _04730_ _04732_ net202 vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__o31a_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _05558_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__buf_6
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _07129_ vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__clkbuf_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11651_ _07093_ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10602_ _06076_ _06372_ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14370_ fifo_bank_register.bank\[5\]\[90\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[90\]
+ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11582_ fifo_bank_register.bank\[6\]\[0\] _05248_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ _05382_ fifo_bank_register.bank\[0\]\[53\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07975_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10533_ _06312_ _06313_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ net230 ks1.key_reg\[75\] _03918_ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ _05311_ fifo_bank_register.bank\[0\]\[20\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07939_ sky130_fd_sc_hd__mux2_1
X_10464_ mix1.data_o\[70\] _06217_ _06241_ _06242_ sub1.data_o\[70\] vssd1 vssd1 vccd1
+ vccd1 _06253_ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ _07384_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13183_ _07901_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__clkbuf_1
X_10395_ _06190_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _05280_ fifo_bank_register.bank\[4\]\[5\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17991_ net438 _01434_ net597 vssd1 vssd1 vccd1 vccd1 fifo_bank_register.read_ptr\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12065_ _07311_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__clkbuf_1
X_16942_ net463 _00385_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11016_ addroundkey_data_o\[125\] _06749_ _05696_ vssd1 vssd1 vccd1 vccd1 _06750_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16873_ net428 _00316_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18612_ clknet_leaf_12_clk _02041_ net628 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ _03844_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__clkbuf_1
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18543_ clknet_leaf_79_clk _01972_ net579 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[70\]
+ sky130_fd_sc_hd__dfrtp_1
X_15755_ _03741_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__buf_4
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ fifo_bank_register.bank\[1\]\[14\] _05299_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14706_ sub1.data_o\[49\] sub1.data_o\[113\] _05598_ vssd1 vssd1 vccd1 vccd1 _03013_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _07234_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__clkbuf_1
X_18474_ clknet_leaf_56_clk _01903_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_197_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15686_ mix1.data_o\[46\] net730 _03764_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__mux2_1
X_12898_ _07651_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__clkbuf_4
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17425_ net552 _00868_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
X_14637_ _02953_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__clkbuf_1
X_11849_ _07196_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17356_ net477 _00799_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14568_ fifo_bank_register.bank\[1\]\[111\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[111\]
+ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16307_ net821 _04096_ _04222_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13519_ _08089_ vssd1 vssd1 vccd1 vccd1 _08090_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17287_ net521 _00730_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14499_ fifo_bank_register.bank\[7\]\[104\] _02785_ _02794_ fifo_bank_register.bank\[2\]\[104\]
+ _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__a221o_1
X_16238_ ks1.col\[30\] _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16169_ net209 ks1.key_reg\[56\] _03982_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08991_ _04873_ _04923_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09612_ fifo_bank_register.bank\[9\]\[111\] _05504_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09543_ fifo_bank_register.bank\[9\]\[89\] _05457_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09474_ net221 vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__buf_2
XFILLER_0_176_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08425_ _04528_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__buf_1
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08356_ _04492_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08287_ _04438_ _04441_ _04442_ _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__or4_2
XFILLER_0_190_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10180_ net193 ks1.key_reg\[41\] _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ fifo_bank_register.bank\[7\]\[35\] _02218_ _02227_ fifo_bank_register.bank\[2\]\[35\]
+ _02270_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12821_ fifo_bank_register.bank\[2\]\[73\] _05424_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15540_ _03689_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__clkbuf_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ fifo_bank_register.bank\[2\]\[40\] _05354_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07675_ sky130_fd_sc_hd__mux2_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11703_ _07120_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__clkbuf_1
X_15471_ sub1.data_o\[69\] _05227_ _03633_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__mux2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ fifo_bank_register.bank\[2\]\[8\] _05286_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _02762_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__clkbuf_1
X_17210_ net411 _00653_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
X_11634_ _07084_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18190_ clknet_leaf_24_clk _01621_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[84\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14353_ fifo_bank_register.bank\[9\]\[88\] _02631_ _02698_ _02699_ _02700_ vssd1
+ vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__a2111o_1
X_17141_ net396 _00584_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11565_ fifo_bank_register.bank\[7\]\[121\] _05524_ _06912_ vssd1 vssd1 vccd1 vccd1
+ _07047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _05365_ fifo_bank_register.bank\[0\]\[45\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10516_ net231 ks1.key_reg\[76\] _06245_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__mux2_1
X_17072_ net464 _00515_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
X_14284_ _02151_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__clkbuf_4
X_11496_ fifo_bank_register.bank\[7\]\[88\] _05455_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13235_ _07929_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__clkbuf_1
X_16023_ _05553_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__xnor2_2
X_10447_ _05749_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13166_ _07892_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__clkbuf_1
X_10378_ net214 ks1.key_reg\[60\] _06166_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__mux2_1
X_12117_ fifo_bank_register.bank\[5\]\[126\] _05534_ _07198_ vssd1 vssd1 vccd1 vccd1
+ _07338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17974_ net433 _01417_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
X_13097_ _07856_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ _07302_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__clkbuf_1
X_16925_ net561 _00368_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16856_ net532 _00299_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15807_ _03835_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16787_ clknet_leaf_80_clk _00231_ net579 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[78\]
+ sky130_fd_sc_hd__dfrtp_4
X_13999_ fifo_bank_register.bank\[0\]\[49\] _02385_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18526_ clknet_leaf_66_clk _01955_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15738_ _03799_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18457_ clknet_leaf_30_clk _01887_ net642 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[97\]
+ sky130_fd_sc_hd__dfrtp_4
X_15669_ mix1.data_o\[38\] net762 _03753_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_190 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08210_ _04369_ vssd1 vssd1 vccd1 vccd1 sub1.next_ready_o sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17408_ net558 _00851_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_09190_ _04624_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__buf_4
XFILLER_0_111_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18388_ clknet_leaf_12_clk _01818_ net622 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[73\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17339_ net434 _00782_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08974_ _04653_ _04972_ _04985_ _04997_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__a211o_1
Xhold16 ks1.key_reg\[109\] vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold27 mix1.data_reg\[70\] vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 ks1.key_reg\[10\] vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold49 mix1.data_reg\[99\] vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ _05446_ vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09457_ fifo_bank_register.bank\[9\]\[61\] _05399_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08408_ _04519_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09388_ fifo_bank_register.bank\[9\]\[39\] _05352_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08339_ _04483_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11350_ fifo_bank_register.bank\[7\]\[19\] _05309_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10301_ _06076_ _06102_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_160_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11281_ _05512_ fifo_bank_register.bank\[8\]\[115\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13020_ fifo_bank_register.bank\[1\]\[39\] _05352_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07816_ sky130_fd_sc_hd__mux2_1
X_10232_ addroundkey_data_o\[47\] _06043_ _05980_ vssd1 vssd1 vccd1 vccd1 _06044_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10163_ net63 mix1.data_o\[40\] _05817_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10094_ _05899_ _05912_ _05918_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__o21ai_2
X_14971_ _03241_ _03244_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__nor2_8
X_16710_ clknet_leaf_41_clk _00154_ net658 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13922_ fifo_bank_register.bank\[1\]\[40\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[40\]
+ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17690_ net536 _01133_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ net563 _00089_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
X_13853_ fifo_bank_register.bank\[5\]\[33\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[33\]
+ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12804_ fifo_bank_register.bank\[2\]\[65\] _05407_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07702_ sky130_fd_sc_hd__mux2_1
X_16572_ net504 _00020_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10996_ mix1.data_o\[123\] _05676_ _05758_ _05620_ sub1.data_o\[123\] vssd1 vssd1
+ vccd1 vccd1 _06732_ sky130_fd_sc_hd__a32o_1
X_13784_ _02194_ fifo_bank_register.data_out\[25\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18311_ clknet_leaf_5_clk _01742_ net624 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[77\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15523_ _03668_ _04777_ _05236_ _03680_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__a31o_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12735_ fifo_bank_register.bank\[2\]\[32\] _05338_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07666_ sky130_fd_sc_hd__mux2_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ clknet_leaf_10_clk _01673_ net623 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15454_ sub1.data_o\[64\] _05547_ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__mux2_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12666_ _07628_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14405_ _02747_ fifo_bank_register.data_out\[93\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02748_ sky130_fd_sc_hd__mux2_1
X_11617_ fifo_bank_register.bank\[6\]\[17\] _05305_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07075_ sky130_fd_sc_hd__mux2_1
X_18173_ clknet_leaf_20_clk _01604_ net640 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15385_ _03590_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__clkbuf_1
X_12597_ _07592_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17124_ net430 _00567_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11548_ _07038_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__clkbuf_1
X_14336_ fifo_bank_register.bank\[9\]\[86\] _02631_ _02683_ _02684_ _02685_ vssd1
+ vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_29_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14267_ fifo_bank_register.bank\[5\]\[79\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[79\]
+ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__a22o_1
X_17055_ net536 _00498_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ _06935_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__buf_4
XFILLER_0_208_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13218_ _07920_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__clkbuf_1
X_16006_ _05007_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__or2_1
XFILLER_0_204_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14198_ fifo_bank_register.bank\[0\]\[70\] _02562_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02564_ sky130_fd_sc_hd__mux2_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ fifo_bank_register.bank\[1\]\[100\] _05480_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07884_ sky130_fd_sc_hd__mux2_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ net402 _01400_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16908_ net519 _00351_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08690_ addroundkey_data_o\[68\] mix1.data_o\[68\] _04663_ vssd1 vssd1 vccd1 vccd1
+ _04714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17888_ net510 _01331_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16839_ net439 _00282_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09311_ _05300_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18509_ clknet_leaf_62_clk _01938_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09242_ ks1.state\[1\] _04723_ _04749_ _04737_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__o31a_1
XFILLER_0_180_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09173_ _05145_ _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_56_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput106 data_i[7] vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_4
XTAP_5328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput117 data_i[8] vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__buf_2
Xinput128 data_i[9] vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_4
XTAP_5339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput139 key_i[108] vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ _04677_ _04979_ _04980_ _04682_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_216_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ ks1.key_reg\[8\] _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__or3_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ mix1.data_o\[108\] _06463_ _06575_ _06576_ sub1.data_o\[108\] vssd1 vssd1
+ vccd1 vccd1 _06601_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ fifo_bank_register.bank\[9\]\[78\] _05434_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05435_ sky130_fd_sc_hd__mux2_1
X_10781_ sub1.data_o\[101\] _06513_ _06537_ _06538_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06539_ sky130_fd_sc_hd__a221o_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12520_ fifo_bank_register.bank\[3\]\[59\] _05394_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07552_ sky130_fd_sc_hd__mux2_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12451_ fifo_bank_register.bank\[3\]\[26\] _05325_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11402_ fifo_bank_register.bank\[7\]\[43\] _05361_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15170_ net727 _03435_ _03425_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12382_ _05528_ fifo_bank_register.bank\[4\]\[123\] _07341_ vssd1 vssd1 vccd1 vccd1
+ _07478_ sky130_fd_sc_hd__mux2_1
XANTENNA_90 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14121_ fifo_bank_register.bank\[1\]\[62\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[62\]
+ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__a22o_1
X_11333_ _06925_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ fifo_bank_register.bank\[7\]\[55\] _02380_ _02389_ fifo_bank_register.bank\[2\]\[55\]
+ _02432_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__a221o_1
X_11264_ _05495_ fifo_bank_register.bank\[8\]\[107\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06888_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13003_ _07807_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__clkbuf_1
X_10215_ _06027_ _06028_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__xor2_1
X_11195_ _05426_ fifo_bank_register.bank\[8\]\[74\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17811_ net553 _01254_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
X_10146_ _05965_ _05966_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_182_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17742_ net477 _01185_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10077_ _05201_ _05754_ sub1.data_o\[33\] _05902_ vssd1 vssd1 vccd1 vccd1 _05903_
+ sky130_fd_sc_hd__a31o_1
X_14954_ addroundkey_data_o\[81\] _03209_ _03067_ addroundkey_data_o\[49\] vssd1 vssd1
+ vccd1 vccd1 _03229_ sky130_fd_sc_hd__a22o_1
XTAP_5884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13905_ fifo_bank_register.bank\[6\]\[39\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[39\]
+ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17673_ net515 _01116_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14885_ sub1.data_o\[95\] _03061_ _03065_ sub1.data_o\[63\] vssd1 vssd1 vccd1 vccd1
+ _03161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16624_ net514 _00072_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13836_ _02241_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16555_ clknet_leaf_28_clk _00003_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[118\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10979_ sub1.data_o\[121\] _06716_ _06573_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__mux2_1
X_13767_ fifo_bank_register.bank\[0\]\[23\] _02179_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15506_ _05103_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_174_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12718_ fifo_bank_register.bank\[2\]\[24\] _05321_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16486_ _04326_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__clkbuf_1
X_13698_ fifo_bank_register.bank\[9\]\[17\] _08190_ _02114_ _02115_ _02116_ vssd1
+ vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18225_ clknet_leaf_36_clk _01656_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[55\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_170_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15437_ sub1.data_o\[24\] _05547_ _04879_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ _07619_ vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18156_ clknet_leaf_67_clk _01587_ net610 vssd1 vssd1 vccd1 vccd1 ks1.col\[26\] sky130_fd_sc_hd__dfrtp_2
X_15368_ sub1.data_o\[1\] _03578_ _03576_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17107_ net505 _00550_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14319_ fifo_bank_register.bank\[1\]\[84\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[84\]
+ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__a22o_1
X_18087_ net472 _01530_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15299_ _03541_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17038_ net546 _00481_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ net141 ks1.key_reg\[10\] _05708_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ addroundkey_data_o\[22\] mix1.data_o\[22\] _04662_ vssd1 vssd1 vccd1 vccd1
+ _04835_ sky130_fd_sc_hd__mux2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ mix1.data_o\[3\] _05586_ _05618_ _05621_ sub1.data_o\[3\] vssd1 vssd1 vccd1
+ vccd1 _05647_ sky130_fd_sc_hd__a32o_1
XFILLER_0_175_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _04713_ _04764_ _04668_ _04765_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__a22o_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08673_ addroundkey_data_o\[44\] _04693_ _04695_ addroundkey_data_o\[36\] vssd1 vssd1
+ vccd1 vccd1 _04697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09225_ _05145_ _05224_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__xor2_4
XFILLER_0_146_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09156_ _05109_ _05110_ sbox1.ah_reg\[1\] vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ sbox1.ah\[1\] _05067_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ net174 ks1.key_reg\[24\] _05825_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09989_ _05707_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__buf_4
XTAP_5147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _07251_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10902_ addroundkey_data_o\[113\] _06647_ _06612_ vssd1 vssd1 vccd1 vccd1 _06648_
+ sky130_fd_sc_hd__mux2_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14670_ fifo_bank_register.bank\[5\]\[124\] _08096_ _08099_ fifo_bank_register.bank\[3\]\[124\]
+ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__a22o_1
X_11882_ fifo_bank_register.bank\[5\]\[14\] _05299_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10833_ mix1.data_o\[106\] _06463_ _06575_ _06576_ sub1.data_o\[106\] vssd1 vssd1
+ vccd1 vccd1 _06586_ sky130_fd_sc_hd__a32o_1
X_13621_ fifo_bank_register.bank\[5\]\[9\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[9\]
+ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_196_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16340_ _04245_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13552_ _08122_ fifo_bank_register.data_out\[0\] _08064_ vssd1 vssd1 vccd1 vccd1
+ _08123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10764_ _06523_ vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ _07543_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__clkbuf_1
X_13483_ _08057_ _08058_ _08059_ _08060_ _08061_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__a221o_1
X_16271_ _04208_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10695_ _06460_ vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18010_ net500 _01453_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_15222_ _03188_ _03417_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__xor2_1
X_12434_ _07506_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ _03417_ _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12365_ _07469_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11316_ _06916_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__clkbuf_1
X_14104_ fifo_bank_register.bank\[1\]\[60\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[60\]
+ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__a22o_1
X_15084_ sub1.data_o\[12\] _04378_ _03059_ _03355_ vssd1 vssd1 vccd1 vccd1 _03356_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ _07433_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14035_ fifo_bank_register.bank\[5\]\[53\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[53\]
+ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11247_ _05478_ fifo_bank_register.bank\[8\]\[99\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11178_ _05409_ fifo_bank_register.bank\[8\]\[66\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ _05949_ _05948_ _05950_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ _04961_ _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17725_ net430 _01168_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14937_ sub1.data_o\[96\] _03056_ _03211_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ net556 _01099_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_14868_ _03072_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__buf_6
XFILLER_0_37_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16607_ net396 _00055_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_13819_ _02225_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17587_ net458 _01030_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
X_14799_ addroundkey_data_o\[112\] _03057_ _03074_ vssd1 vssd1 vccd1 vccd1 _03075_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16538_ _04353_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16469_ _04317_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09010_ addroundkey_data_o\[42\] _04692_ _04694_ addroundkey_data_o\[34\] vssd1 vssd1
+ vccd1 vccd1 _05032_ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18208_ clknet_leaf_15_clk _01639_ net629 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18139_ clknet_leaf_53_clk sbox1.next_alph\[1\] net656 vssd1 vssd1 vccd1 vccd1 sbox1.alph\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold102 mix1.data_reg\[33\] vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold113 mix1.data_reg\[84\] vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold124 ks1.key_reg\[114\] vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold135 ks1.key_reg\[86\] vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 ks1.key_reg\[51\] vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 ks1.key_reg\[97\] vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 ks1.key_reg\[65\] vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _05201_ _05754_ sub1.data_o\[16\] _05585_ vssd1 vssd1 vccd1 vccd1 _05755_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold179 ks1.key_reg\[127\] vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout604 net607 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_4
Xfanout615 net617 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout626 net635 vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__buf_2
Xfanout637 net638 vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__buf_2
X_09843_ _05629_ _05691_ _05692_ _05633_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__a22o_1
Xfanout648 net649 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_4
Xfanout659 net660 vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ mix1.data_o\[1\] _05586_ _05618_ _05621_ sub1.data_o\[1\] vssd1 vssd1 vccd1
+ vccd1 _05632_ sky130_fd_sc_hd__a32o_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _04644_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__inv_2
XFILLER_0_197_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08656_ sub1.state\[1\] _04673_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__or2_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08587_ round\[3\] _04614_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09208_ _05214_ _05217_ _04649_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__mux2_8
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ sub1.data_o\[72\] _06266_ _06239_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09139_ sbox1.alph\[2\] _05111_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12150_ _07356_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11101_ _06802_ vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12081_ _07319_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11032_ addroundkey_data_o\[127\] _06763_ _05696_ vssd1 vssd1 vccd1 vccd1 _06764_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15840_ _03852_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__clkbuf_1
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _03816_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__clkbuf_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ fifo_bank_register.bank\[1\]\[21\] _05315_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07797_ sky130_fd_sc_hd__mux2_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ net419 _00953_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_14722_ sub1.data_o\[54\] sub1.data_o\[118\] _05598_ vssd1 vssd1 vccd1 vccd1 _03024_
+ sky130_fd_sc_hd__mux2_1
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _07242_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__clkbuf_1
X_18490_ clknet_leaf_54_clk _01919_ net615 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17441_ net401 _00884_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
X_14653_ _02967_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__clkbuf_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ fifo_bank_register.bank\[5\]\[6\] _05282_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07206_ sky130_fd_sc_hd__mux2_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ fifo_bank_register.bank\[6\]\[7\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17372_ net500 _00815_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10816_ _06570_ vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__clkbuf_1
X_14584_ fifo_bank_register.bank\[1\]\[113\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[113\]
+ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__a22o_1
X_11796_ _07169_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16323_ _04189_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13535_ _08069_ _08094_ vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10747_ net255 ks1.key_reg\[98\] _06402_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16254_ net217 ks1.key_reg\[63\] _03982_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__mux2_1
X_13466_ _08050_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__clkbuf_1
X_10678_ addroundkey_data_o\[91\] _06445_ _06431_ vssd1 vssd1 vccd1 vccd1 _06446_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15205_ net780 _03467_ _03425_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12417_ fifo_bank_register.bank\[3\]\[10\] _05290_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07498_ sky130_fd_sc_hd__mux2_1
X_16185_ _04761_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_211_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13397_ _08014_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ _03099_ _03131_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12348_ _07460_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15067_ sub1.data_o\[116\] _03057_ _03338_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__a21oi_2
X_12279_ _07424_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _02403_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15969_ ks1.key_reg\[3\] _03940_ _04373_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__mux2_1
X_08510_ addroundkey_data_o\[94\] fifo_bank_register.data_out\[94\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__mux2_4
XFILLER_0_222_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17708_ net464 _01151_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09490_ net227 vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08441_ addroundkey_data_o\[61\] fifo_bank_register.data_out\[61\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ net424 _01082_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08372_ _04500_ vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_176_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout401 net404 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__buf_2
Xfanout412 net413 vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_2
Xfanout423 net427 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__buf_2
XFILLER_0_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout434 net436 vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_2
XFILLER_0_10_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout445 net449 vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__buf_2
Xfanout456 net460 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__buf_2
XFILLER_0_201_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09826_ mix1.data_o\[7\] _05677_ _05618_ _05621_ sub1.data_o\[7\] vssd1 vssd1 vccd1
+ vccd1 _05678_ sky130_fd_sc_hd__a32o_1
Xfanout467 net468 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
Xfanout478 net481 vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__clkbuf_2
Xfanout489 net530 vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_214_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09757_ _04618_ _04629_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__nor2_2
XFILLER_0_213_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _04731_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__buf_2
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09688_ _05213_ _05557_ _04649_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _04662_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__buf_4
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11650_ fifo_bank_register.bank\[6\]\[32\] _05338_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07093_ sky130_fd_sc_hd__mux2_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10601_ sub1.data_o\[84\] _06341_ _06374_ _06375_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06376_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11581_ _07055_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13320_ _07974_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10532_ net233 ks1.key_reg\[78\] _06245_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10463_ sub1.data_o\[70\] _06251_ _06239_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__mux2_1
X_13251_ _07937_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__buf_4
XFILLER_0_134_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12202_ _05348_ fifo_bank_register.bank\[4\]\[37\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13182_ fifo_bank_register.bank\[1\]\[116\] _05514_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10394_ net216 ks1.key_reg\[62\] _06166_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_206_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12133_ _07347_ vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17990_ net442 _01433_ net596 vssd1 vssd1 vccd1 vccd1 fifo_bank_register.read_ptr\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_202_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12064_ fifo_bank_register.bank\[5\]\[100\] _05480_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07311_ sky130_fd_sc_hd__mux2_1
X_16941_ net467 _00384_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11015_ _06747_ _06748_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16872_ net430 _00315_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18611_ clknet_leaf_12_clk _02040_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[104\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ mix1.data_o\[111\] net745 _03841_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ clknet_leaf_79_clk _01971_ net579 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[69\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _03807_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__clkbuf_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12966_ _07787_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__clkbuf_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _05104_ _04927_ _05548_ _03012_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a31o_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ fifo_bank_register.bank\[5\]\[30\] _05333_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07234_ sky130_fd_sc_hd__mux2_1
X_18473_ clknet_leaf_57_clk _01902_ net602 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15685_ _03771_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__clkbuf_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_350 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ _07750_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__clkbuf_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17424_ net546 _00867_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14636_ _02952_ fifo_bank_register.data_out\[119\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _02953_ sky130_fd_sc_hd__mux2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11848_ fifo_bank_register.bank\[6\]\[127\] _05536_ _07055_ vssd1 vssd1 vccd1 vccd1
+ _07196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ net474 _00798_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14567_ fifo_bank_register.bank\[6\]\[111\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[111\]
+ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__a22o_1
X_11779_ _07160_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16306_ _04227_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__clkbuf_1
X_13518_ _08088_ vssd1 vssd1 vccd1 vccd1 _08089_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17286_ net512 _00729_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14498_ fifo_bank_register.bank\[5\]\[104\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[104\]
+ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16237_ _04111_ _04112_ _04126_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__or3_2
XFILLER_0_10_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13449_ _05510_ fifo_bank_register.bank\[0\]\[114\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16168_ _04117_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15119_ _03385_ _03387_ _03388_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__o21a_2
XFILLER_0_140_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08990_ _04649_ _05009_ _05011_ _05012_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__o2bb2a_4
X_16099_ _04754_ _04056_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09611_ net143 vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09542_ net245 vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__buf_2
XFILLER_0_222_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09473_ _05410_ vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08424_ addroundkey_data_o\[53\] fifo_bank_register.data_out\[53\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08355_ addroundkey_data_o\[20\] fifo_bank_register.data_out\[20\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__mux2_4
XFILLER_0_188_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08286_ net167 net170 net171 net168 vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09809_ net213 ks1.key_reg\[5\] _05625_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__mux2_2
XFILLER_0_96_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12820_ _07710_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12751_ _07651_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__buf_4
XFILLER_0_201_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_81_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_210_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ fifo_bank_register.bank\[6\]\[57\] _05390_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07120_ sky130_fd_sc_hd__mux2_1
X_15470_ _03645_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _07637_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__clkbuf_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _02761_ fifo_bank_register.data_out\[95\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11633_ fifo_bank_register.bank\[6\]\[24\] _05321_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07084_ sky130_fd_sc_hd__mux2_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17140_ net390 _00583_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14352_ fifo_bank_register.bank\[1\]\[88\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[88\]
+ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11564_ _07046_ vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13303_ _07965_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__clkbuf_1
X_10515_ _06250_ _06295_ _06297_ _06254_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__a22o_2
X_17071_ net467 _00514_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
X_14283_ fifo_bank_register.bank\[6\]\[80\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[80\]
+ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11495_ _07010_ vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16022_ net136 ks1.key_reg\[105\] _03976_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__mux2_1
X_10446_ _06236_ vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__clkbuf_1
X_13234_ _05295_ fifo_bank_register.bank\[0\]\[12\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10377_ _06171_ _06173_ _06174_ _06175_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__a22o_1
X_13165_ fifo_bank_register.bank\[1\]\[108\] _05497_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ _07337_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__clkbuf_1
X_17973_ net411 _01416_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
X_13096_ fifo_bank_register.bank\[1\]\[75\] _05428_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12047_ fifo_bank_register.bank\[5\]\[92\] _05464_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07302_ sky130_fd_sc_hd__mux2_1
X_16924_ net547 _00367_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16855_ net532 _00298_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15806_ mix1.data_o\[103\] net728 _03830_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16786_ clknet_leaf_73_clk _00230_ net590 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[77\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_204_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13998_ fifo_bank_register.bank\[9\]\[49\] _02307_ _02382_ _02383_ _02384_ vssd1
+ vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_220_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18525_ clknet_leaf_67_clk _01954_ net606 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
X_15737_ mix1.data_o\[70\] net697 _03797_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__mux2_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ _07778_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18456_ clknet_leaf_27_clk _01886_ net642 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[96\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_158_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15668_ _03762_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_180 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_173_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_191 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17407_ net550 _00850_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14619_ _08063_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__clkbuf_8
X_18387_ clknet_leaf_12_clk _01817_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[72\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15599_ _03725_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17338_ net412 _00781_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17269_ net396 _00712_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08973_ _04988_ _04990_ _04993_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__or4_2
XFILLER_0_228_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold17 mix1.data_reg\[105\] vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 ks1.key_reg\[21\] vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_227_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold39 mix1.data_reg\[100\] vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09525_ fifo_bank_register.bank\[9\]\[83\] _05445_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_63_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk
+ sky130_fd_sc_hd__clkbuf_16
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ net215 vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__clkbuf_4
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08407_ addroundkey_data_o\[45\] fifo_bank_register.data_out\[45\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__mux2_2
XFILLER_0_136_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09387_ net190 vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08338_ addroundkey_data_o\[12\] fifo_bank_register.data_out\[12\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__mux2_4
XFILLER_0_163_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ net134 net133 net136 net135 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__and4b_1
XFILLER_0_229_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ sub1.data_o\[53\] _05971_ _06104_ _06105_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _06106_ sky130_fd_sc_hd__a221o_1
XFILLER_0_166_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11280_ _06896_ vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10231_ _06041_ _06042_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10162_ _05981_ vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10093_ sub1.data_o\[34\] _05753_ _05915_ _05917_ _04611_ vssd1 vssd1 vccd1 vccd1
+ _05918_ sky130_fd_sc_hd__a221o_1
X_14970_ addroundkey_data_o\[111\] _03078_ _03243_ vssd1 vssd1 vccd1 vccd1 _03244_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13921_ _02153_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ net565 _00088_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ _02255_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12803_ _07701_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__clkbuf_1
X_16571_ net533 _00019_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_13783_ fifo_bank_register.bank\[0\]\[25\] _02193_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10995_ sub1.data_o\[123\] _06730_ _05609_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18310_ clknet_leaf_2_clk _01741_ net624 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[76\]
+ sky130_fd_sc_hd__dfrtp_2
X_15522_ sub1.data_o\[54\] _03663_ _03679_ _03673_ vssd1 vssd1 vccd1 vccd1 _03680_
+ sky130_fd_sc_hd__a22o_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12734_ _07665_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18241_ clknet_leaf_35_clk _01672_ net662 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _05198_ _04368_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__nand2_4
XFILLER_0_132_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12665_ _07627_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__buf_4
XFILLER_0_167_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14404_ fifo_bank_register.bank\[0\]\[93\] _02746_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02747_ sky130_fd_sc_hd__mux2_1
X_18172_ clknet_leaf_20_clk _01603_ net640 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11616_ _07074_ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15384_ sub1.data_o\[6\] _03589_ _03581_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12596_ fifo_bank_register.bank\[3\]\[95\] _05470_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17123_ net499 _00566_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14335_ fifo_bank_register.bank\[1\]\[86\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[86\]
+ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11547_ fifo_bank_register.bank\[7\]\[112\] _05506_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17054_ net541 _00497_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14266_ _08181_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11478_ _07001_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16005_ _03971_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__xor2_2
XFILLER_0_208_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13217_ _05278_ fifo_bank_register.bank\[0\]\[4\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07920_ sky130_fd_sc_hd__mux2_1
X_10429_ addroundkey_data_o\[66\] _06221_ _06169_ vssd1 vssd1 vccd1 vccd1 _06222_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14197_ _02157_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _07794_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__buf_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ fifo_bank_register.bank\[1\]\[67\] _05411_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07847_ sky130_fd_sc_hd__mux2_1
X_17956_ net455 _01399_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16907_ net518 _00350_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
X_17887_ net508 _01330_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16838_ net421 _00281_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16769_ clknet_leaf_48_clk _00213_ net611 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[60\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_177_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_221_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09310_ fifo_bank_register.bank\[9\]\[14\] _05299_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18508_ clknet_leaf_67_clk _01937_ net606 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09241_ _05104_ _04946_ _05245_ _05247_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__a31o_1
X_18439_ clknet_leaf_36_clk _01869_ net666 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[124\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09172_ _05175_ _05182_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput107 data_i[80] vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput118 data_i[90] vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_228_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08956_ addroundkey_data_o\[119\] mix1.data_o\[119\] _04778_ vssd1 vssd1 vccd1 vccd1
+ _04980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput129 decrypt_i vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_4
XTAP_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08887_ _04738_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__buf_4
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09508_ net233 vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__clkbuf_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ mix1.data_o\[101\] _06494_ _06398_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _05387_ vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__clkbuf_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ _07515_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ _06961_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12381_ _07477_ vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_80 addroundkey_data_o\[69\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_91 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ fifo_bank_register.bank\[6\]\[62\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[62\]
+ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__a22o_1
X_11332_ fifo_bank_register.bank\[7\]\[10\] _05290_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14051_ fifo_bank_register.bank\[5\]\[55\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[55\]
+ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a22o_1
X_11263_ _06887_ vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13002_ fifo_bank_register.bank\[1\]\[30\] _05333_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10214_ net197 ks1.key_reg\[45\] _05997_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__mux2_1
X_11194_ _06851_ vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17810_ net545 _01253_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
X_10145_ net189 ks1.key_reg\[38\] _05920_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__mux2_4
XTAP_5830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17741_ net477 _01184_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10076_ _05584_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__buf_2
X_14953_ sub1.data_o\[113\] _03056_ _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a21oi_1
XTAP_5874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ fifo_bank_register.bank\[7\]\[39\] _02299_ _02227_ fifo_bank_register.bank\[2\]\[39\]
+ _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17672_ net521 _01115_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14884_ _03156_ _03159_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__nor2_8
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16623_ net524 _00071_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _02240_ fifo_bank_register.data_out\[30\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_203_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16554_ clknet_leaf_28_clk _00002_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[117\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ fifo_bank_register.bank\[9\]\[23\] _02137_ _02176_ _02177_ _02178_ vssd1
+ vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ net25 mix1.data_o\[121\] _06571_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15505_ _03652_ _04777_ _05554_ _03667_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a31o_1
XFILLER_0_186_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12717_ _07656_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__clkbuf_1
X_16485_ net709 _03363_ _04321_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13697_ fifo_bank_register.bank\[1\]\[17\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18224_ clknet_leaf_36_clk _01655_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[54\]
+ sky130_fd_sc_hd__dfrtp_1
X_15436_ _03603_ _04949_ _05245_ _03624_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a31o_1
X_12648_ fifo_bank_register.bank\[3\]\[120\] _05522_ _07485_ vssd1 vssd1 vccd1 vccd1
+ _07619_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18155_ clknet_leaf_48_clk _01586_ net610 vssd1 vssd1 vccd1 vccd1 ks1.col\[25\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15367_ sub1.data_o\[33\] sub1.data_o\[97\] _03574_ vssd1 vssd1 vccd1 vccd1 _03578_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12579_ fifo_bank_register.bank\[3\]\[87\] _05453_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17106_ net504 _00549_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14318_ fifo_bank_register.bank\[6\]\[84\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[84\]
+ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
X_18086_ net541 _01529_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[88\]
+ sky130_fd_sc_hd__dfxtp_2
X_15298_ net772 _03236_ _03539_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17037_ net519 _00480_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14249_ fifo_bank_register.bank\[5\]\[77\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[77\]
+ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08810_ addroundkey_data_o\[126\] mix1.data_o\[126\] _04657_ vssd1 vssd1 vccd1 vccd1
+ _04834_ sky130_fd_sc_hd__mux2_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ sub1.data_o\[3\] _05645_ _05610_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__mux2_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ addroundkey_data_o\[73\] mix1.data_o\[73\] _04655_ vssd1 vssd1 vccd1 vccd1
+ _04765_ sky130_fd_sc_hd__mux2_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ net555 _01382_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08672_ mix1.data_o\[44\] _04693_ _04695_ mix1.data_o\[36\] vssd1 vssd1 vccd1 vccd1
+ _04696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09224_ _05145_ _05171_ _05060_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09155_ _05124_ _05125_ _05126_ sbox1.ah_reg\[2\] vssd1 vssd1 vccd1 vccd1 _05166_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09086_ _05092_ _05098_ vssd1 vssd1 vccd1 vccd1 sbox1.intermediate_to_invert_var\[1\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09988_ _05712_ _05820_ _05823_ _05716_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_216_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08939_ ks1.key_reg\[29\] _04725_ _04962_ net179 vssd1 vssd1 vccd1 vccd1 _04963_
+ sky130_fd_sc_hd__a22o_1
XTAP_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ fifo_bank_register.bank\[5\]\[46\] _05367_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10901_ _06645_ _06646_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__xnor2_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ _07214_ vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13620_ _08181_ vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__buf_4
XFILLER_0_200_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10832_ sub1.data_o\[106\] _06584_ _06573_ vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13551_ fifo_bank_register.bank\[0\]\[0\] _08117_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10763_ addroundkey_data_o\[99\] _06521_ _06522_ vssd1 vssd1 vccd1 vccd1 _06523_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_165_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ fifo_bank_register.bank\[3\]\[50\] _05375_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16270_ ks1.key_reg\[37\] _03955_ _04206_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__mux2_1
X_13482_ fifo_bank_register.read_ptr\[1\] _05250_ vssd1 vssd1 vccd1 vccd1 _08061_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10694_ addroundkey_data_o\[93\] _06459_ _06431_ vssd1 vssd1 vccd1 vccd1 _06460_
+ sky130_fd_sc_hd__mux2_1
X_15221_ _03480_ _03481_ _05198_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__a21o_2
XFILLER_0_129_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12433_ fifo_bank_register.bank\[3\]\[18\] _05307_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15152_ _03245_ _03418_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__xnor2_2
X_12364_ _05510_ fifo_bank_register.bank\[4\]\[114\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14103_ _02153_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__buf_4
XFILLER_0_121_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11315_ fifo_bank_register.bank\[7\]\[2\] _05274_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06916_ sky130_fd_sc_hd__mux2_1
X_15083_ sub1.data_o\[76\] _03072_ _03068_ sub1.data_o\[44\] vssd1 vssd1 vccd1 vccd1
+ _03355_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12295_ _05441_ fifo_bank_register.bank\[4\]\[81\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14034_ _02417_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11246_ _06878_ vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ _06842_ vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10128_ _05913_ _05754_ sub1.data_o\[37\] _05902_ vssd1 vssd1 vccd1 vccd1 _05950_
+ sky130_fd_sc_hd__a31o_1
X_15985_ _03953_ _03954_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__xor2_2
XTAP_5660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14936_ sub1.data_o\[0\] _03208_ _03081_ _03210_ vssd1 vssd1 vccd1 vccd1 _03211_
+ sky130_fd_sc_hd__a211o_1
X_10059_ _05885_ _05886_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__xor2_1
X_17724_ net407 _01167_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14867_ _03057_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__buf_8
X_17655_ net407 _01098_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16606_ net394 _00054_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_13818_ _02224_ fifo_bank_register.data_out\[29\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17586_ net451 _01029_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
X_14798_ addroundkey_data_o\[16\] _04378_ _05607_ _03073_ vssd1 vssd1 vccd1 vccd1
+ _03074_ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16537_ net729 _03529_ _04343_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__mux2_1
X_13749_ fifo_bank_register.bank\[1\]\[21\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16468_ ks1.key_reg\[126\] _04316_ _03957_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15419_ sub1.data_o\[114\] sub1.data_o\[50\] _03609_ vssd1 vssd1 vccd1 vccd1 _03613_
+ sky130_fd_sc_hd__mux2_1
X_18207_ clknet_leaf_15_clk _01638_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16399_ ks1.key_reg\[95\] _04278_ _04264_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18138_ clknet_leaf_42_clk sbox1.next_alph\[0\] net656 vssd1 vssd1 vccd1 vccd1 sbox1.alph\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_131_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold103 mix1.data_reg\[93\] vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold114 mix1.data_reg\[101\] vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18069_ net527 _01512_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[71\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold125 ks1.key_reg\[27\] vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold136 ks1.col\[0\] vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold147 ks1.key_reg\[78\] vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 ks1.key_reg\[98\] vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09911_ sub1.ready_o vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__buf_2
XFILLER_0_229_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold169 mix1.data_reg\[68\] vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout605 net607 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_4
Xfanout616 net617 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__buf_2
X_09842_ mix1.data_o\[9\] _05677_ _05618_ _05621_ sub1.data_o\[9\] vssd1 vssd1 vccd1
+ vccd1 _05692_ sky130_fd_sc_hd__a32o_1
Xfanout627 net634 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout638 net639 vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__buf_2
XFILLER_0_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout649 net650 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_4
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09773_ sub1.data_o\[1\] _05630_ _05610_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__mux2_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08724_ ks1.key_reg\[28\] _04735_ _04747_ net178 vssd1 vssd1 vccd1 vccd1 _04748_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08655_ addroundkey_data_o\[116\] mix1.data_o\[116\] _04666_ vssd1 vssd1 vccd1 vccd1
+ _04679_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08586_ round\[1\] _04613_ round\[2\] vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__or3_2
XFILLER_0_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09207_ _05215_ _05216_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_107_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09138_ sbox1.alph\[1\] _05119_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_162_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09069_ _05057_ _05071_ _04971_ _05016_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__and4b_1
XFILLER_0_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11100_ _05331_ fifo_bank_register.bank\[8\]\[29\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12080_ fifo_bank_register.bank\[5\]\[108\] _05497_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11031_ _06761_ _06762_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__xor2_1
XFILLER_0_216_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15770_ mix1.data_o\[86\] net792 _03808_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _07796_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__clkbuf_1
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _03019_ _04927_ _05228_ _03023_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a31o_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ fifo_bank_register.bank\[5\]\[38\] _05350_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ net409 _00883_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _02966_ fifo_bank_register.data_out\[121\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _02967_ sky130_fd_sc_hd__mux2_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11864_ _07205_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__clkbuf_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13603_ fifo_bank_register.bank\[7\]\[7\] _08078_ _08093_ fifo_bank_register.bank\[2\]\[7\]
+ _08166_ vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__a221o_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17371_ net482 _00814_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ addroundkey_data_o\[104\] _06569_ _06522_ vssd1 vssd1 vccd1 vccd1 _06570_
+ sky130_fd_sc_hd__mux2_1
X_14583_ fifo_bank_register.bank\[6\]\[113\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[113\]
+ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11795_ fifo_bank_register.bank\[6\]\[101\] _05483_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16322_ _04215_ _04179_ _04235_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__o21ai_1
X_13534_ _08104_ vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__clkbuf_4
X_10746_ _06381_ _06502_ _06506_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16253_ _04195_ _04196_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__xor2_4
X_13465_ _05526_ fifo_bank_register.bank\[0\]\[122\] _07914_ vssd1 vssd1 vccd1 vccd1
+ _08050_ sky130_fd_sc_hd__mux2_1
X_10677_ _06443_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15204_ _03464_ _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__xor2_4
X_12416_ _07485_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__buf_4
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16184_ _04132_ _04133_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__xor2_2
XFILLER_0_140_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13396_ _05457_ fifo_bank_register.bank\[0\]\[89\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08014_ sky130_fd_sc_hd__mux2_1
X_15135_ _03403_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12347_ _05493_ fifo_bank_register.bank\[4\]\[106\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15066_ sub1.data_o\[20\] _04378_ _03059_ _03337_ vssd1 vssd1 vccd1 vccd1 _03338_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12278_ _05424_ fifo_bank_register.bank\[4\]\[73\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07424_ sky130_fd_sc_hd__mux2_1
X_14017_ _02402_ fifo_bank_register.data_out\[50\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02403_ sky130_fd_sc_hd__mux2_1
X_11229_ _05459_ fifo_bank_register.bank\[8\]\[90\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15968_ _04800_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__xnor2_1
X_17707_ net450 _01150_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
X_14919_ addroundkey_data_o\[110\] _03055_ _03193_ vssd1 vssd1 vccd1 vccd1 _03194_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15899_ _03885_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08440_ _04536_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17638_ net419 _01081_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08371_ addroundkey_data_o\[28\] fifo_bank_register.data_out\[28\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17569_ net401 _01012_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout402 net404 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__buf_2
Xfanout413 net444 vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_2
Xfanout424 net427 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_2
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_2
Xfanout446 net449 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_2
X_09825_ _05676_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__clkbuf_4
Xfanout457 net460 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__clkbuf_2
Xfanout468 net472 vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout479 net481 vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_2
XFILLER_0_214_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09756_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08707_ _04641_ _04722_ addroundkey_start_i vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__o21a_4
XFILLER_0_119_1256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09687_ _05191_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__xnor2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08638_ _04654_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08569_ _04603_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10600_ mix1.data_o\[84\] _06129_ _06093_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11580_ _07054_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__buf_4
XFILLER_0_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10531_ _06250_ _06310_ _06311_ _06254_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__a22o_2
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _07913_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__clkbuf_8
X_10462_ net96 mix1.data_o\[70\] _06237_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12201_ _07383_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13181_ _07900_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__clkbuf_1
X_10393_ _06171_ _06188_ _06189_ _06175_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12132_ _05278_ fifo_bank_register.bank\[4\]\[4\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12063_ _07221_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__buf_4
X_16940_ net465 _00383_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
X_11014_ net158 ks1.key_reg\[125\] _05762_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16871_ net423 _00314_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18610_ clknet_leaf_13_clk _02039_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[103\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _03843_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__clkbuf_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ mix1.data_o\[78\] net737 _03797_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__mux2_1
X_18541_ clknet_leaf_62_clk _01970_ net601 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[68\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ fifo_bank_register.bank\[1\]\[13\] _05297_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07787_ sky130_fd_sc_hd__mux2_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ sub1.data_o\[80\] _03010_ _03011_ sub1.next_ready_o vssd1 vssd1 vccd1 vccd1
+ _03012_ sky130_fd_sc_hd__a22o_1
X_11916_ _07221_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__buf_4
X_18472_ clknet_leaf_33_clk mix1.next_ready_o net660 vssd1 vssd1 vccd1 vccd1 mix1.ready_o
+ sky130_fd_sc_hd__dfrtp_2
X_15684_ mix1.data_o\[45\] net718 _03764_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__mux2_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_340 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12896_ fifo_bank_register.bank\[2\]\[109\] _05499_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_351 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14635_ fifo_bank_register.bank\[0\]\[119\] _02951_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02952_ sky130_fd_sc_hd__mux2_1
X_17423_ net552 _00866_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11847_ _07195_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__clkbuf_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17354_ net474 _00797_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_14566_ fifo_bank_register.bank\[7\]\[111\] _02866_ _02875_ fifo_bank_register.bank\[2\]\[111\]
+ _02890_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a221o_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11778_ fifo_bank_register.bank\[6\]\[93\] _05466_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07160_ sky130_fd_sc_hd__mux2_1
X_13517_ _08056_ _08087_ vssd1 vssd1 vccd1 vccd1 _08088_ sky130_fd_sc_hd__and2_1
X_16305_ net810 _04088_ _04222_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__mux2_1
X_10729_ _05574_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17285_ net522 _00728_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14497_ _02829_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16236_ _04181_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13448_ _08041_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ net244 ks1.key_reg\[88\] _03906_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__mux2_1
X_13379_ _08005_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15118_ _03385_ _03387_ _05198_ vssd1 vssd1 vccd1 vccd1 _03388_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_224_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16098_ _04054_ _04055_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__xor2_2
XFILLER_0_103_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15049_ _03314_ _03321_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_220_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09610_ _05503_ vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09541_ _05456_ vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09472_ fifo_bank_register.bank\[9\]\[66\] _05409_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08423_ _04527_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ _04491_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08285_ net164 net166 net165 net163 vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_172_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09808_ _05629_ _05660_ _05661_ _05633_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_213_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09739_ _05598_ addroundkey_ready_o _04618_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12750_ _07673_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11701_ _07119_ vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__clkbuf_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ fifo_bank_register.bank\[2\]\[7\] _05284_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ fifo_bank_register.bank\[0\]\[95\] _02760_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02761_ sky130_fd_sc_hd__mux2_1
X_11632_ _07083_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__clkbuf_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14351_ fifo_bank_register.bank\[6\]\[88\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[88\]
+ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11563_ fifo_bank_register.bank\[7\]\[120\] _05522_ _06912_ vssd1 vssd1 vccd1 vccd1
+ _07046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13302_ _05363_ fifo_bank_register.bank\[0\]\[44\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07965_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10514_ mix1.data_o\[76\] _06296_ _06241_ _06242_ sub1.data_o\[76\] vssd1 vssd1 vccd1
+ vccd1 _06297_ sky130_fd_sc_hd__a32o_1
X_17070_ net462 _00513_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14282_ _02148_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__clkbuf_4
X_11494_ fifo_bank_register.bank\[7\]\[87\] _05453_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16021_ net228 ks1.key_reg\[73\] _03979_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ _07928_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ addroundkey_data_o\[68\] _06235_ _06169_ vssd1 vssd1 vccd1 vccd1 _06236_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13164_ _07891_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__clkbuf_1
X_10376_ _04609_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12115_ fifo_bank_register.bank\[5\]\[125\] _05532_ _07198_ vssd1 vssd1 vccd1 vccd1
+ _07337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17972_ net434 _01415_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
X_13095_ _07855_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__clkbuf_1
X_16923_ net566 _00366_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
X_12046_ _07301_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16854_ net497 _00297_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _03834_ vssd1 vssd1 vccd1 vccd1 _01847_ sky130_fd_sc_hd__clkbuf_1
X_13997_ fifo_bank_register.bank\[1\]\[49\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[49\]
+ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a22o_1
X_16785_ clknet_leaf_80_clk _00229_ net578 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[76\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_217_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18524_ clknet_leaf_67_clk _01953_ net610 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_15736_ _03798_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__clkbuf_1
X_12948_ fifo_bank_register.bank\[1\]\[5\] _05280_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18455_ clknet_leaf_70_clk _01885_ net609 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[95\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15667_ mix1.data_o\[37\] net789 _03753_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__mux2_1
XANTENNA_170 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _07741_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_181 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_192 net118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17406_ net574 _00849_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14618_ fifo_bank_register.bank\[0\]\[117\] _02936_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15598_ mix1.data_o\[5\] _03382_ mix1.next_ready_o vssd1 vssd1 vccd1 vccd1 _03725_
+ sky130_fd_sc_hd__mux2_1
X_18386_ clknet_leaf_0_clk _01816_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[71\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17337_ net429 _00780_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
X_14549_ _02138_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17268_ net391 _00711_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16219_ net249 ks1.key_reg\[92\] _03979_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17199_ net467 _00642_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08972_ _04713_ _04994_ _04995_ _04716_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__a22o_1
XFILLER_0_227_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold18 mix1.data_reg\[116\] vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 ks1.key_reg\[14\] vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_194_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09524_ net239 vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09455_ _05398_ vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ _04518_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09386_ _05351_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08337_ _04482_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08268_ net139 net140 net138 net137 vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__and4b_1
XFILLER_0_166_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10230_ net199 ks1.key_reg\[47\] _05997_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ addroundkey_data_o\[39\] _05979_ _05980_ vssd1 vssd1 vccd1 vccd1 _05981_
+ sky130_fd_sc_hd__mux2_1
Xoutput380 net380 vssd1 vssd1 vccd1 vccd1 data_o[93] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10092_ mix1.data_o\[34\] _05576_ _05916_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__o21a_1
XFILLER_0_195_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13920_ _02151_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13851_ _02254_ fifo_bank_register.data_out\[32\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ fifo_bank_register.bank\[2\]\[64\] _05405_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13782_ fifo_bank_register.bank\[9\]\[25\] _02137_ _02190_ _02191_ _02192_ vssd1
+ vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__a2111o_1
X_16570_ net504 _00018_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_201_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10994_ net27 mix1.data_o\[123\] _05603_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15521_ sub1.data_o\[22\] sub1.data_o\[86\] _03671_ vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__mux2_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ fifo_bank_register.bank\[2\]\[31\] _05336_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18240_ clknet_leaf_39_clk _01671_ net663 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_15452_ _03632_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__clkbuf_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _05249_ _05250_ _07483_ net597 vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__and4b_1
XFILLER_0_182_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14403_ fifo_bank_register.bank\[9\]\[93\] _02712_ _02743_ _02744_ _02745_ vssd1
+ vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11615_ fifo_bank_register.bank\[6\]\[16\] _05303_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07074_ sky130_fd_sc_hd__mux2_1
X_15383_ sub1.data_o\[38\] sub1.data_o\[102\] _05202_ vssd1 vssd1 vccd1 vccd1 _03589_
+ sky130_fd_sc_hd__mux2_1
X_18171_ clknet_leaf_17_clk _01602_ net633 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12595_ _07591_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17122_ net485 _00565_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14334_ fifo_bank_register.bank\[6\]\[86\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[86\]
+ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11546_ _07037_ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17053_ net538 _00496_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14265_ _02622_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__clkbuf_1
X_11477_ fifo_bank_register.bank\[7\]\[79\] _05436_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _07001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16004_ net190 ks1.key_reg\[39\] _03910_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13216_ _07919_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10428_ _06219_ _06220_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__xor2_1
X_14196_ fifo_bank_register.bank\[9\]\[70\] _02550_ _02555_ _02558_ _02561_ vssd1
+ vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13147_ _07882_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10359_ net83 mix1.data_o\[59\] _06158_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ net399 _01398_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_13078_ _07846_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16906_ net511 _00349_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
X_12029_ _07292_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_174_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17886_ net482 _01329_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16837_ clknet_leaf_44_clk next_first_round_reg net663 vssd1 vssd1 vccd1 vccd1 first_round_reg
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16768_ clknet_leaf_47_clk _00212_ net651 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[59\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_220_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18507_ clknet_leaf_61_clk _01936_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_15719_ _03789_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16699_ clknet_leaf_72_clk _00146_ net635 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[126\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_111_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09240_ sub1.data_o\[119\] _05197_ _05246_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18438_ clknet_leaf_36_clk _01868_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[123\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09171_ _05180_ _05181_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18369_ clknet_leaf_37_clk _01799_ net666 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[54\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_6009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput108 data_i[81] vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_2
XTAP_5319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08955_ addroundkey_data_o\[87\] mix1.data_o\[87\] _04656_ vssd1 vssd1 vccd1 vccd1
+ _04979_ sky130_fd_sc_hd__mux2_1
Xinput119 data_i[91] vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_4
XFILLER_0_122_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08886_ _04653_ _04878_ _04896_ _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__a211o_2
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09507_ _05433_ vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09438_ fifo_bank_register.bank\[9\]\[55\] _05386_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05387_ sky130_fd_sc_hd__mux2_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ net184 vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ fifo_bank_register.bank\[7\]\[42\] _05359_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12380_ _05526_ fifo_bank_register.bank\[4\]\[122\] _07341_ vssd1 vssd1 vccd1 vccd1
+ _07477_ sky130_fd_sc_hd__mux2_1
XANTENNA_70 addroundkey_data_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_81 addroundkey_data_o\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11331_ _06912_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__buf_4
XANTENNA_92 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ _02431_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11262_ _05493_ fifo_bank_register.bank\[8\]\[106\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06887_ sky130_fd_sc_hd__mux2_1
X_13001_ _07794_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__buf_4
X_10213_ _06001_ _06025_ _06026_ _06005_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__a22o_1
X_11193_ _05424_ fifo_bank_register.bank\[8\]\[73\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10144_ _05899_ _05960_ _05964_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_101_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17740_ net477 _01183_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14952_ sub1.data_o\[17\] _04377_ _03081_ _03226_ vssd1 vssd1 vccd1 vccd1 _03227_
+ sky130_fd_sc_hd__a211o_1
X_10075_ sub1.data_o\[33\] _05900_ _05751_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ fifo_bank_register.bank\[5\]\[39\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[39\]
+ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a22o_1
X_17671_ net526 _01114_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
X_14883_ addroundkey_data_o\[103\] _03054_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_202_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16622_ net523 _00070_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_13834_ fifo_bank_register.bank\[0\]\[30\] _02238_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16553_ clknet_leaf_21_clk _00001_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[116\]
+ sky130_fd_sc_hd__dfrtp_4
X_13765_ fifo_bank_register.bank\[1\]\[23\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__a22o_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10977_ _06715_ vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__clkbuf_1
X_15504_ sub1.data_o\[49\] _03663_ _03666_ _03611_ vssd1 vssd1 vccd1 vccd1 _03667_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12716_ fifo_bank_register.bank\[2\]\[23\] _05319_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16484_ _04325_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__clkbuf_1
X_13696_ fifo_bank_register.bank\[6\]\[17\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__a22o_1
XFILLER_0_214_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18223_ clknet_leaf_37_clk _01654_ net666 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[53\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15435_ sub1.data_o\[23\] _03606_ _03623_ _03611_ vssd1 vssd1 vccd1 vccd1 _03624_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12647_ _07618_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15366_ _03577_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18154_ clknet_leaf_49_clk _01585_ net615 vssd1 vssd1 vccd1 vccd1 ks1.col\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12578_ _07582_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17105_ net535 _00548_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14317_ fifo_bank_register.bank\[7\]\[84\] _02623_ _02632_ fifo_bank_register.bank\[2\]\[84\]
+ _02668_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a221o_1
X_11529_ _07028_ vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__clkbuf_1
X_15297_ _03540_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__clkbuf_1
X_18085_ net542 _01528_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[87\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_1_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14248_ _02607_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__clkbuf_1
X_17036_ net518 _00479_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ fifo_bank_register.bank\[1\]\[69\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[69\]
+ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ addroundkey_data_o\[65\] mix1.data_o\[65\] _04655_ vssd1 vssd1 vccd1 vccd1
+ _04764_ sky130_fd_sc_hd__mux2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ net545 _01381_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08671_ _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__clkbuf_4
X_17869_ net425 _01312_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09223_ _05145_ _05171_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09154_ sbox1.ah_reg\[0\] _05119_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09085_ _05093_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput90 data_i[65] vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_4
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09987_ mix1.data_o\[23\] _05797_ _05821_ _05822_ sub1.data_o\[23\] vssd1 vssd1 vccd1
+ vccd1 _05823_ sky130_fd_sc_hd__a32o_1
XTAP_5127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08938_ ks1.key_reg\[29\] _04729_ _04731_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__or3_1
XTAP_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ addroundkey_data_o\[56\] mix1.data_o\[56\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04893_ sky130_fd_sc_hd__mux2_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ net145 ks1.key_reg\[113\] _04639_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__mux2_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11880_ fifo_bank_register.bank\[5\]\[13\] _05297_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10831_ net8 mix1.data_o\[106\] _06571_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13550_ _08120_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10762_ _05792_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12501_ _07508_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13481_ _05262_ fifo_bank_register.write_ptr\[2\] vssd1 vssd1 vccd1 vccd1 _08060_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10693_ _06457_ _06458_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__xor2_1
XFILLER_0_168_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15220_ _03466_ _03479_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12432_ _07505_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15151_ _03124_ _03179_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_106_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12363_ _07468_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14102_ _02151_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__buf_4
XFILLER_0_205_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ _06915_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__clkbuf_1
X_15082_ _03168_ _03353_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__xnor2_2
X_12294_ _07432_ vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ _02416_ fifo_bank_register.data_out\[52\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02417_ sky130_fd_sc_hd__mux2_1
X_11245_ _05476_ fifo_bank_register.bank\[8\]\[98\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11176_ _05407_ fifo_bank_register.bank\[8\]\[65\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10127_ _05574_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15984_ net188 ks1.key_reg\[37\] _03937_ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__mux2_1
XTAP_5661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17723_ net434 _01166_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14935_ sub1.data_o\[64\] _03209_ _03067_ sub1.data_o\[32\] vssd1 vssd1 vccd1 vccd1
+ _03210_ sky130_fd_sc_hd__a22o_1
X_10058_ net182 ks1.key_reg\[31\] _05825_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__mux2_2
XTAP_5694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17654_ net397 _01097_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14866_ _04617_ _03141_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__or2_1
XFILLER_0_159_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16605_ net405 _00053_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13817_ fifo_bank_register.bank\[0\]\[29\] _02223_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02224_ sky130_fd_sc_hd__mux2_1
X_17585_ net462 _01028_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14797_ addroundkey_data_o\[80\] _03072_ _03068_ addroundkey_data_o\[48\] vssd1 vssd1
+ vccd1 vccd1 _03073_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16536_ _04352_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__clkbuf_1
X_13748_ fifo_bank_register.bank\[6\]\[21\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16467_ _04185_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__inv_2
X_13679_ fifo_bank_register.bank\[7\]\[15\] _08182_ _08191_ fifo_bank_register.bank\[2\]\[15\]
+ _02099_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a221o_1
XFILLER_0_186_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18206_ clknet_leaf_18_clk _01637_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15418_ _03603_ _04949_ _05554_ _03612_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__a31o_1
XFILLER_0_183_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16398_ _04197_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18137_ clknet_leaf_53_clk sbox1.intermediate_to_invert_var\[3\] net656 vssd1 vssd1
+ vccd1 vccd1 sbox1.inversion_to_invert_var\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15349_ _03567_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 mix1.data_reg\[123\] vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold115 mix1.data_reg\[89\] vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18068_ net516 _01511_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[70\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold126 ks1.key_reg\[76\] vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 ks1.key_reg\[56\] vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold148 ks1.key_reg\[45\] vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09910_ _05613_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold159 ks1.key_reg\[71\] vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ net562 _00462_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout606 net607 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
X_09841_ sub1.data_o\[9\] _05690_ _05610_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout617 net618 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout628 net634 vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
Xfanout639 net640 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__clkbuf_2
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09772_ net40 mix1.data_o\[1\] _05604_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__mux2_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ ks1.key_reg\[28\] _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__or3_1
XFILLER_0_193_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08654_ addroundkey_data_o\[84\] mix1.data_o\[84\] _04663_ vssd1 vssd1 vccd1 vccd1
+ _04678_ sky130_fd_sc_hd__mux2_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08585_ round\[0\] vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__buf_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09206_ _05153_ _05214_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09137_ _05146_ _05147_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__xor2_4
X_09068_ _05016_ sbox1.ah\[0\] _05071_ sbox1.ah\[1\] vssd1 vssd1 vccd1 vccd1 _05082_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_130_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11030_ net160 ks1.key_reg\[127\] _05762_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_216_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ fifo_bank_register.bank\[1\]\[20\] _05311_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ sub1.data_o\[85\] _03010_ _03022_ sub1.next_ready_o vssd1 vssd1 vccd1 vccd1
+ _03023_ sky130_fd_sc_hd__a22o_1
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _07241_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__clkbuf_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ fifo_bank_register.bank\[5\]\[5\] _05280_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07205_ sky130_fd_sc_hd__mux2_1
X_14651_ fifo_bank_register.bank\[0\]\[121\] _02965_ _08120_ vssd1 vssd1 vccd1 vccd1
+ _02966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ fifo_bank_register.bank\[5\]\[7\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[7\]
+ vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _06567_ _06568_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__xor2_1
XFILLER_0_200_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17370_ net501 _00813_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14582_ fifo_bank_register.bank\[7\]\[113\] _02866_ _02875_ fifo_bank_register.bank\[2\]\[113\]
+ _02904_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11794_ _07168_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16321_ net672 _04136_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__nand2_1
X_10745_ sub1.data_o\[98\] _06341_ _06504_ _06505_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06506_ sky130_fd_sc_hd__a221o_1
X_13533_ _08103_ vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13464_ _08049_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__clkbuf_1
X_16252_ net252 ks1.key_reg\[95\] _03979_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__mux2_2
XFILLER_0_192_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10676_ net248 ks1.key_reg\[91\] _06324_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_200_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15203_ _03138_ _03465_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__xnor2_4
X_12415_ _07496_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13395_ _08013_ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__clkbuf_1
X_16183_ net210 ks1.key_reg\[57\] _03937_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__mux2_1
X_15134_ net720 _03402_ _03171_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__mux2_1
X_12346_ _07459_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15065_ sub1.data_o\[84\] _03072_ _03068_ sub1.data_o\[52\] vssd1 vssd1 vccd1 vccd1
+ _03337_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12277_ _07423_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ fifo_bank_register.bank\[0\]\[50\] _02400_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02402_ sky130_fd_sc_hd__mux2_1
X_11228_ _06791_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__buf_4
XFILLER_0_226_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ _05390_ fifo_bank_register.bank\[8\]\[57\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ _03936_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__xor2_2
XTAP_5491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_164_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17706_ net452 _01149_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
X_14918_ addroundkey_data_o\[14\] _03100_ _05606_ _03192_ vssd1 vssd1 vccd1 vccd1
+ _03193_ sky130_fd_sc_hd__a211o_1
XTAP_4790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15898_ sub1.data_o\[100\] _03884_ _03876_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17637_ net423 _01080_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14849_ sub1.data_o\[69\] _03108_ _03066_ sub1.data_o\[37\] vssd1 vssd1 vccd1 vccd1
+ _03125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08370_ _04499_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17568_ net402 _01011_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16519_ net688 _03502_ _04343_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17499_ net485 _00942_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_2__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_171_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout403 net404 vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__buf_1
Xfanout414 net419 vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__buf_2
Xfanout425 net427 vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_2
Xfanout436 net444 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_2
X_09824_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__buf_4
Xfanout447 net449 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout458 net460 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_2
Xfanout469 net470 vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_214_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09755_ _04627_ _05613_ _04609_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_216_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08706_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__buf_2
X_09686_ _05153_ _05243_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__xnor2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__clkbuf_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ addroundkey_data_o\[122\] fifo_bank_register.data_out\[122\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08499_ _04478_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__buf_6
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10530_ mix1.data_o\[78\] _06296_ _06241_ _06242_ sub1.data_o\[78\] vssd1 vssd1 vccd1
+ vccd1 _06311_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10461_ _05614_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12200_ _05346_ fifo_bank_register.bank\[4\]\[36\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13180_ fifo_bank_register.bank\[1\]\[115\] _05512_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07900_ sky130_fd_sc_hd__mux2_1
X_10392_ mix1.data_o\[62\] _06138_ _06162_ _06163_ sub1.data_o\[62\] vssd1 vssd1 vccd1
+ vccd1 _06189_ sky130_fd_sc_hd__a32o_1
XFILLER_0_27_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12131_ _07346_ vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12062_ _07309_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11013_ _05615_ _06745_ _06746_ _05567_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__a22o_1
X_16870_ net417 _00313_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ mix1.data_o\[110\] net711 _03841_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__mux2_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18540_ clknet_leaf_66_clk _01969_ net606 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[67\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _03806_ vssd1 vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__clkbuf_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12964_ _07786_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__clkbuf_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14703_ sub1.data_o\[48\] sub1.data_o\[112\] _05598_ vssd1 vssd1 vccd1 vccd1 _03011_
+ sky130_fd_sc_hd__mux2_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18471_ clknet_leaf_83_clk _01901_ net584 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[111\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _07232_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15683_ _03770_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__clkbuf_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_330 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _07749_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_341 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_352 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17422_ net553 _00865_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
X_14634_ fifo_bank_register.bank\[9\]\[119\] _02874_ _02948_ _02949_ _02950_ vssd1
+ vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__a2111o_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ fifo_bank_register.bank\[6\]\[126\] _05534_ _07055_ vssd1 vssd1 vccd1 vccd1
+ _07195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17353_ net473 _00796_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14565_ fifo_bank_register.bank\[5\]\[111\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[111\]
+ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__a22o_1
X_11777_ _07159_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _04226_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__clkbuf_1
X_10728_ sub1.data_o\[97\] _06489_ _06478_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__mux2_1
X_13516_ _05262_ _08065_ vssd1 vssd1 vccd1 vccd1 _08087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17284_ net521 _00727_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14496_ _02828_ fifo_bank_register.data_out\[103\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16235_ ks1.key_reg\[29\] _04180_ _04106_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ net245 ks1.key_reg\[89\] _06324_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__mux2_1
X_13447_ _05508_ fifo_bank_register.bank\[0\]\[113\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13378_ _05438_ fifo_bank_register.bank\[0\]\[80\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08005_ sky130_fd_sc_hd__mux2_1
X_16166_ _04115_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__xor2_2
XFILLER_0_224_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15117_ _03354_ _03386_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ _07450_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16097_ net201 ks1.key_reg\[49\] _03937_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15048_ _03317_ _03320_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__nor2_8
XFILLER_0_227_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16999_ net424 _00442_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09540_ fifo_bank_register.bank\[9\]\[88\] _05455_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09471_ net220 vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__buf_2
XFILLER_0_222_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08422_ addroundkey_data_o\[52\] fifo_bank_register.data_out\[52\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__mux2_2
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08353_ addroundkey_data_o\[19\] fifo_bank_register.data_out\[19\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__mux2_2
XFILLER_0_163_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08284_ _04439_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09807_ mix1.data_o\[5\] _05586_ _05618_ _05621_ sub1.data_o\[5\] vssd1 vssd1 vccd1
+ vccd1 _05661_ sky130_fd_sc_hd__a32o_1
XFILLER_0_214_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09738_ _05202_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09669_ addroundkey_round\[2\] _04637_ _04642_ _05542_ vssd1 vssd1 vccd1 vccd1 _00138_
+ sky130_fd_sc_hd__a31o_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ fifo_bank_register.bank\[6\]\[56\] _05388_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07119_ sky130_fd_sc_hd__mux2_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12680_ _07636_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__clkbuf_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11631_ fifo_bank_register.bank\[6\]\[23\] _05319_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07083_ sky130_fd_sc_hd__mux2_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14350_ fifo_bank_register.bank\[7\]\[88\] _02623_ _02632_ fifo_bank_register.bank\[2\]\[88\]
+ _02697_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a221o_1
X_11562_ _07045_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10513_ _05585_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__clkbuf_4
X_13301_ _07964_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14281_ _02146_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11493_ _07009_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__clkbuf_1
X_13232_ _05293_ fifo_bank_register.bank\[0\]\[11\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07928_ sky130_fd_sc_hd__mux2_1
X_16020_ _03986_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ _06233_ _06234_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13163_ fifo_bank_register.bank\[1\]\[107\] _05495_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07891_ sky130_fd_sc_hd__mux2_1
X_10375_ mix1.data_o\[60\] _06138_ _06162_ _06163_ sub1.data_o\[60\] vssd1 vssd1 vccd1
+ vccd1 _06174_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ _07336_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13094_ fifo_bank_register.bank\[1\]\[74\] _05426_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07855_ sky130_fd_sc_hd__mux2_1
X_17971_ net458 _01414_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12045_ fifo_bank_register.bank\[5\]\[91\] _05462_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07301_ sky130_fd_sc_hd__mux2_1
X_16922_ net548 _00365_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16853_ net505 _00296_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_15804_ mix1.data_o\[102\] net717 _03830_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16784_ clknet_leaf_73_clk _00228_ net593 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[75\]
+ sky130_fd_sc_hd__dfrtp_4
X_13996_ fifo_bank_register.bank\[6\]\[49\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[49\]
+ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18523_ clknet_leaf_67_clk _01952_ net606 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15735_ mix1.data_o\[69\] net750 _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12947_ _07777_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__clkbuf_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ clknet_leaf_72_clk _01884_ net594 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[94\]
+ sky130_fd_sc_hd__dfrtp_1
X_15666_ _03761_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12878_ fifo_bank_register.bank\[2\]\[100\] _05480_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07741_ sky130_fd_sc_hd__mux2_1
XANTENNA_171 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_182 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17405_ net574 _00848_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_193 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617_ fifo_bank_register.bank\[9\]\[117\] _02874_ _02933_ _02934_ _02935_ vssd1
+ vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_157_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18385_ clknet_leaf_12_clk _01815_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[70\]
+ sky130_fd_sc_hd__dfrtp_4
X_11829_ _07186_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__clkbuf_1
X_15597_ _03724_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__clkbuf_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ net408 _00779_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
X_14548_ _02136_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17267_ net394 _00710_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_14479_ fifo_bank_register.bank\[0\]\[101\] _02813_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16218_ _04163_ _04164_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17198_ net463 _00641_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16149_ net243 ks1.key_reg\[87\] _03906_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ addroundkey_data_o\[95\] mix1.data_o\[95\] _04663_ vssd1 vssd1 vccd1 vccd1
+ _04995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold19 ks1.key_reg\[30\] vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09523_ _05444_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09454_ fifo_bank_register.bank\[9\]\[60\] _05396_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08405_ addroundkey_data_o\[44\] fifo_bank_register.data_out\[44\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__mux2_2
XFILLER_0_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09385_ fifo_bank_register.bank\[9\]\[38\] _05350_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08336_ addroundkey_data_o\[11\] fifo_bank_register.data_out\[11\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__mux2_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08267_ _04420_ _04421_ _04422_ _04423_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10160_ _05792_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput370 net370 vssd1 vssd1 vccd1 vccd1 data_o[84] sky130_fd_sc_hd__clkbuf_4
Xoutput381 net381 vssd1 vssd1 vccd1 vccd1 data_o[94] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10091_ _05757_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13850_ fifo_bank_register.bank\[0\]\[32\] _02253_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _07700_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__clkbuf_1
X_13781_ fifo_bank_register.bank\[1\]\[25\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__a22o_1
X_10993_ _06729_ vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15520_ _03668_ _04777_ _05228_ _03678_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a31o_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _07664_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_214_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15451_ sub1.data_o\[31\] _05244_ _04879_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__mux2_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _07626_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ fifo_bank_register.bank\[1\]\[93\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[93\]
+ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__a22o_1
X_18170_ clknet_leaf_11_clk _01601_ net631 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_11614_ _07073_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15382_ _03588_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__clkbuf_1
X_12594_ fifo_bank_register.bank\[3\]\[94\] _05468_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17121_ net499 _00564_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14333_ fifo_bank_register.bank\[7\]\[86\] _02623_ _02632_ fifo_bank_register.bank\[2\]\[86\]
+ _02682_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11545_ fifo_bank_register.bank\[7\]\[111\] _05504_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17052_ net536 _00495_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11476_ _07000_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__clkbuf_1
X_14264_ _02621_ fifo_bank_register.data_out\[78\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16003_ _03969_ _03970_ vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__xor2_4
X_13215_ _05276_ fifo_bank_register.bank\[0\]\[3\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07919_ sky130_fd_sc_hd__mux2_1
X_10427_ net220 ks1.key_reg\[66\] _06166_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14195_ fifo_bank_register.bank\[1\]\[70\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[70\]
+ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10358_ _05603_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ fifo_bank_register.bank\[1\]\[99\] _05478_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07882_ sky130_fd_sc_hd__mux2_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ fifo_bank_register.bank\[1\]\[66\] _05409_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07846_ sky130_fd_sc_hd__mux2_1
X_17954_ net410 _01397_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
X_10289_ _06076_ _06089_ _06095_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_40_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16905_ net509 _00348_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_12028_ fifo_bank_register.bank\[5\]\[83\] _05445_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17885_ net483 _01328_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16836_ clknet_leaf_69_clk _00280_ net608 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[127\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16767_ clknet_leaf_68_clk _00211_ net611 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[58\]
+ sky130_fd_sc_hd__dfrtp_4
X_13979_ fifo_bank_register.bank\[1\]\[47\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[47\]
+ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18506_ clknet_leaf_59_clk _01935_ net606 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15718_ mix1.data_o\[61\] net724 _03786_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16698_ clknet_leaf_71_clk _00145_ net652 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18437_ clknet_leaf_24_clk _01867_ net645 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[122\]
+ sky130_fd_sc_hd__dfrtp_4
X_15649_ _03752_ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_173_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_158_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09170_ sbox1.ah_reg\[1\] _05142_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18368_ clknet_leaf_37_clk _01798_ net666 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[53\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17319_ net448 _00762_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18299_ clknet_leaf_29_clk _01730_ net642 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[65\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08954_ _04670_ _04976_ _04977_ _04675_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a22o_1
Xinput109 data_i[82] vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_4
XFILLER_0_122_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08885_ _04899_ _04902_ _04905_ _04908_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__or4_1
XFILLER_0_192_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09506_ fifo_bank_register.bank\[9\]\[77\] _05432_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ net208 vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__clkbuf_4
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09368_ _05339_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08319_ _04472_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_164_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09299_ _05292_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_60 addroundkey_data_o\[19\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 addroundkey_data_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_82 addroundkey_data_o\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _06923_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_93 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ _06886_ vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10212_ mix1.data_o\[45\] _05876_ _05993_ _05994_ sub1.data_o\[45\] vssd1 vssd1 vccd1
+ vccd1 _06026_ sky130_fd_sc_hd__a32o_1
X_13000_ _07805_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__clkbuf_1
X_11192_ _06850_ vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10143_ sub1.data_o\[38\] _05753_ _05962_ _05963_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _05964_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14951_ sub1.data_o\[81\] _03209_ _03067_ sub1.data_o\[49\] vssd1 vssd1 vccd1 vccd1
+ _03226_ sky130_fd_sc_hd__a22o_1
X_10074_ net55 mix1.data_o\[33\] _05749_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__mux2_1
XTAP_5854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13902_ _08181_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__clkbuf_4
XTAP_5887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17670_ net512 _01113_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14882_ addroundkey_data_o\[7\] _04374_ _04900_ _03157_ vssd1 vssd1 vccd1 vccd1 _03158_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_215_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16621_ net527 _00069_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13833_ _02157_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__buf_4
XFILLER_0_187_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16552_ clknet_leaf_28_clk _00000_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[115\]
+ sky130_fd_sc_hd__dfrtp_4
X_13764_ fifo_bank_register.bank\[6\]\[23\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__a22o_1
X_10976_ addroundkey_data_o\[120\] _06714_ _05696_ vssd1 vssd1 vccd1 vccd1 _06715_
+ sky130_fd_sc_hd__mux2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15503_ sub1.data_o\[17\] sub1.data_o\[81\] _03609_ vssd1 vssd1 vccd1 vccd1 _03666_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12715_ _07655_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16483_ net719 _03324_ _04321_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13695_ fifo_bank_register.bank\[7\]\[17\] _08182_ _08191_ fifo_bank_register.bank\[2\]\[17\]
+ _02113_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a221o_1
X_18222_ clknet_leaf_37_clk _01653_ net666 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[52\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15434_ sub1.data_o\[119\] sub1.data_o\[55\] _03609_ vssd1 vssd1 vccd1 vccd1 _03623_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ fifo_bank_register.bank\[3\]\[119\] _05520_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18153_ clknet_leaf_81_clk _01584_ net578 vssd1 vssd1 vccd1 vccd1 ks1.col\[7\] sky130_fd_sc_hd__dfrtp_4
X_15365_ sub1.data_o\[0\] _03575_ _03576_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12577_ fifo_bank_register.bank\[3\]\[86\] _05451_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17104_ net504 _00547_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ fifo_bank_register.bank\[5\]\[84\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[84\]
+ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11528_ fifo_bank_register.bank\[7\]\[103\] _05487_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07028_ sky130_fd_sc_hd__mux2_1
X_18084_ net560 _01527_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[86\]
+ sky130_fd_sc_hd__dfxtp_2
X_15296_ net694 _03170_ _03539_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17035_ net516 _00478_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
X_14247_ _02606_ fifo_bank_register.data_out\[76\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02607_ sky130_fd_sc_hd__mux2_1
X_11459_ fifo_bank_register.bank\[7\]\[70\] _05417_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _06992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14178_ fifo_bank_register.bank\[6\]\[69\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[69\]
+ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__a22o_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _07873_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__clkbuf_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ net552 _01380_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08670_ sub1.state\[2\] _04687_ _04364_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__and3b_2
XFILLER_0_79_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17868_ net425 _01311_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16819_ clknet_leaf_4_clk _00263_ net591 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[110\]
+ sky130_fd_sc_hd__dfrtp_4
X_17799_ net518 _01242_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09222_ _05104_ _04946_ _05228_ _05230_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09153_ sbox1.ah_reg\[3\] _05134_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__nand2_2
XFILLER_0_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _05095_ _05096_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__xor2_1
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput80 data_i[56] vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_4
Xinput91 data_i[66] vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__buf_4
XFILLER_0_226_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09986_ _05620_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__buf_2
XFILLER_0_228_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08937_ ks1.key_reg\[5\] _04735_ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08868_ _04888_ _04889_ _04890_ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08799_ addroundkey_data_o\[99\] mix1.data_o\[99\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _04823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10830_ _05614_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10761_ _06519_ _06520_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_211_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12500_ _07541_ vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13480_ _05262_ fifo_bank_register.write_ptr\[2\] vssd1 vssd1 vccd1 vccd1 _08059_
+ sky130_fd_sc_hd__or2_1
X_10692_ net250 ks1.key_reg\[93\] _06324_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12431_ fifo_bank_register.bank\[3\]\[17\] _05305_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15150_ _03167_ _03416_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__xor2_4
XFILLER_0_168_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ _05508_ fifo_bank_register.bank\[4\]\[113\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14101_ fifo_bank_register.bank\[6\]\[60\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[60\]
+ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a22o_1
X_11313_ fifo_bank_register.bank\[7\]\[1\] _05272_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06915_ sky130_fd_sc_hd__mux2_1
X_15081_ _03314_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__xnor2_4
X_12293_ _05438_ fifo_bank_register.bank\[4\]\[80\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14032_ fifo_bank_register.bank\[0\]\[52\] _02415_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02416_ sky130_fd_sc_hd__mux2_1
X_11244_ _06877_ vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ _06841_ vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10126_ sub1.data_o\[37\] _05947_ _05936_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15983_ _03951_ _03952_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__xor2_4
XFILLER_0_175_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17722_ net412 _01165_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14934_ _03108_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__buf_4
X_10057_ _05829_ _05883_ _05884_ _05833_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a22o_1
XTAP_5684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ net396 _01096_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865_ _03117_ _03140_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__xor2_4
XFILLER_0_203_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ net389 _00052_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_13816_ fifo_bank_register.bank\[9\]\[29\] _02137_ _02220_ _02221_ _02222_ vssd1
+ vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17584_ net462 _01027_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14796_ _03064_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__buf_4
XFILLER_0_212_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16535_ net766 _03527_ _04343_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13747_ fifo_bank_register.bank\[7\]\[21\] _02128_ _02139_ fifo_bank_register.bank\[2\]\[21\]
+ _02161_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__a221o_1
X_10959_ net22 mix1.data_o\[119\] _05602_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16466_ _04315_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13678_ fifo_bank_register.bank\[5\]\[15\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18205_ clknet_leaf_18_clk _01636_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_15417_ sub1.data_o\[17\] _03606_ _03610_ _03611_ vssd1 vssd1 vccd1 vccd1 _03612_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12629_ _07609_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16397_ _04277_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18136_ clknet_leaf_53_clk sbox1.intermediate_to_invert_var\[2\] net656 vssd1 vssd1
+ vccd1 vccd1 sbox1.inversion_to_invert_var\[2\] sky130_fd_sc_hd__dfrtp_1
X_15348_ net715 _03516_ _03560_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold105 mix1.data_reg\[85\] vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18067_ net516 _01510_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[69\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_223_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold116 mix1.data_reg\[83\] vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ _03452_ _03472_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold127 ks1.key_reg\[107\] vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold138 ks1.key_reg\[83\] vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17018_ net563 _00461_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold149 ks1.key_reg\[124\] vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_223_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1094 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09840_ net128 mix1.data_o\[9\] _05604_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__mux2_1
Xfanout607 net617 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__buf_2
Xfanout618 net259 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__buf_2
Xfanout629 net630 vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ _05615_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__clkbuf_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _04731_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__buf_2
XFILLER_0_217_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08653_ _04362_ _04364_ _04365_ _04363_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_96_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08584_ _04612_ vssd1 vssd1 vccd1 vccd1 next_first_round_reg sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09205_ _05163_ _05184_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09136_ sbox1.alph\[3\] _05127_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__nand2_2
XFILLER_0_228_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _05075_ _05081_ vssd1 vssd1 vccd1 vccd1 sbox1.intermediate_to_invert_var\[3\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ net171 ks1.key_reg\[21\] _05708_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__mux2_2
XFILLER_0_228_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__buf_4
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ fifo_bank_register.bank\[5\]\[37\] _05348_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07241_ sky130_fd_sc_hd__mux2_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ fifo_bank_register.bank\[9\]\[121\] _08089_ _02962_ _02963_ _02964_ vssd1
+ vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__a2111o_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11862_ _07204_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__clkbuf_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _08165_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ net135 ks1.key_reg\[104\] _06324_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__mux2_1
X_14581_ fifo_bank_register.bank\[5\]\[113\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[113\]
+ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__a22o_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ fifo_bank_register.bank\[6\]\[100\] _05480_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07168_ sky130_fd_sc_hd__mux2_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16320_ _04215_ _04169_ _04234_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13532_ _08066_ _08094_ vssd1 vssd1 vccd1 vccd1 _08103_ sky130_fd_sc_hd__nor2_1
X_10744_ mix1.data_o\[98\] _06494_ _06398_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16251_ _04193_ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__xnor2_4
X_13463_ _05524_ fifo_bank_register.bank\[0\]\[121\] _07914_ vssd1 vssd1 vccd1 vccd1
+ _08049_ sky130_fd_sc_hd__mux2_1
X_10675_ _06416_ _06441_ _06442_ _06420_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15202_ _03361_ _03371_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ fifo_bank_register.bank\[3\]\[9\] _05288_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16182_ _04130_ _04131_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__xor2_4
X_13394_ _05455_ fifo_bank_register.bank\[0\]\[88\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15133_ _03394_ _03401_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_129_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12345_ _05491_ fifo_bank_register.bank\[4\]\[105\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15064_ _03332_ _03335_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__nor2_8
XFILLER_0_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12276_ _05422_ fifo_bank_register.bank\[4\]\[72\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14015_ _02157_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__buf_4
X_11227_ _06868_ vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ _06832_ vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10109_ addroundkey_data_o\[35\] _05932_ _05872_ vssd1 vssd1 vccd1 vccd1 _05933_
+ sky130_fd_sc_hd__mux2_1
X_11089_ _06796_ vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__clkbuf_1
X_15966_ net186 ks1.key_reg\[35\] _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__mux2_1
XTAP_5470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14917_ addroundkey_data_o\[78\] _03108_ _03066_ addroundkey_data_o\[46\] vssd1 vssd1
+ vccd1 vccd1 _03192_ sky130_fd_sc_hd__a22o_1
X_17705_ net446 _01148_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15897_ _05218_ sub1.data_o\[68\] _05200_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14848_ _03120_ _03123_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__nor2_8
X_17636_ net418 _01079_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17567_ net536 _01010_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
X_14779_ _03054_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__buf_6
XFILLER_0_105_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ _03143_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17498_ net501 _00941_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16449_ net801 _04100_ _04295_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18119_ net490 _01562_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_197_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout404 net444 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_2
Xfanout415 net419 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout426 net427 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_2
X_09823_ _05584_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__clkbuf_4
Xfanout437 net443 vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__buf_2
Xfanout448 net449 vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_2
Xfanout459 net460 vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__buf_1
XFILLER_0_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09754_ _05612_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08705_ _04728_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_213_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09685_ _05555_ vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__clkbuf_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ sub1.state\[1\] _04363_ sub1.state\[3\] sub1.state\[2\] vssd1 vssd1 vccd1
+ vccd1 _04660_ sky130_fd_sc_hd__and4b_1
XFILLER_0_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08567_ _04602_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__buf_1
XFILLER_0_193_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08498_ _04566_ vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10460_ _06249_ vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ sbox1.inversion_to_invert_var\[1\] _05105_ sbox1.inversion_to_invert_var\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10391_ sub1.data_o\[62\] _06187_ _06160_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12130_ _05276_ fifo_bank_register.bank\[4\]\[3\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ fifo_bank_register.bank\[5\]\[99\] _05478_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11012_ mix1.data_o\[125\] _05676_ _05758_ _05620_ sub1.data_o\[125\] vssd1 vssd1
+ vccd1 vccd1 _06746_ sky130_fd_sc_hd__a32o_1
XFILLER_0_99_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15820_ _03842_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15751_ mix1.data_o\[77\] net780 _03797_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__mux2_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12963_ fifo_bank_register.bank\[1\]\[12\] _05295_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07786_ sky130_fd_sc_hd__mux2_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_clk clknet_3_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _04369_ _04927_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__nor2_4
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18470_ clknet_leaf_3_clk _01900_ net583 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[110\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ fifo_bank_register.bank\[5\]\[29\] _05331_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07232_ sky130_fd_sc_hd__mux2_1
X_15682_ mix1.data_o\[44\] net767 _03764_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__mux2_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_320 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12894_ fifo_bank_register.bank\[2\]\[108\] _05497_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07749_ sky130_fd_sc_hd__mux2_1
XANTENNA_331 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_342 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ net525 _00864_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14633_ fifo_bank_register.bank\[1\]\[119\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[119\]
+ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__a22o_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_353 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11845_ _07194_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__clkbuf_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17352_ net474 _00795_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _02889_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__clkbuf_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ fifo_bank_register.bank\[6\]\[92\] _05464_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16303_ ks1.key_reg\[52\] _04080_ _04222_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13515_ _08086_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10727_ net125 mix1.data_o\[97\] _06476_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17283_ net526 _00726_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14495_ fifo_bank_register.bank\[0\]\[103\] _02827_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16234_ _04963_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__xnor2_1
X_13446_ _08040_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__clkbuf_1
X_10658_ _06416_ _06426_ _06427_ _06420_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__a22o_2
XFILLER_0_183_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16165_ net153 ks1.key_reg\[120\] _03976_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13377_ _07937_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__buf_4
X_10589_ mix1.data_o\[83\] _06129_ _06093_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15116_ _03343_ _03371_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_51_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12328_ _05474_ fifo_bank_register.bank\[4\]\[97\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07450_ sky130_fd_sc_hd__mux2_1
X_16096_ _04052_ _04053_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__xor2_4
XFILLER_0_220_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ addroundkey_data_o\[107\] _03079_ _03319_ vssd1 vssd1 vccd1 vccd1 _03320_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_43_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12259_ _05405_ fifo_bank_register.bank\[4\]\[64\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16998_ net414 _00441_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_15949_ _04759_ _03922_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__and2_1
XFILLER_0_211_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09470_ _05408_ vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__clkbuf_1
X_08421_ _04526_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__buf_1
XFILLER_0_8_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17619_ net505 _01062_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18599_ clknet_leaf_68_clk _02028_ net608 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[126\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_176_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08352_ _04478_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08283_ net235 net224 net257 net246 vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__and4b_1
XFILLER_0_74_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09806_ sub1.data_o\[5\] _05659_ _05610_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09737_ round\[3\] _05587_ _05596_ _05576_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_214_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09668_ _04644_ _05540_ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__nor3_2
XFILLER_0_97_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08619_ _04637_ _04636_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__or2b_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ fifo_bank_register.bank\[9\]\[107\] _05495_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05496_ sky130_fd_sc_hd__mux2_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11630_ _07082_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ fifo_bank_register.bank\[7\]\[119\] _05520_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13300_ _05361_ fifo_bank_register.bank\[0\]\[43\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07964_ sky130_fd_sc_hd__mux2_1
X_10512_ sub1.data_o\[76\] _06294_ _06239_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14280_ fifo_bank_register.bank\[7\]\[80\] _02623_ _02632_ fifo_bank_register.bank\[2\]\[80\]
+ _02635_ vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__a221o_1
XFILLER_0_208_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11492_ fifo_bank_register.bank\[7\]\[86\] _05451_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13231_ _07927_ vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10443_ net222 ks1.key_reg\[68\] _06166_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ _07890_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__clkbuf_1
X_10374_ sub1.data_o\[60\] _06172_ _06160_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12113_ fifo_bank_register.bank\[5\]\[124\] _05530_ _07198_ vssd1 vssd1 vccd1 vccd1
+ _07336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13093_ _07854_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__clkbuf_1
X_17970_ net452 _01413_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
X_12044_ _07300_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__clkbuf_1
X_16921_ net561 _00364_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16852_ net534 _00295_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15803_ _03833_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__clkbuf_1
X_16783_ clknet_leaf_74_clk _00227_ net591 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13995_ fifo_bank_register.bank\[7\]\[49\] _02380_ _02308_ fifo_bank_register.bank\[2\]\[49\]
+ _02381_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a221o_1
XFILLER_0_205_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_57_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15734_ _03741_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18522_ clknet_leaf_67_clk _01951_ net606 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
X_12946_ fifo_bank_register.bank\[1\]\[4\] _05278_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07777_ sky130_fd_sc_hd__mux2_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15665_ mix1.data_o\[36\] net700 _03753_ vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__mux2_1
X_18453_ clknet_leaf_70_clk _01883_ net609 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[93\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_150 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _07651_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_161 net94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_172 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14616_ fifo_bank_register.bank\[1\]\[117\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[117\]
+ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__a22o_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ net556 _00847_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18384_ clknet_leaf_12_clk _01814_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[69\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11828_ fifo_bank_register.bank\[6\]\[117\] _05516_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07186_ sky130_fd_sc_hd__mux2_1
XANTENNA_183 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15596_ mix1.data_o\[4\] _03363_ mix1.next_ready_o vssd1 vssd1 vccd1 vccd1 _03724_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_194 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ net429 _00778_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14547_ _02873_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__clkbuf_1
X_11759_ fifo_bank_register.bank\[6\]\[84\] _05447_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17266_ net391 _00709_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
X_14478_ fifo_bank_register.bank\[9\]\[101\] _02793_ _02810_ _02811_ _02812_ vssd1
+ vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_102_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16217_ net157 ks1.key_reg\[124\] _03976_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__mux2_2
XFILLER_0_148_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13429_ _08031_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17197_ net467 _00640_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16148_ ks1.col\[23\] _04099_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08970_ addroundkey_data_o\[71\] mix1.data_o\[71\] _04778_ vssd1 vssd1 vccd1 vccd1
+ _04994_ sky130_fd_sc_hd__mux2_1
X_16079_ _04036_ _04038_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_227_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 data_i[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_4
XFILLER_0_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09522_ fifo_bank_register.bank\[9\]\[82\] _05443_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05444_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09453_ _05312_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08404_ _04517_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09384_ net189 vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08335_ _04481_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08266_ net62 net51 net84 net73 vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__or4_1
XFILLER_0_85_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput360 net360 vssd1 vssd1 vccd1 vccd1 data_o[75] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput371 net371 vssd1 vssd1 vccd1 vccd1 data_o[85] sky130_fd_sc_hd__buf_2
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput382 net382 vssd1 vssd1 vccd1 vccd1 data_o[95] sky130_fd_sc_hd__clkbuf_4
X_10090_ _05575_ _05912_ _05914_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__a21o_1
XFILLER_0_203_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_39_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12800_ fifo_bank_register.bank\[2\]\[63\] _05403_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13780_ fifo_bank_register.bank\[6\]\[25\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__a22o_1
X_10992_ addroundkey_data_o\[122\] _06728_ _05696_ vssd1 vssd1 vccd1 vccd1 _06729_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ fifo_bank_register.bank\[2\]\[30\] _05333_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15450_ _03631_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__clkbuf_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12662_ fifo_bank_register.bank\[3\]\[127\] _05536_ _07485_ vssd1 vssd1 vccd1 vccd1
+ _07626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401_ fifo_bank_register.bank\[6\]\[93\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[93\]
+ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__a22o_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ fifo_bank_register.bank\[6\]\[15\] _05301_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07073_ sky130_fd_sc_hd__mux2_1
X_15381_ sub1.data_o\[5\] _03587_ _03581_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12593_ _07590_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__clkbuf_1
X_17120_ net510 _00563_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14332_ fifo_bank_register.bank\[5\]\[86\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[86\]
+ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a22o_1
X_11544_ _07036_ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17051_ net540 _00494_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14263_ fifo_bank_register.bank\[0\]\[78\] _02620_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02621_ sky130_fd_sc_hd__mux2_1
X_11475_ fifo_bank_register.bank\[7\]\[78\] _05434_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _07000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16002_ net226 ks1.key_reg\[71\] _03907_ vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__mux2_2
XFILLER_0_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ _07918_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10426_ _06171_ _06216_ _06218_ _06175_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14194_ _02153_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13145_ _07881_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10357_ _06157_ vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _07845_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__clkbuf_1
X_17953_ net403 _01396_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10288_ sub1.data_o\[52\] _05971_ _06092_ _06094_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _06095_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16904_ net526 _00347_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
X_12027_ _07291_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17884_ net502 _01327_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16835_ clknet_leaf_68_clk _00279_ net608 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[126\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_178_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16766_ clknet_leaf_48_clk _00210_ net610 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[57\]
+ sky130_fd_sc_hd__dfrtp_4
X_13978_ fifo_bank_register.bank\[6\]\[47\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[47\]
+ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18505_ clknet_leaf_58_clk _01934_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_15717_ _03788_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__clkbuf_1
X_12929_ fifo_bank_register.bank\[2\]\[125\] _05532_ _07628_ vssd1 vssd1 vccd1 vccd1
+ _07767_ sky130_fd_sc_hd__mux2_1
X_16697_ clknet_leaf_71_clk _00144_ net608 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[124\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_220_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18436_ clknet_leaf_25_clk _01866_ net650 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[121\]
+ sky130_fd_sc_hd__dfrtp_4
X_15648_ mix1.data_o\[28\] _03527_ _03742_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18367_ clknet_leaf_37_clk _01797_ net667 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[52\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_173_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15579_ sub1.data_o\[12\] _03660_ _03710_ sub1.data_o\[76\] vssd1 vssd1 vccd1 vccd1
+ _03715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17318_ net401 _00761_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
X_18298_ clknet_leaf_27_clk _01729_ net642 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[64\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17249_ net488 _00692_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08953_ addroundkey_data_o\[31\] mix1.data_o\[31\] _04778_ vssd1 vssd1 vccd1 vccd1
+ _04977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ _04713_ _04906_ _04907_ _04716_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09505_ net232 vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_211_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09436_ _05385_ vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09367_ fifo_bank_register.bank\[9\]\[32\] _05338_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08318_ addroundkey_data_o\[3\] fifo_bank_register.data_out\[3\] _04468_ vssd1 vssd1
+ vccd1 vccd1 _04472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09298_ fifo_bank_register.bank\[9\]\[10\] _05290_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05292_ sky130_fd_sc_hd__mux2_1
XANTENNA_50 _06401_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_61 addroundkey_data_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_72 addroundkey_data_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ net88 net87 net90 net89 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__or4_1
XANTENNA_83 addroundkey_data_o\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_94 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ _05491_ fifo_bank_register.bank\[8\]\[105\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10211_ sub1.data_o\[45\] _06024_ _05991_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ _05422_ fifo_bank_register.bank\[8\]\[72\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10142_ mix1.data_o\[38\] _05952_ _05916_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__o21a_1
XTAP_5800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10073_ _05567_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__clkbuf_8
X_14950_ _03221_ _03224_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__nor2_8
XTAP_5844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ _02298_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__clkbuf_1
XTAP_5888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14881_ addroundkey_data_o\[71\] _03061_ _03065_ addroundkey_data_o\[39\] vssd1 vssd1
+ vccd1 vccd1 _03157_ sky130_fd_sc_hd__a22o_1
XTAP_5899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13832_ fifo_bank_register.bank\[9\]\[30\] _02226_ _02231_ _02234_ _02237_ vssd1
+ vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a2111o_1
X_16620_ net515 _00068_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16551_ _05103_ _04946_ _05560_ _04361_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a31o_1
XFILLER_0_168_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ fifo_bank_register.bank\[7\]\[23\] _02128_ _02139_ fifo_bank_register.bank\[2\]\[23\]
+ _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a221o_1
XFILLER_0_202_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10975_ _06712_ _06713_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15502_ _03652_ _04777_ _05548_ _03665_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__a31o_1
X_12714_ fifo_bank_register.bank\[2\]\[22\] _05317_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07655_ sky130_fd_sc_hd__mux2_1
X_16482_ _04324_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__clkbuf_1
X_13694_ fifo_bank_register.bank\[5\]\[17\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18221_ clknet_leaf_36_clk _01652_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[51\]
+ sky130_fd_sc_hd__dfrtp_1
X_15433_ _03603_ _04949_ _05236_ _03622_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__a31o_1
X_12645_ _07617_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15364_ _04368_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__buf_4
X_18152_ clknet_leaf_81_clk _01583_ net586 vssd1 vssd1 vccd1 vccd1 ks1.col\[6\] sky130_fd_sc_hd__dfrtp_2
X_12576_ _07581_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14315_ _02667_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__clkbuf_1
X_17103_ net478 _00546_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18083_ net568 _01526_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[85\]
+ sky130_fd_sc_hd__dfxtp_1
X_11527_ _07027_ vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__clkbuf_1
X_15295_ _03145_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17034_ net521 _00477_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14246_ fifo_bank_register.bank\[0\]\[76\] _02605_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ _06935_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ _06171_ _06202_ _06203_ _06175_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14177_ fifo_bank_register.bank\[7\]\[69\] _02542_ _02470_ fifo_bank_register.bank\[2\]\[69\]
+ _02543_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a221o_1
X_11389_ fifo_bank_register.bank\[7\]\[37\] _05348_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ fifo_bank_register.bank\[1\]\[90\] _05459_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07873_ sky130_fd_sc_hd__mux2_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ net549 _01379_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
X_13059_ _07836_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17867_ net421 _01310_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16818_ clknet_leaf_4_clk _00262_ net591 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[109\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17798_ net509 _01241_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16749_ clknet_leaf_68_clk _00193_ net608 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[40\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09221_ sub1.data_o\[117\] _05197_ _05229_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18419_ clknet_leaf_12_clk _01849_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[104\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_185_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09152_ _05159_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_56_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_185_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09083_ _05085_ sbox1.ah\[2\] vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput70 data_i[47] vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_4
Xinput81 data_i[57] vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_2
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput92 data_i[67] vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09985_ _05757_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__buf_2
XTAP_5107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08936_ ks1.key_reg\[5\] _04745_ _04746_ net213 vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__o31a_1
XFILLER_0_200_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08867_ _04682_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__clkbuf_8
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08798_ mix1.data_o\[43\] _04698_ _04693_ _04821_ vssd1 vssd1 vccd1 vccd1 _04822_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10760_ net256 ks1.key_reg\[99\] _06402_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09419_ fifo_bank_register.bank\[9\]\[49\] _05373_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10691_ _06416_ _06455_ _06456_ _06420_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12430_ _07504_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12361_ _07467_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14100_ _02148_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_200_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _06914_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__clkbuf_1
X_15080_ _03348_ _03351_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__nor2_4
XFILLER_0_133_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12292_ _07364_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__buf_4
XFILLER_0_105_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14031_ fifo_bank_register.bank\[9\]\[52\] _02388_ _02412_ _02413_ _02414_ vssd1
+ vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__a2111o_1
X_11243_ _05474_ fifo_bank_register.bank\[8\]\[97\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06877_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11174_ _05405_ fifo_bank_register.bank\[8\]\[64\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10125_ net59 mix1.data_o\[37\] _05934_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__mux2_1
XTAP_5630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15982_ net223 ks1.key_reg\[69\] _03906_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__mux2_2
XTAP_5641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17721_ net430 _01164_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
X_14933_ _04376_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__buf_4
X_10056_ mix1.data_o\[31\] _05876_ _05821_ _05822_ sub1.data_o\[31\] vssd1 vssd1 vccd1
+ vccd1 _05884_ sky130_fd_sc_hd__a32o_1
XTAP_5674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17652_ net391 _01095_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14864_ _03124_ _03139_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16603_ net393 _00051_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_13815_ fifo_bank_register.bank\[1\]\[29\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__a22o_1
X_14795_ sub1.data_o\[112\] _03057_ _03070_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_159_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17583_ net464 _01026_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16534_ _04351_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__clkbuf_1
X_13746_ fifo_bank_register.bank\[5\]\[21\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[21\]
+ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__a22o_1
X_10958_ _06698_ vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13677_ _02098_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__clkbuf_1
X_16465_ net840 _04314_ _03957_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__mux2_1
X_10889_ net144 ks1.key_reg\[112\] _04639_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18204_ clknet_leaf_18_clk _01635_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15416_ _03581_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__clkbuf_4
X_12628_ fifo_bank_register.bank\[3\]\[110\] _05501_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16396_ ks1.key_reg\[94\] _04276_ _04264_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15347_ _03566_ vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18135_ clknet_leaf_53_clk sbox1.intermediate_to_invert_var\[1\] net656 vssd1 vssd1
+ vccd1 vccd1 sbox1.inversion_to_invert_var\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12559_ _07572_ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15278_ _03526_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__clkbuf_1
Xhold106 mix1.data_reg\[117\] vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__dlygate4sd3_1
X_18066_ net509 _01509_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold117 mix1.data_reg\[109\] vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold128 mix1.data_reg\[58\] vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14229_ fifo_bank_register.bank\[9\]\[74\] _02550_ _02588_ _02589_ _02590_ vssd1
+ vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__a2111o_1
Xhold139 ks1.key_reg\[55\] vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ net573 _00460_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout608 net612 vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_4
Xfanout619 net626 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09770_ _05628_ vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__clkbuf_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _04729_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ net549 _01362_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08652_ _04670_ _04671_ _04672_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__a22o_1
XFILLER_0_221_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08583_ _04611_ net258 vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__and2_1
XFILLER_0_194_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09204_ _05212_ _05213_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__xor2_2
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ sbox1.alph\[0\] _05142_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__nand2_2
XFILLER_0_45_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09066_ _05076_ _05080_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ _05712_ _05804_ _05805_ _05716_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__a22o_1
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _04701_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__clkbuf_4
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ sub1.data_o\[15\] _05742_ _05701_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__mux2_1
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _07240_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__clkbuf_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11861_ fifo_bank_register.bank\[5\]\[4\] _05278_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07204_ sky130_fd_sc_hd__mux2_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _08164_ fifo_bank_register.data_out\[6\] _08064_ vssd1 vssd1 vccd1 vccd1
+ _08165_ sky130_fd_sc_hd__mux2_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10812_ _06416_ _06565_ _06566_ _06420_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14580_ _02903_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__clkbuf_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11792_ _07078_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__buf_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ fifo_bank_register.bank\[7\]\[0\] _08078_ _08093_ fifo_bank_register.bank\[2\]\[0\]
+ _08101_ vssd1 vssd1 vccd1 vccd1 _08102_ sky130_fd_sc_hd__a221o_1
X_10743_ _06491_ _06502_ _06503_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ net160 ks1.key_reg\[127\] _04742_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__mux2_2
X_13462_ _08048_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__clkbuf_1
X_10674_ mix1.data_o\[91\] _06296_ _06320_ _06321_ sub1.data_o\[91\] vssd1 vssd1 vccd1
+ vccd1 _06442_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15201_ _03395_ _03463_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__xnor2_4
X_12413_ _07495_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16181_ net245 ks1.key_reg\[89\] _03918_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__mux2_2
XFILLER_0_153_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13393_ _08012_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15132_ _03180_ _03400_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__xor2_2
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12344_ _07458_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15063_ addroundkey_data_o\[124\] _03143_ _03334_ vssd1 vssd1 vccd1 vccd1 _03335_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12275_ _07422_ vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14014_ fifo_bank_register.bank\[9\]\[50\] _02388_ _02393_ _02396_ _02399_ vssd1
+ vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_120_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11226_ _05457_ fifo_bank_register.bank\[8\]\[89\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11157_ _05388_ fifo_bank_register.bank\[8\]\[56\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10108_ _05930_ _05931_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_218_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11088_ _05319_ fifo_bank_register.bank\[8\]\[23\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06796_ sky130_fd_sc_hd__mux2_1
X_15965_ _03918_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__buf_4
XTAP_5471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17704_ net446 _01147_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10039_ _05829_ _05867_ _05868_ _05833_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a22o_1
X_14916_ sub1.data_o\[110\] _03055_ _03190_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_175_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15896_ _03883_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__clkbuf_1
XTAP_4770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17635_ net499 _01078_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_14847_ addroundkey_data_o\[118\] _03077_ _03122_ vssd1 vssd1 vccd1 vccd1 _03123_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_81_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17566_ net540 _01009_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14778_ mix1.state\[1\] _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__nor2_4
XFILLER_0_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16517_ _04342_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13729_ fifo_bank_register.bank\[7\]\[20\] _02128_ _02139_ fifo_bank_register.bank\[2\]\[20\]
+ _02144_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17497_ net502 _00940_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16448_ _04304_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_186_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16379_ net822 _04119_ _04264_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18118_ net471 _01561_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[120\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18049_ net574 _01492_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout405 net413 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
XFILLER_0_226_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout416 net419 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__buf_2
XFILLER_0_201_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09822_ sub1.data_o\[7\] _05673_ _05610_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__mux2_1
Xfanout427 net444 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout438 net443 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_225_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout449 net461 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09753_ _04618_ _04629_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__or2_1
XFILLER_0_193_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08704_ _04722_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09684_ sub1.data_o\[121\] _05554_ _04891_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08635_ addroundkey_data_o\[124\] mix1.data_o\[124\] _04658_ vssd1 vssd1 vccd1 vccd1
+ _04659_ sky130_fd_sc_hd__mux2_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ addroundkey_data_o\[121\] fifo_bank_register.data_out\[121\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08497_ addroundkey_data_o\[88\] fifo_bank_register.data_out\[88\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__mux2_2
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09118_ _05105_ sbox1.inversion_to_invert_var\[0\] vssd1 vssd1 vccd1 vccd1 _05129_
+ sky130_fd_sc_hd__and2b_1
X_10390_ net87 mix1.data_o\[62\] _06158_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ _05058_ _05067_ vssd1 vssd1 vccd1 vccd1 sbox1.next_alph\[3\] sky130_fd_sc_hd__xor2_1
XFILLER_0_102_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12060_ _07308_ vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11011_ sub1.data_o\[125\] _06744_ _05609_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _03805_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__clkbuf_1
X_12962_ _07785_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__clkbuf_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _07231_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__clkbuf_1
X_14701_ _03009_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_310 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15681_ _03769_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__clkbuf_1
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _07748_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_321 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_332 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17420_ net519 _00863_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_343 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ fifo_bank_register.bank\[6\]\[125\] _05532_ _07055_ vssd1 vssd1 vccd1 vccd1
+ _07194_ sky130_fd_sc_hd__mux2_1
X_14632_ fifo_bank_register.bank\[6\]\[119\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[119\]
+ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_354 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17351_ net490 _00794_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _02888_ fifo_bank_register.data_out\[110\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11775_ _07158_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__clkbuf_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _04225_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__clkbuf_1
X_13514_ fifo_bank_register.write_ptr\[3\] _08085_ _05266_ vssd1 vssd1 vccd1 vccd1
+ _08086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10726_ _06488_ vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17282_ net512 _00725_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_14494_ fifo_bank_register.bank\[9\]\[103\] _02793_ _02824_ _02825_ _02826_ vssd1
+ vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ _05506_ fifo_bank_register.bank\[0\]\[112\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08040_ sky130_fd_sc_hd__mux2_1
X_16233_ _04177_ _04178_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__xor2_2
X_10657_ mix1.data_o\[89\] _06296_ _06320_ _06321_ sub1.data_o\[89\] vssd1 vssd1 vccd1
+ vccd1 _06427_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16164_ ks1.col\[24\] _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13376_ _08003_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__clkbuf_1
X_10588_ _06126_ _06362_ _06363_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15115_ _03321_ _03384_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_140_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12327_ _07449_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16095_ net237 ks1.key_reg\[81\] _03906_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__mux2_2
XFILLER_0_80_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15046_ addroundkey_data_o\[11\] _03208_ _03086_ _03318_ vssd1 vssd1 vccd1 vccd1
+ _03319_ sky130_fd_sc_hd__a211o_1
XFILLER_0_220_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12258_ _07413_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11209_ _06859_ vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__clkbuf_1
X_12189_ _07377_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16997_ net423 _00440_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ _03920_ _03921_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__xor2_2
XFILLER_0_190_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15879_ sub1.data_o\[94\] _05235_ _04888_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ addroundkey_data_o\[51\] fifo_bank_register.data_out\[51\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17618_ net500 _01061_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18598_ clknet_leaf_68_clk _02027_ net608 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[125\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08351_ _04489_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17549_ net517 _00992_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08282_ net161 net162 net152 net141 vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__and4b_1
XFILLER_0_184_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09805_ net84 mix1.data_o\[5\] _05604_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09736_ _05588_ round\[2\] round\[3\] vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__or3b_1
XFILLER_0_213_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09667_ addroundkey_round\[0\] addroundkey_round\[1\] addroundkey_round\[2\] vssd1
+ vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_213_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08618_ addroundkey_start_i _04641_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__nand2_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ net138 vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__buf_2
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _04593_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _07044_ vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10511_ net102 mix1.data_o\[76\] _06237_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11491_ _07008_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13230_ _05290_ fifo_bank_register.bank\[0\]\[10\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07927_ sky130_fd_sc_hd__mux2_1
X_10442_ _06171_ _06231_ _06232_ _06175_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13161_ fifo_bank_register.bank\[1\]\[106\] _05493_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07890_ sky130_fd_sc_hd__mux2_1
X_10373_ net85 mix1.data_o\[60\] _06158_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12112_ _07335_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13092_ fifo_bank_register.bank\[1\]\[73\] _05424_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12043_ fifo_bank_register.bank\[5\]\[90\] _05459_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07300_ sky130_fd_sc_hd__mux2_1
X_16920_ net560 _00363_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
X_16851_ net517 _00294_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15802_ mix1.data_o\[101\] net784 _03830_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16782_ clknet_leaf_73_clk _00226_ net593 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[73\]
+ sky130_fd_sc_hd__dfrtp_4
X_13994_ fifo_bank_register.bank\[5\]\[49\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[49\]
+ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18521_ clknet_leaf_66_clk _01950_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
X_15733_ _03796_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__clkbuf_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _07776_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__clkbuf_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ clknet_leaf_70_clk _01882_ net608 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[92\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15664_ _03760_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__clkbuf_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_140 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _07739_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_151 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_162 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17403_ net567 _00846_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_173 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ fifo_bank_register.bank\[6\]\[117\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[117\]
+ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__a22o_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_213_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18383_ clknet_leaf_25_clk _01813_ net648 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[68\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_185_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_184 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11827_ _07185_ vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__clkbuf_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _03723_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__clkbuf_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_195 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ net412 _00777_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
X_14546_ _02872_ fifo_bank_register.data_out\[109\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02873_ sky130_fd_sc_hd__mux2_1
X_11758_ _07149_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10709_ net252 ks1.key_reg\[95\] _06324_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17265_ net392 _00708_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
X_14477_ fifo_bank_register.bank\[1\]\[101\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[101\]
+ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__a22o_1
X_11689_ _07113_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16216_ ks1.col\[28\] _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__xor2_4
XFILLER_0_181_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13428_ _05489_ fifo_bank_register.bank\[0\]\[104\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17196_ net465 _00639_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13359_ _05420_ fifo_bank_register.bank\[0\]\[71\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _07995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16147_ net151 ks1.key_reg\[119\] _03976_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16078_ _05244_ _04037_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__xor2_2
XFILLER_0_228_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15029_ addroundkey_data_o\[2\] _04375_ _04900_ _03301_ vssd1 vssd1 vccd1 vccd1 _03302_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput2 data_i[100] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__buf_2
XFILLER_0_194_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09521_ net238 vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_196_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09452_ net214 vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ addroundkey_data_o\[43\] fifo_bank_register.data_out\[43\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__mux2_4
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09383_ _05349_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ addroundkey_data_o\[10\] fifo_bank_register.data_out\[10\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__mux2_2
XFILLER_0_164_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08265_ net160 net40 net1 net159 vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__or4b_1
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput350 net350 vssd1 vssd1 vccd1 vccd1 data_o[66] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput361 net361 vssd1 vssd1 vccd1 vccd1 data_o[76] sky130_fd_sc_hd__clkbuf_4
Xoutput372 net372 vssd1 vssd1 vccd1 vccd1 data_o[86] sky130_fd_sc_hd__clkbuf_4
Xoutput383 net383 vssd1 vssd1 vccd1 vccd1 data_o[96] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09719_ _05198_ net258 _05568_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__a21oi_1
X_10991_ _06726_ _06727_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__xor2_1
XFILLER_0_214_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _07651_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _07625_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ fifo_bank_register.bank\[7\]\[93\] _02704_ _02713_ fifo_bank_register.bank\[2\]\[93\]
+ _02742_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__a221o_1
X_11612_ _07072_ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ sub1.data_o\[37\] sub1.data_o\[101\] _05202_ vssd1 vssd1 vccd1 vccd1 _03587_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12592_ fifo_bank_register.bank\[3\]\[93\] _05466_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14331_ _02681_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__clkbuf_1
X_11543_ fifo_bank_register.bank\[7\]\[110\] _05501_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14262_ fifo_bank_register.bank\[9\]\[78\] _02550_ _02617_ _02618_ _02619_ vssd1
+ vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a2111o_1
X_17050_ net536 _00493_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11474_ _06999_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13213_ _05274_ fifo_bank_register.bank\[0\]\[2\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07918_ sky130_fd_sc_hd__mux2_1
X_16001_ ks1.col\[7\] _03968_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__xor2_4
X_10425_ mix1.data_o\[66\] _06217_ _06162_ _06163_ sub1.data_o\[66\] vssd1 vssd1 vccd1
+ vccd1 _06218_ sky130_fd_sc_hd__a32o_1
X_14193_ _02151_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13144_ fifo_bank_register.bank\[1\]\[98\] _05476_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07881_ sky130_fd_sc_hd__mux2_1
X_10356_ addroundkey_data_o\[58\] _06156_ _06064_ vssd1 vssd1 vccd1 vccd1 _06157_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17952_ net406 _01395_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
X_13075_ fifo_bank_register.bank\[1\]\[65\] _05407_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07845_ sky130_fd_sc_hd__mux2_1
X_10287_ mix1.data_o\[52\] _05952_ _06093_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16903_ net518 _00346_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12026_ fifo_bank_register.bank\[5\]\[82\] _05443_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17883_ net482 _01326_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16834_ clknet_leaf_47_clk _00278_ net651 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[125\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16765_ clknet_leaf_48_clk _00209_ net611 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[56\]
+ sky130_fd_sc_hd__dfrtp_4
X_13977_ fifo_bank_register.bank\[7\]\[47\] _02299_ _02308_ fifo_bank_register.bank\[2\]\[47\]
+ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18504_ clknet_leaf_61_clk _01933_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_15716_ mix1.data_o\[60\] net742 _03786_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__mux2_1
X_12928_ _07766_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__clkbuf_1
X_16696_ clknet_leaf_72_clk _00143_ net594 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[123\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18435_ clknet_leaf_23_clk _01865_ net645 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[120\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_185_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15647_ _03751_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ fifo_bank_register.bank\[2\]\[91\] _05462_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07731_ sky130_fd_sc_hd__mux2_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18366_ clknet_leaf_36_clk _01796_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[51\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_150_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15578_ _03700_ _03709_ _05196_ _03714_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17317_ net400 _00760_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
X_14529_ _02856_ fifo_bank_register.data_out\[107\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18297_ clknet_leaf_46_clk _01728_ net652 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17248_ net508 _00691_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17179_ net567 _00622_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08952_ addroundkey_data_o\[55\] mix1.data_o\[55\] _04656_ vssd1 vssd1 vccd1 vccd1
+ _04976_ sky130_fd_sc_hd__mux2_1
X_08883_ addroundkey_data_o\[88\] mix1.data_o\[88\] _04702_ vssd1 vssd1 vccd1 vccd1
+ _04907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09504_ _05431_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09435_ fifo_bank_register.bank\[9\]\[54\] _05384_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05385_ sky130_fd_sc_hd__mux2_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09366_ net183 vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08317_ _04471_ vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_40 _05553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09297_ _05269_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__buf_4
XFILLER_0_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_51 addroundkey_data_o\[112\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_62 addroundkey_data_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08248_ net79 net78 net81 net80 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__or4_1
XANTENNA_73 addroundkey_data_o\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 addroundkey_data_o\[73\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_95 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10210_ net68 mix1.data_o\[45\] _05989_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ _06849_ vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10141_ _05949_ _05960_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10072_ _05898_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__clkbuf_1
XTAP_5834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13900_ _02297_ fifo_bank_register.data_out\[38\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02298_ sky130_fd_sc_hd__mux2_1
XTAP_5867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14880_ sub1.data_o\[103\] _03054_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__a21oi_2
XTAP_5889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13831_ fifo_bank_register.bank\[1\]\[30\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16550_ sub1.data_o\[114\] _05197_ _04360_ _03594_ vssd1 vssd1 vccd1 vccd1 _04361_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13762_ fifo_bank_register.bank\[5\]\[23\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[23\]
+ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__a22o_1
X_10974_ net153 ks1.key_reg\[120\] _06579_ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15501_ sub1.data_o\[48\] _03663_ _03664_ _03611_ vssd1 vssd1 vccd1 vccd1 _03665_
+ sky130_fd_sc_hd__a22o_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12713_ _07654_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__clkbuf_1
X_16481_ net722 _03283_ _04321_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13693_ _02112_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__clkbuf_1
X_18220_ clknet_leaf_19_clk _01651_ net640 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[50\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15432_ sub1.data_o\[22\] _03606_ _03621_ _03611_ vssd1 vssd1 vccd1 vccd1 _03622_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12644_ fifo_bank_register.bank\[3\]\[118\] _05518_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18151_ clknet_leaf_81_clk _01582_ net578 vssd1 vssd1 vccd1 vccd1 ks1.col\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15363_ sub1.data_o\[32\] sub1.data_o\[96\] _03574_ vssd1 vssd1 vccd1 vccd1 _03575_
+ sky130_fd_sc_hd__mux2_1
X_12575_ fifo_bank_register.bank\[3\]\[85\] _05449_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17102_ net478 _00545_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_14314_ _02666_ fifo_bank_register.data_out\[83\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18082_ net537 _01525_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[84\]
+ sky130_fd_sc_hd__dfxtp_2
X_11526_ fifo_bank_register.bank\[7\]\[102\] _05485_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07027_ sky130_fd_sc_hd__mux2_1
X_15294_ _03538_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17033_ net515 _00476_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11457_ _06990_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__clkbuf_1
X_14245_ fifo_bank_register.bank\[9\]\[76\] _02550_ _02602_ _02603_ _02604_ vssd1
+ vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_123_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10408_ mix1.data_o\[64\] _06138_ _06162_ _06163_ sub1.data_o\[64\] vssd1 vssd1 vccd1
+ vccd1 _06203_ sky130_fd_sc_hd__a32o_1
XFILLER_0_1_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14176_ fifo_bank_register.bank\[5\]\[69\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[69\]
+ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11388_ _06954_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10339_ _06140_ _06141_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13127_ _07794_ vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__buf_4
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ net554 _01378_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
X_13058_ fifo_bank_register.bank\[1\]\[57\] _05390_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12009_ fifo_bank_register.bank\[5\]\[74\] _05426_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07282_ sky130_fd_sc_hd__mux2_1
X_17866_ net420 _01309_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16817_ clknet_leaf_82_clk _00261_ net585 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[108\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17797_ net524 _01240_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16748_ clknet_leaf_65_clk _00192_ net604 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16679_ net435 _00127_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09220_ sub1.data_o\[21\] _05200_ _05203_ sub1.data_o\[85\] vssd1 vssd1 vccd1 vccd1
+ _05229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18418_ clknet_leaf_13_clk _01848_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[103\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_173_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ _05160_ _05161_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__xnor2_2
X_18349_ clknet_leaf_15_clk _01779_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09082_ _05016_ _05058_ _05094_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput60 data_i[38] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_2
Xinput71 data_i[48] vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_2
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput82 data_i[58] vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_4
Xinput93 data_i[68] vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09984_ sub1.data_o\[23\] _05818_ _05819_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08935_ ks1.key_reg\[13\] _04726_ _04958_ net162 vssd1 vssd1 vccd1 vccd1 _04959_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_228_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08866_ addroundkey_data_o\[112\] mix1.data_o\[112\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ addroundkey_data_o\[43\] _04663_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__or2_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09418_ net201 vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10690_ mix1.data_o\[93\] _06296_ _06320_ _06321_ sub1.data_o\[93\] vssd1 vssd1 vccd1
+ vccd1 _06456_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09349_ _05326_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12360_ _05506_ fifo_bank_register.bank\[4\]\[112\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ fifo_bank_register.bank\[7\]\[0\] _05248_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12291_ _07430_ vssd1 vssd1 vccd1 vccd1 _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14030_ fifo_bank_register.bank\[1\]\[52\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[52\]
+ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__a22o_1
X_11242_ _06876_ vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11173_ _06840_ vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10124_ _05946_ vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__clkbuf_1
XTAP_5620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15981_ ks1.col\[5\] _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__xor2_4
XTAP_5631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17720_ net408 _01163_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10055_ sub1.data_o\[31\] _05882_ _05819_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__mux2_1
X_14932_ _03203_ _03206_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__nor2_8
XTAP_5664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ net405 _01094_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _03131_ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__xnor2_4
XTAP_4974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16602_ net405 _00050_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13814_ fifo_bank_register.bank\[6\]\[29\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__a22o_1
X_17582_ net462 _01025_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14794_ sub1.data_o\[16\] _04378_ _03059_ _03069_ vssd1 vssd1 vccd1 vccd1 _03070_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_159_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16533_ net774 _03525_ _04343_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__mux2_1
X_13745_ _02160_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10957_ addroundkey_data_o\[118\] _06697_ _06612_ vssd1 vssd1 vccd1 vccd1 _06698_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16464_ _04175_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13676_ _02097_ fifo_bank_register.data_out\[14\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _02098_ sky130_fd_sc_hd__mux2_1
X_10888_ _05623_ _06629_ _06634_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_167_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18203_ clknet_leaf_15_clk _01634_ net637 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15415_ sub1.data_o\[113\] sub1.data_o\[49\] _03609_ vssd1 vssd1 vccd1 vccd1 _03610_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12627_ _07508_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16395_ _04187_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18134_ clknet_leaf_53_clk sbox1.intermediate_to_invert_var\[0\] net656 vssd1 vssd1
+ vccd1 vccd1 sbox1.inversion_to_invert_var\[0\] sky130_fd_sc_hd__dfrtp_2
X_15346_ net756 _03514_ _03560_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12558_ fifo_bank_register.bank\[3\]\[77\] _05432_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18065_ net508 _01508_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_11509_ fifo_bank_register.bank\[7\]\[94\] _05468_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07018_ sky130_fd_sc_hd__mux2_1
X_15277_ net736 _03525_ _03498_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold107 mix1.data_reg\[76\] vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ fifo_bank_register.bank\[3\]\[44\] _05363_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold118 mix1.data_reg\[49\] vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17016_ net558 _00459_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold129 ks1.key_reg\[99\] vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14228_ fifo_bank_register.bank\[1\]\[74\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[74\]
+ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14159_ fifo_bank_register.bank\[7\]\[67\] _02461_ _02470_ fifo_bank_register.bank\[2\]\[67\]
+ _02527_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a221o_1
Xfanout609 net612 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__buf_2
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08720_ ks1.key_reg\[20\] _04742_ _04743_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__a21oi_1
X_17918_ net574 _01361_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08651_ _04674_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__clkbuf_4
X_17849_ net469 _01292_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08582_ _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09203_ _05170_ _05192_ vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_130_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09134_ _05140_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_228_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09065_ sbox1.ah\[3\] sbox1.ah\[0\] _05067_ _05074_ _05079_ vssd1 vssd1 vccd1 vccd1
+ _05080_ sky130_fd_sc_hd__a41o_1
XFILLER_0_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09967_ mix1.data_o\[21\] _05797_ _05703_ _05704_ sub1.data_o\[21\] vssd1 vssd1 vccd1
+ vccd1 _05805_ sky130_fd_sc_hd__a32o_1
XFILLER_0_228_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08918_ _04940_ _04941_ _04900_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__mux2_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ net35 mix1.data_o\[15\] _05699_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__mux2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _04833_ _04872_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__xnor2_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _07203_ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10811_ mix1.data_o\[104\] _06463_ _06320_ _06321_ sub1.data_o\[104\] vssd1 vssd1
+ vccd1 vccd1 _06566_ sky130_fd_sc_hd__a32o_1
X_11791_ _07166_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__clkbuf_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13530_ fifo_bank_register.bank\[5\]\[0\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08101_ sky130_fd_sc_hd__a22o_1
X_10742_ _06395_ _06342_ sub1.data_o\[98\] _06384_ vssd1 vssd1 vccd1 vccd1 _06503_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10673_ sub1.data_o\[91\] _06440_ _06318_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__mux2_1
X_13461_ _05522_ fifo_bank_register.bank\[0\]\[120\] _07914_ vssd1 vssd1 vccd1 vccd1
+ _08048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ _03420_ _03461_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__o21a_1
XFILLER_0_180_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12412_ fifo_bank_register.bank\[3\]\[8\] _05286_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16180_ _04128_ _04129_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13392_ _05453_ fifo_bank_register.bank\[0\]\[87\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15131_ _03245_ _03399_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12343_ _05489_ fifo_bank_register.bank\[4\]\[104\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15062_ addroundkey_data_o\[28\] _04379_ _05607_ _03333_ vssd1 vssd1 vccd1 vccd1
+ _03334_ sky130_fd_sc_hd__a211o_1
X_12274_ _05420_ fifo_bank_register.bank\[4\]\[71\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11225_ _06867_ vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__clkbuf_1
X_14013_ fifo_bank_register.bank\[1\]\[50\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[50\]
+ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11156_ _06831_ vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__clkbuf_1
XTAP_6140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10107_ net186 ks1.key_reg\[35\] _05920_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__mux2_2
XTAP_5450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11087_ _06795_ vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__clkbuf_1
X_15964_ _03934_ _03935_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__xor2_2
XTAP_5461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput250 key_i[93] vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17703_ net448 _01146_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10038_ mix1.data_o\[29\] _05797_ _05821_ _05822_ sub1.data_o\[29\] vssd1 vssd1 vccd1
+ vccd1 _05868_ sky130_fd_sc_hd__a32o_1
X_14915_ sub1.data_o\[14\] _03100_ _03058_ _03189_ vssd1 vssd1 vccd1 vccd1 _03190_
+ sky130_fd_sc_hd__a211o_1
XTAP_5494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_216_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15895_ sub1.data_o\[99\] _03882_ _03876_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__mux2_1
XTAP_4760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17634_ net486 _01077_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14846_ addroundkey_data_o\[22\] _04375_ _04900_ _03121_ vssd1 vssd1 vccd1 vccd1
+ _03122_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17565_ net538 _01008_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
X_14777_ state _04622_ _03052_ mix1.state\[0\] vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a211o_1
XFILLER_0_105_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11989_ _07271_ vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16516_ net696 _03497_ _04332_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13728_ fifo_bank_register.bank\[5\]\[20\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17496_ net497 _00939_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16447_ net835 _04092_ _04295_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__mux2_1
X_13659_ fifo_bank_register.bank\[0\]\[12\] _02082_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16378_ _04265_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18117_ net431 _01560_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15329_ net741 _03487_ _03549_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18048_ net557 _01491_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout406 net413 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_1
X_09821_ net106 mix1.data_o\[7\] _05604_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__mux2_1
Xfanout417 net419 vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_2
XFILLER_0_226_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout428 net431 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__buf_2
Xfanout439 net443 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_2
XFILLER_0_201_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09752_ sub1.data_o\[0\] _05605_ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08703_ ks1.ready_o _04636_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_213_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09683_ _05553_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _04657_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _04601_ vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08496_ _04565_ vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__buf_1
XFILLER_0_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09117_ sbox1.alph\[1\] _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09048_ _04877_ _05065_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11010_ net29 mix1.data_o\[125\] _05603_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12961_ fifo_bank_register.bank\[1\]\[11\] _05293_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07785_ sky130_fd_sc_hd__mux2_1
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _03008_ fifo_bank_register.data_out\[127\] _08068_ vssd1 vssd1 vccd1 vccd1
+ _03009_ sky130_fd_sc_hd__mux2_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ fifo_bank_register.bank\[5\]\[28\] _05329_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07231_ sky130_fd_sc_hd__mux2_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ mix1.data_o\[43\] net723 _03764_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__mux2_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ fifo_bank_register.bank\[2\]\[107\] _05495_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07748_ sky130_fd_sc_hd__mux2_1
XANTENNA_311 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_322 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_333 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ fifo_bank_register.bank\[7\]\[119\] _08077_ _02875_ fifo_bank_register.bank\[2\]\[119\]
+ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__a221o_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _07193_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__clkbuf_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_344 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ net473 _00793_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ fifo_bank_register.bank\[0\]\[110\] _02886_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02888_ sky130_fd_sc_hd__mux2_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ fifo_bank_register.bank\[6\]\[91\] _05462_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07158_ sky130_fd_sc_hd__mux2_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ net816 _04072_ _04222_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__mux2_1
X_13513_ _05256_ vssd1 vssd1 vccd1 vccd1 _08085_ sky130_fd_sc_hd__inv_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ addroundkey_data_o\[96\] _06487_ _06431_ vssd1 vssd1 vccd1 vccd1 _06488_
+ sky130_fd_sc_hd__mux2_1
X_17281_ net570 _00724_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14493_ fifo_bank_register.bank\[1\]\[103\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[103\]
+ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16232_ net215 ks1.key_reg\[61\] _03982_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__mux2_1
X_13444_ _08039_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10656_ sub1.data_o\[89\] _06425_ _06318_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16163_ _04111_ _04112_ _04113_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__and3_1
X_10587_ _06090_ _06342_ sub1.data_o\[83\] _06079_ vssd1 vssd1 vccd1 vccd1 _06363_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13375_ _05436_ fifo_bank_register.bank\[0\]\[79\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _08003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15114_ _03246_ _03297_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12326_ _05472_ fifo_bank_register.bank\[4\]\[96\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16094_ ks1.col\[17\] _04051_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__xor2_4
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ addroundkey_data_o\[75\] _03064_ _03084_ addroundkey_data_o\[43\] vssd1 vssd1
+ vccd1 vccd1 _03318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12257_ _05403_ fifo_bank_register.bank\[4\]\[63\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ _05438_ fifo_bank_register.bank\[8\]\[80\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06859_ sky130_fd_sc_hd__mux2_1
X_12188_ _05333_ fifo_bank_register.bank\[4\]\[30\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11139_ _06822_ vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__clkbuf_1
X_16996_ net424 _00439_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15947_ net184 ks1.key_reg\[33\] _03910_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__mux2_1
XTAP_5280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15878_ _03871_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14829_ addroundkey_data_o\[6\] _03100_ _05606_ _03104_ vssd1 vssd1 vccd1 vccd1 _03105_
+ sky130_fd_sc_hd__a211o_1
X_17617_ net503 _01060_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_18597_ clknet_leaf_67_clk _02026_ net610 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[124\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08350_ addroundkey_data_o\[18\] fifo_bank_register.data_out\[18\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17548_ net517 _00991_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08281_ net130 net169 _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17479_ net492 _00922_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09804_ _05658_ vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09735_ round\[3\] _05590_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_158_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09666_ addroundkey_round\[0\] addroundkey_round\[1\] addroundkey_round\[2\] vssd1
+ vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08617_ round\[3\] _04614_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__or2_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09597_ _05494_ vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ addroundkey_data_o\[112\] fifo_bank_register.data_out\[112\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__mux2_4
XFILLER_0_33_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08479_ addroundkey_data_o\[79\] fifo_bank_register.data_out\[79\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10510_ _06293_ vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__clkbuf_1
X_11490_ fifo_bank_register.bank\[7\]\[85\] _05449_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10441_ mix1.data_o\[68\] _06217_ _06162_ _06163_ sub1.data_o\[68\] vssd1 vssd1 vccd1
+ vccd1 _06232_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10372_ _05615_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13160_ _07889_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12111_ fifo_bank_register.bank\[5\]\[123\] _05528_ _07198_ vssd1 vssd1 vccd1 vccd1
+ _07335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13091_ _07853_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12042_ _07221_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__buf_4
X_16850_ net504 _00293_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15801_ _03832_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__clkbuf_1
X_16781_ clknet_leaf_77_clk _00225_ net590 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[72\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_217_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13993_ _08181_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_176_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18520_ clknet_leaf_66_clk _01949_ net606 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_1
X_15732_ mix1.data_o\[68\] net839 _03786_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__mux2_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12944_ fifo_bank_register.bank\[1\]\[3\] _05276_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07776_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ clknet_leaf_73_clk _01881_ net593 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[91\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15663_ mix1.data_o\[35\] net735 _03753_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_130 mix1.data_o\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ fifo_bank_register.bank\[2\]\[99\] _05478_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07739_ sky130_fd_sc_hd__mux2_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_141 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_152 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17402_ net567 _00845_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14614_ fifo_bank_register.bank\[7\]\[117\] _02866_ _02875_ fifo_bank_register.bank\[2\]\[117\]
+ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__a221o_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ clknet_leaf_26_clk _01812_ net648 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[67\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_185_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_163 net96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ fifo_bank_register.bank\[6\]\[116\] _05514_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07185_ sky130_fd_sc_hd__mux2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15594_ mix1.data_o\[3\] _03324_ mix1.next_ready_o vssd1 vssd1 vccd1 vccd1 _03723_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_174 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_185 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_196 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ net412 _00776_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14545_ fifo_bank_register.bank\[0\]\[109\] _02871_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02872_ sky130_fd_sc_hd__mux2_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ fifo_bank_register.bank\[6\]\[83\] _05445_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07149_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10708_ _06416_ _06470_ _06471_ _06420_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__a22o_2
X_17264_ net390 _00707_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14476_ fifo_bank_register.bank\[6\]\[101\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[101\]
+ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__a22o_1
X_11688_ fifo_bank_register.bank\[6\]\[50\] _05375_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16215_ _04112_ _04113_ _04124_ _04151_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13427_ _08030_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__clkbuf_1
X_10639_ sub1.data_o\[87\] _06341_ _06409_ _06410_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06411_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17195_ net450 _00638_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16146_ _04098_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _07994_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12309_ _05455_ fifo_bank_register.bank\[4\]\[88\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16077_ net143 ks1.key_reg\[111\] _03905_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13289_ _05350_ fifo_bank_register.bank\[0\]\[38\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15028_ addroundkey_data_o\[66\] _03062_ _03091_ addroundkey_data_o\[34\] vssd1 vssd1
+ vccd1 vccd1 _03301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_220_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput3 data_i[101] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_4
X_16979_ net506 _00422_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09520_ _05442_ vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09451_ _05395_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08402_ _04516_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09382_ fifo_bank_register.bank\[9\]\[37\] _05348_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08333_ _04480_ vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08264_ net151 net154 net153 net150 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__or4b_1
XFILLER_0_7_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput340 net340 vssd1 vssd1 vccd1 vccd1 data_o[57] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput351 net351 vssd1 vssd1 vccd1 vccd1 data_o[67] sky130_fd_sc_hd__clkbuf_4
Xoutput362 net362 vssd1 vssd1 vccd1 vccd1 data_o[77] sky130_fd_sc_hd__clkbuf_4
Xoutput373 net373 vssd1 vssd1 vccd1 vccd1 data_o[87] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput384 net384 vssd1 vssd1 vccd1 vccd1 data_o[97] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09718_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_173_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10990_ net155 ks1.key_reg\[122\] _06579_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09649_ _05529_ vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__clkbuf_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ fifo_bank_register.bank\[3\]\[126\] _05534_ _07485_ vssd1 vssd1 vccd1 vccd1
+ _07625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ fifo_bank_register.bank\[6\]\[14\] _05299_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12591_ _07589_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14330_ _02680_ fifo_bank_register.data_out\[85\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _06935_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14261_ fifo_bank_register.bank\[1\]\[78\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[78\]
+ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11473_ fifo_bank_register.bank\[7\]\[77\] _05432_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _06999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16000_ net134 ks1.key_reg\[103\] _03902_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__mux2_2
XFILLER_0_208_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13212_ _07917_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10424_ _05585_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14192_ fifo_bank_register.bank\[6\]\[70\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[70\]
+ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ _07880_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__clkbuf_1
X_10355_ _06154_ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _05757_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__clkbuf_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _07844_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__clkbuf_1
X_17951_ net547 _01394_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16902_ net509 _00345_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
X_12025_ _07290_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__clkbuf_1
X_17882_ net513 _01325_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16833_ clknet_leaf_47_clk _00277_ net612 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[124\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_79_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16764_ clknet_leaf_39_clk _00208_ net668 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[55\]
+ sky130_fd_sc_hd__dfrtp_4
X_13976_ fifo_bank_register.bank\[5\]\[47\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[47\]
+ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a22o_1
XFILLER_0_219_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15715_ _03787_ vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18503_ clknet_leaf_59_clk _01932_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12927_ fifo_bank_register.bank\[2\]\[124\] _05530_ _07628_ vssd1 vssd1 vccd1 vccd1
+ _07766_ sky130_fd_sc_hd__mux2_1
X_16695_ clknet_leaf_5_clk _00142_ net592 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18434_ clknet_leaf_24_clk _01864_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[119\]
+ sky130_fd_sc_hd__dfrtp_2
X_15646_ mix1.data_o\[27\] _03525_ _03742_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12858_ _07730_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18365_ clknet_leaf_35_clk _01795_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[50\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_158_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11809_ fifo_bank_register.bank\[6\]\[108\] _05497_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15577_ sub1.data_o\[11\] _03660_ _03710_ sub1.data_o\[75\] vssd1 vssd1 vccd1 vccd1
+ _03714_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12789_ fifo_bank_register.bank\[2\]\[58\] _05392_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17316_ net448 _00759_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ _08063_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__buf_4
X_18296_ clknet_leaf_51_clk _01727_ net651 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[62\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17247_ net487 _00690_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_14459_ _02140_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17178_ net547 _00621_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16129_ net149 ks1.key_reg\[117\] _03902_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ _04661_ _04973_ _04974_ _04668_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08882_ addroundkey_data_o\[64\] mix1.data_o\[64\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ fifo_bank_register.bank\[9\]\[76\] _05430_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09434_ net207 vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09365_ _05337_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08316_ addroundkey_data_o\[2\] fifo_bank_register.data_out\[2\] _04468_ vssd1 vssd1
+ vccd1 vccd1 _04471_ sky130_fd_sc_hd__mux2_2
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09296_ net141 vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_41 _05553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_52 addroundkey_data_o\[112\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_63 addroundkey_data_o\[25\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ net83 net82 net86 net85 vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__or4_1
XFILLER_0_144_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_74 addroundkey_data_o\[50\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_85 addroundkey_data_o\[73\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_96 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10140_ _05913_ _05754_ sub1.data_o\[38\] _05902_ vssd1 vssd1 vccd1 vccd1 _05961_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10071_ addroundkey_data_o\[32\] _05897_ _05872_ vssd1 vssd1 vccd1 vccd1 _05898_
+ sky130_fd_sc_hd__mux2_1
XTAP_5824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13830_ _02153_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_215_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13761_ _02174_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__clkbuf_1
X_10973_ _06583_ _06710_ _06711_ _06587_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15500_ sub1.data_o\[16\] sub1.data_o\[80\] _03609_ vssd1 vssd1 vccd1 vccd1 _03664_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12712_ fifo_bank_register.bank\[2\]\[21\] _05315_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16480_ _04323_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__clkbuf_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13692_ _02111_ fifo_bank_register.data_out\[16\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _02112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15431_ sub1.data_o\[118\] sub1.data_o\[54\] _03609_ vssd1 vssd1 vccd1 vccd1 _03621_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12643_ _07616_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18150_ clknet_leaf_81_clk _01581_ net586 vssd1 vssd1 vccd1 vccd1 ks1.col\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ _05202_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__buf_4
XFILLER_0_136_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12574_ _07580_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17101_ net477 _00544_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14313_ fifo_bank_register.bank\[0\]\[83\] _02665_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18081_ net568 _01524_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[83\]
+ sky130_fd_sc_hd__dfxtp_1
X_11525_ _07026_ vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__clkbuf_1
X_15293_ net725 _03537_ _03144_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17032_ net526 _00475_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14244_ fifo_bank_register.bank\[1\]\[76\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[76\]
+ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11456_ fifo_bank_register.bank\[7\]\[69\] _05415_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10407_ sub1.data_o\[64\] _06201_ _06160_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14175_ _08181_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11387_ fifo_bank_register.bank\[7\]\[36\] _05346_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13126_ _07871_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ net209 ks1.key_reg\[56\] _05997_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__mux2_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ net554 _01377_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
X_13057_ _07835_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__clkbuf_1
X_10269_ net75 mix1.data_o\[51\] _05934_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__mux2_1
X_12008_ _07281_ vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17865_ net420 _01308_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16816_ clknet_leaf_82_clk _00260_ net585 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[107\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17796_ net511 _01239_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16747_ clknet_leaf_45_clk _00191_ net653 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[38\]
+ sky130_fd_sc_hd__dfrtp_4
X_13959_ _02350_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16678_ net456 _00126_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18417_ clknet_leaf_11_clk _01847_ net628 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[102\]
+ sky130_fd_sc_hd__dfrtp_2
X_15629_ _03741_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_185_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09150_ sbox1.ah_reg\[2\] _05134_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__nand2_1
X_18348_ clknet_leaf_16_clk _01778_ net637 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[33\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09081_ sbox1.ah\[3\] _05071_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__and2_1
X_18279_ clknet_leaf_5_clk _01710_ net592 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[45\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput50 data_i[29] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput61 data_i[39] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_4
Xinput72 data_i[49] vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__buf_2
XFILLER_0_163_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput83 data_i[59] vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput94 data_i[69] vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_4
XFILLER_0_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ _05609_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ ks1.key_reg\[13\] _04730_ _04732_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__or3_1
XTAP_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08865_ addroundkey_data_o\[80\] mix1.data_o\[80\] _04666_ vssd1 vssd1 vccd1 vccd1
+ _04889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08796_ _04818_ _04819_ _04702_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09417_ _05372_ vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09348_ fifo_bank_register.bank\[9\]\[26\] _05325_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09279_ fifo_bank_register.bank\[9\]\[4\] _05278_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ _06912_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12290_ _05436_ fifo_bank_register.bank\[4\]\[79\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ _05472_ fifo_bank_register.bank\[8\]\[96\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ _05403_ fifo_bank_register.bank\[8\]\[63\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ addroundkey_data_o\[36\] _05945_ _05872_ vssd1 vssd1 vccd1 vccd1 _05946_
+ sky130_fd_sc_hd__mux2_1
X_15980_ net132 ks1.key_reg\[101\] _03905_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__mux2_2
XTAP_5610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10054_ net53 mix1.data_o\[31\] _05817_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__mux2_1
X_14931_ addroundkey_data_o\[121\] _03078_ _03205_ vssd1 vssd1 vccd1 vccd1 _03206_
+ sky130_fd_sc_hd__a21oi_2
XTAP_5654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14862_ _03134_ _03137_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__nor2_8
X_17650_ net391 _01093_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16601_ net398 _00049_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_13813_ fifo_bank_register.bank\[7\]\[29\] _02218_ _02139_ fifo_bank_register.bank\[2\]\[29\]
+ _02219_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__a221o_1
XFILLER_0_188_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17581_ net464 _01024_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14793_ sub1.data_o\[80\] _03064_ _03068_ sub1.data_o\[48\] vssd1 vssd1 vccd1 vccd1
+ _03069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16532_ _04350_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13744_ _02159_ fifo_bank_register.data_out\[20\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02160_ sky130_fd_sc_hd__mux2_1
X_10956_ _06695_ _06696_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16463_ _04313_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13675_ fifo_bank_register.bank\[0\]\[14\] _02096_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02097_ sky130_fd_sc_hd__mux2_1
X_10887_ sub1.data_o\[112\] _06513_ _06632_ _06633_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06634_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15414_ _05202_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__clkbuf_4
X_18202_ clknet_leaf_16_clk _01633_ net637 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12626_ _07607_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__clkbuf_1
X_16394_ _04275_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18133_ clknet_leaf_28_clk _01576_ net643 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[87\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15345_ _03565_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12557_ _07571_ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11508_ _07017_ vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__clkbuf_1
X_18064_ net573 _01507_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[66\]
+ sky130_fd_sc_hd__dfxtp_1
X_15276_ _03441_ _03524_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__xnor2_4
X_12488_ _07535_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 mix1.data_reg\[80\] vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17015_ net407 _00458_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold119 mix1.data_reg\[37\] vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__dlygate4sd3_1
X_14227_ fifo_bank_register.bank\[6\]\[74\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[74\]
+ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a22o_1
X_11439_ _06981_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14158_ fifo_bank_register.bank\[5\]\[67\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[67\]
+ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13109_ fifo_bank_register.bank\[1\]\[81\] _05441_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14089_ fifo_bank_register.bank\[9\]\[59\] _02388_ _02463_ _02464_ _02465_ vssd1
+ vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_225_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ net575 _01360_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08650_ sub1.state\[1\] _04673_ sub1.state\[3\] sub1.state\[2\] vssd1 vssd1 vccd1
+ vccd1 _04674_ sky130_fd_sc_hd__and4b_1
X_17848_ net457 _01291_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08581_ _04609_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_135_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17779_ net405 _01222_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09202_ _05206_ _05211_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09133_ _05141_ _05143_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09064_ _05058_ _05077_ _05078_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09966_ sub1.data_o\[21\] _05803_ _05701_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08917_ addroundkey_data_o\[45\] _04693_ _04695_ addroundkey_data_o\[37\] vssd1 vssd1
+ vccd1 vccd1 _04941_ sky130_fd_sc_hd__a22o_1
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _05741_ vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__clkbuf_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__inv_2
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _04655_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10810_ sub1.data_o\[104\] _06564_ _06318_ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__mux2_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11790_ fifo_bank_register.bank\[6\]\[99\] _05478_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07166_ sky130_fd_sc_hd__mux2_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10741_ sub1.data_o\[98\] _06501_ _06478_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _08047_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__clkbuf_1
X_10672_ net119 mix1.data_o\[91\] _06316_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12411_ _07494_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13391_ _08011_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_20_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15130_ _03372_ _03397_ _03398_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__a21oi_1
X_12342_ _07457_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15061_ addroundkey_data_o\[92\] _03144_ _03145_ addroundkey_data_o\[60\] vssd1 vssd1
+ vccd1 vccd1 _03333_ sky130_fd_sc_hd__a22o_1
X_12273_ _07421_ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14012_ _02153_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11224_ _05455_ fifo_bank_register.bank\[8\]\[88\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ _05386_ fifo_bank_register.bank\[8\]\[55\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06831_ sky130_fd_sc_hd__mux2_1
XTAP_6141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10106_ _05899_ _05925_ _05929_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_207_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11086_ _05317_ fifo_bank_register.bank\[8\]\[22\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15963_ net221 ks1.key_reg\[67\] _03918_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput240 key_i[84] vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__buf_4
XTAP_5462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput251 key_i[94] vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_4
XFILLER_0_216_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17702_ net445 _01145_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
X_10037_ sub1.data_o\[29\] _05866_ _05819_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__mux2_1
X_14914_ sub1.data_o\[78\] _03108_ _03066_ sub1.data_o\[46\] vssd1 vssd1 vccd1 vccd1
+ _03189_ sky130_fd_sc_hd__a22o_1
XTAP_5484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15894_ _05195_ sub1.data_o\[67\] _05200_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17633_ net486 _01076_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14845_ addroundkey_data_o\[86\] _03062_ _03091_ addroundkey_data_o\[54\] vssd1 vssd1
+ vccd1 vccd1 _03121_ sky130_fd_sc_hd__a22o_1
XFILLER_0_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14776_ _04617_ sub1.ready_o _04666_ addroundkey_ready_o vssd1 vssd1 vccd1 vccd1
+ _03052_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_81_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17564_ net538 _01007_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11988_ fifo_bank_register.bank\[5\]\[64\] _05405_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16515_ _04341_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__clkbuf_1
X_13727_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__clkbuf_4
X_10939_ _06630_ sub1.ready_o sub1.data_o\[117\] _05675_ vssd1 vssd1 vccd1 vccd1 _06681_
+ sky130_fd_sc_hd__a31o_1
X_17495_ net497 _00938_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13658_ fifo_bank_register.bank\[9\]\[12\] _08190_ _02079_ _02080_ _02081_ vssd1
+ vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__a2111o_1
X_16446_ _04303_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ fifo_bank_register.bank\[3\]\[101\] _05483_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16377_ net831 _04102_ _04264_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13589_ fifo_bank_register.bank\[1\]\[5\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_11_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15328_ _03556_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18116_ net457 _01559_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[118\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15259_ _03511_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__clkbuf_1
X_18047_ net429 _01490_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[49\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_160_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09820_ _05672_ vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__clkbuf_1
Xfanout407 net413 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__buf_2
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_201_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout429 net431 vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09751_ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08702_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09682_ _05170_ _05552_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_193_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08633_ _04656_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ addroundkey_data_o\[120\] fifo_bank_register.data_out\[120\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__mux2_4
XFILLER_0_221_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08495_ addroundkey_data_o\[87\] fifo_bank_register.data_out\[87\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__mux2_2
XFILLER_0_193_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09116_ _05124_ _05125_ _05126_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__o21a_2
XFILLER_0_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09047_ _05061_ _05066_ vssd1 vssd1 vccd1 vccd1 sbox1.ah\[2\] sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09949_ _05712_ _05787_ _05788_ _05716_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__a22o_1
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _07784_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__clkbuf_1
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _07230_ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__clkbuf_1
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _07747_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__clkbuf_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_301 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ fifo_bank_register.bank\[5\]\[119\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[119\]
+ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__a22o_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_212_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11842_ fifo_bank_register.bank\[6\]\[124\] _05530_ _07055_ vssd1 vssd1 vccd1 vccd1
+ _07193_ sky130_fd_sc_hd__mux2_1
XANTENNA_323 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_334 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_345 _04566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14561_ _02157_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__buf_4
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _07157_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__clkbuf_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _08084_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__clkbuf_1
X_16300_ _04224_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__clkbuf_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _06485_ _06486_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__xnor2_1
X_17280_ net555 _00723_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14492_ fifo_bank_register.bank\[6\]\[103\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[103\]
+ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16231_ _04175_ _04176_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__xor2_2
XFILLER_0_64_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13443_ _05504_ fifo_bank_register.bank\[0\]\[111\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08039_ sky130_fd_sc_hd__mux2_1
X_10655_ net116 mix1.data_o\[89\] _06316_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16162_ addroundkey_round\[0\] _04109_ _05538_ _04723_ vssd1 vssd1 vccd1 vccd1 _04113_
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13374_ _08002_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__clkbuf_1
X_10586_ sub1.data_o\[83\] _06361_ _06113_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15113_ _03383_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12325_ _07448_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16093_ net145 ks1.key_reg\[113\] _03905_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__mux2_2
XFILLER_0_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15044_ sub1.data_o\[107\] _03079_ _03316_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_121_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12256_ _07412_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ _06791_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__buf_4
X_12187_ _07364_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__buf_4
XFILLER_0_222_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11138_ _05369_ fifo_bank_register.bank\[8\]\[47\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16995_ net499 _00438_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11069_ _06785_ vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__clkbuf_1
X_15946_ _03917_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__xor2_2
XTAP_5281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_5292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15877_ sub1.data_o\[93\] _05227_ _04888_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__mux2_1
XTAP_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17616_ net496 _01059_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_14828_ addroundkey_data_o\[70\] _03062_ _03091_ addroundkey_data_o\[38\] vssd1 vssd1
+ vccd1 vccd1 _03104_ sky130_fd_sc_hd__a22o_1
X_18596_ clknet_leaf_65_clk _02025_ net604 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[123\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17547_ net513 _00990_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14759_ _03043_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08280_ net202 net213 net191 net180 vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__and4b_1
XFILLER_0_188_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17478_ net475 _00921_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16429_ _04215_ _04022_ _04294_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_229_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09803_ addroundkey_data_o\[4\] _05657_ next_addroundkey_ready_o vssd1 vssd1 vccd1
+ vccd1 _05658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09734_ round\[3\] _05590_ _05586_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_213_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09665_ addroundkey_round\[1\] _04637_ _04642_ _04749_ _05539_ vssd1 vssd1 vccd1
+ vccd1 _00137_ sky130_fd_sc_hd__a32o_1
XFILLER_0_213_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ _04640_ vssd1 vssd1 vccd1 vccd1 next_addroundkey_ready_o sky130_fd_sc_hd__buf_4
XFILLER_0_132_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ fifo_bank_register.bank\[9\]\[106\] _05493_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05494_ sky130_fd_sc_hd__mux2_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08547_ _04592_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08478_ _04478_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__buf_8
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10440_ sub1.data_o\[68\] _06230_ _06160_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10371_ _06170_ vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _07334_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13090_ fifo_bank_register.bank\[1\]\[72\] _05422_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12041_ _07298_ vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15800_ mix1.data_o\[100\] net709 _03830_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13992_ _02379_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__clkbuf_1
X_16780_ clknet_leaf_79_clk _00224_ net579 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[71\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_189_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15731_ _03795_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12943_ _07775_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__clkbuf_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ clknet_leaf_70_clk _01880_ net609 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[90\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _03759_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_120 mix1.data_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _07738_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__clkbuf_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_131 sub1.data_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17401_ net575 _00844_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_153 net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14613_ fifo_bank_register.bank\[5\]\[117\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[117\]
+ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__a22o_1
X_11825_ _07184_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18381_ clknet_leaf_36_clk _01811_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[66\]
+ sky130_fd_sc_hd__dfrtp_4
X_15593_ _03722_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_164 net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_175 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_186 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_197 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ net432 _00775_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
X_14544_ fifo_bank_register.bank\[9\]\[109\] _02793_ _02868_ _02869_ _02870_ vssd1
+ vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__a2111o_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11756_ _07148_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10707_ mix1.data_o\[95\] _06463_ _06320_ _06321_ sub1.data_o\[95\] vssd1 vssd1 vccd1
+ vccd1 _06471_ sky130_fd_sc_hd__a32o_1
XFILLER_0_165_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17263_ net398 _00706_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_14475_ fifo_bank_register.bank\[7\]\[101\] _02785_ _02794_ fifo_bank_register.bank\[2\]\[101\]
+ _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11687_ _07078_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__buf_4
XFILLER_0_183_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13426_ _05487_ fifo_bank_register.bank\[0\]\[103\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08030_ sky130_fd_sc_hd__mux2_1
X_16214_ _04161_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__clkbuf_1
X_10638_ mix1.data_o\[87\] _06129_ _06398_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__o21a_1
XFILLER_0_180_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17194_ net453 _00637_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16145_ ks1.key_reg\[22\] _04097_ _03958_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13357_ _05417_ fifo_bank_register.bank\[0\]\[70\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _07994_ sky130_fd_sc_hd__mux2_1
X_10569_ _06076_ _06340_ _06346_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_183_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12308_ _07439_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16076_ net234 ks1.key_reg\[79\] _03979_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13288_ _07957_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15027_ sub1.data_o\[98\] _03077_ _03299_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a21oi_2
X_12239_ _07403_ vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16978_ net500 _00421_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput4 data_i[102] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__buf_4
XFILLER_0_223_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15929_ ks1.col\[0\] _03903_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__xor2_1
XFILLER_0_211_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09450_ fifo_bank_register.bank\[9\]\[59\] _05394_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08401_ addroundkey_data_o\[42\] fifo_bank_register.data_out\[42\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__mux2_2
XFILLER_0_203_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09381_ net188 vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__buf_2
X_18579_ clknet_leaf_77_clk _02008_ net589 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[106\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08332_ addroundkey_data_o\[9\] fifo_bank_register.data_out\[9\] _04479_ vssd1 vssd1
+ vccd1 vccd1 _04480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08263_ net156 net158 net157 net155 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput330 net330 vssd1 vssd1 vccd1 vccd1 data_o[48] sky130_fd_sc_hd__clkbuf_4
Xoutput341 net341 vssd1 vssd1 vccd1 vccd1 data_o[58] sky130_fd_sc_hd__clkbuf_4
Xoutput352 net352 vssd1 vssd1 vccd1 vccd1 data_o[68] sky130_fd_sc_hd__clkbuf_4
Xoutput363 net363 vssd1 vssd1 vccd1 vccd1 data_o[78] sky130_fd_sc_hd__clkbuf_4
Xoutput374 net374 vssd1 vssd1 vccd1 vccd1 data_o[88] sky130_fd_sc_hd__clkbuf_4
Xoutput385 net385 vssd1 vssd1 vccd1 vccd1 data_o[98] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09717_ round\[1\] _04613_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__xor2_1
XFILLER_0_173_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09648_ fifo_bank_register.bank\[9\]\[123\] _05528_ _05269_ vssd1 vssd1 vccd1 vccd1
+ _05529_ sky130_fd_sc_hd__mux2_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _05482_ vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__clkbuf_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11610_ _07071_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__clkbuf_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12590_ fifo_bank_register.bank\[3\]\[92\] _05464_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11541_ _07034_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_175_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ fifo_bank_register.bank\[6\]\[78\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[78\]
+ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _06998_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ _05272_ fifo_bank_register.bank\[0\]\[1\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07917_ sky130_fd_sc_hd__mux2_1
X_10423_ sub1.data_o\[66\] _06215_ _06160_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__mux2_1
X_14191_ _02148_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_180_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13142_ fifo_bank_register.bank\[1\]\[97\] _05474_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10354_ net211 ks1.key_reg\[58\] _05997_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17950_ net541 _01393_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ fifo_bank_register.bank\[1\]\[64\] _05405_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07844_ sky130_fd_sc_hd__mux2_1
X_10285_ _05949_ _06089_ _06091_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16901_ net524 _00344_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_12024_ fifo_bank_register.bank\[5\]\[81\] _05441_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07290_ sky130_fd_sc_hd__mux2_1
X_17881_ net502 _01324_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_228_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16832_ clknet_leaf_69_clk _00276_ net604 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[123\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_206_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout590 net595 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_205_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16763_ clknet_leaf_70_clk _00207_ net608 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[54\]
+ sky130_fd_sc_hd__dfrtp_4
X_13975_ _02364_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18502_ clknet_leaf_58_clk _01931_ net618 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_214_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15714_ mix1.data_o\[59\] net743 _03786_ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12926_ _07765_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__clkbuf_1
X_16694_ clknet_leaf_72_clk _00141_ net594 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[121\]
+ sky130_fd_sc_hd__dfrtp_2
X_18433_ clknet_leaf_23_clk _01863_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[118\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_197_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15645_ _03750_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__clkbuf_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12857_ fifo_bank_register.bank\[2\]\[90\] _05459_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07730_ sky130_fd_sc_hd__mux2_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ clknet_leaf_35_clk _01794_ net667 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[49\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_189_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11808_ _07175_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__clkbuf_1
X_15576_ _03700_ _03709_ _05560_ _03713_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__a31o_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12788_ _07693_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17315_ net400 _00758_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ _07139_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__clkbuf_1
X_14527_ fifo_bank_register.bank\[0\]\[107\] _02855_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02856_ sky130_fd_sc_hd__mux2_1
X_18295_ clknet_leaf_47_clk _01726_ net651 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[61\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17246_ net485 _00689_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14458_ _02138_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13409_ _05470_ fifo_bank_register.bank\[0\]\[95\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14389_ _02733_ fifo_bank_register.data_out\[91\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02734_ sky130_fd_sc_hd__mux2_1
X_17177_ net561 _00620_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16128_ _04082_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08950_ addroundkey_data_o\[79\] mix1.data_o\[79\] _04778_ vssd1 vssd1 vccd1 vccd1
+ _04974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16059_ net140 ks1.key_reg\[109\] _03905_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08881_ _04706_ _04903_ _04904_ _04710_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09502_ net231 vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09433_ _05383_ vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09364_ fifo_bank_register.bank\[9\]\[31\] _05336_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08315_ _04470_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_20 _04541_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_192_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09295_ _05289_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_31 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_42 _05614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08246_ _04399_ _04400_ _04401_ _04402_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__or4_1
XANTENNA_53 addroundkey_data_o\[113\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_64 addroundkey_data_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 addroundkey_data_o\[50\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_86 addroundkey_data_o\[79\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_97 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10070_ _05895_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__xnor2_1
XTAP_5814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13760_ _02173_ fifo_bank_register.data_out\[22\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02174_ sky130_fd_sc_hd__mux2_1
X_10972_ mix1.data_o\[120\] _05676_ _06575_ _06576_ sub1.data_o\[120\] vssd1 vssd1
+ vccd1 vccd1 _06711_ sky130_fd_sc_hd__a32o_1
XFILLER_0_173_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ _07653_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13691_ fifo_bank_register.bank\[0\]\[16\] _02110_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15430_ _03603_ _04949_ _05228_ _03620_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ fifo_bank_register.bank\[3\]\[117\] _05516_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ _03573_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__clkbuf_1
X_12573_ fifo_bank_register.bank\[3\]\[84\] _05447_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17100_ net477 _00543_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11524_ fifo_bank_register.bank\[7\]\[101\] _05483_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07026_ sky130_fd_sc_hd__mux2_1
X_14312_ fifo_bank_register.bank\[9\]\[83\] _02631_ _02662_ _02663_ _02664_ vssd1
+ vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a2111o_1
X_15292_ _03482_ _03536_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__xnor2_2
X_18080_ net568 _01523_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17031_ net526 _00474_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
X_14243_ fifo_bank_register.bank\[6\]\[76\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[76\]
+ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11455_ _06989_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10406_ net89 mix1.data_o\[64\] _06158_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14174_ _02541_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__clkbuf_1
X_11386_ _06953_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13125_ fifo_bank_register.bank\[1\]\[89\] _05457_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07871_ sky130_fd_sc_hd__mux2_1
X_10337_ _06001_ _06137_ _06139_ _06005_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ net528 _01376_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
X_13056_ fifo_bank_register.bank\[1\]\[56\] _05388_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10268_ _05567_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12007_ fifo_bank_register.bank\[5\]\[73\] _05424_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ net420 _01307_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10199_ _06013_ _06014_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__xor2_1
XFILLER_0_206_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16815_ clknet_leaf_4_clk _00259_ net584 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[106\]
+ sky130_fd_sc_hd__dfrtp_4
X_17795_ net527 _01238_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16746_ clknet_leaf_45_clk _00190_ net653 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13958_ _02349_ fifo_bank_register.data_out\[44\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12909_ fifo_bank_register.bank\[2\]\[115\] _05512_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16677_ net435 _00125_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13889_ fifo_bank_register.bank\[9\]\[37\] _02226_ _02285_ _02286_ _02287_ vssd1
+ vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_14_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18416_ clknet_leaf_13_clk _01846_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[101\]
+ sky130_fd_sc_hd__dfrtp_2
X_15628_ _04379_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__buf_4
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18347_ clknet_leaf_18_clk _01777_ net637 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[32\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15559_ _03700_ _04935_ _05219_ _03702_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09080_ sbox1.ah\[1\] _05088_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18278_ clknet_leaf_5_clk _01709_ net592 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[44\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_83_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput40 data_i[1] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_2
XFILLER_0_163_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17229_ net479 _00672_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput51 data_i[2] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_2
Xinput62 data_i[3] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_4
XFILLER_0_163_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput73 data_i[4] vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_4
XFILLER_0_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput84 data_i[5] vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__clkbuf_4
Xinput95 data_i[6] vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09982_ net44 mix1.data_o\[23\] _05817_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08933_ ks1.key_reg\[21\] _04726_ _04956_ net171 vssd1 vssd1 vccd1 vccd1 _04957_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_200_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08864_ _04677_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ mix1.data_o\[83\] _04677_ _04661_ mix1.data_o\[19\] vssd1 vssd1 vccd1 vccd1
+ _04819_ sky130_fd_sc_hd__a22o_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09416_ fifo_bank_register.bank\[9\]\[48\] _05371_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09347_ net176 vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__buf_2
XFILLER_0_165_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ net202 vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__buf_2
X_08229_ net18 net17 net20 net19 vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11240_ _06875_ vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ _06839_ vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10122_ _05943_ _05944_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__xnor2_1
XTAP_5600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10053_ _05881_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__clkbuf_1
X_14930_ addroundkey_data_o\[25\] _04377_ _03086_ _03204_ vssd1 vssd1 vccd1 vccd1
+ _03205_ sky130_fd_sc_hd__a211o_1
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14861_ addroundkey_data_o\[125\] _03055_ _03136_ vssd1 vssd1 vccd1 vccd1 _03137_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_216_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ net395 _00048_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ fifo_bank_register.bank\[5\]\[29\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[29\]
+ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_215_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17580_ net464 _01023_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14792_ _03067_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16531_ net684 _03521_ _04343_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__mux2_1
X_13743_ fifo_bank_register.bank\[0\]\[20\] _02156_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02159_ sky130_fd_sc_hd__mux2_1
X_10955_ net150 ks1.key_reg\[118\] _04639_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__mux2_2
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16462_ net819 _04312_ _03957_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__mux2_1
X_10886_ mix1.data_o\[112\] _06494_ _05617_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13674_ fifo_bank_register.bank\[9\]\[14\] _08190_ _02093_ _02094_ _02095_ vssd1
+ vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_183_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18201_ clknet_leaf_12_clk _01632_ net622 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[95\]
+ sky130_fd_sc_hd__dfrtp_1
X_15413_ _03603_ _04949_ _05548_ _03608_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__a31o_1
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ fifo_bank_register.bank\[3\]\[109\] _05499_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07607_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16393_ ks1.key_reg\[93\] _04274_ _04264_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18132_ clknet_leaf_24_clk _01575_ net643 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[86\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_182_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15344_ net734 _03510_ _03560_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12556_ fifo_bank_register.bank\[3\]\[76\] _05430_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11507_ fifo_bank_register.bank\[7\]\[93\] _05466_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18063_ net567 _01506_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[65\]
+ sky130_fd_sc_hd__dfxtp_2
X_15275_ _03459_ _03523_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__xnor2_2
X_12487_ fifo_bank_register.bank\[3\]\[43\] _05361_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07535_ sky130_fd_sc_hd__mux2_1
Xhold109 mix1.data_reg\[118\] vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ net397 _00457_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11438_ fifo_bank_register.bank\[7\]\[60\] _05396_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06981_ sky130_fd_sc_hd__mux2_1
X_14226_ fifo_bank_register.bank\[7\]\[74\] _02542_ _02551_ fifo_bank_register.bank\[2\]\[74\]
+ _02587_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14157_ _02526_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11369_ _06944_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13108_ _07862_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__clkbuf_1
X_14088_ fifo_bank_register.bank\[1\]\[59\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[59\]
+ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ fifo_bank_register.bank\[1\]\[48\] _05371_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07826_ sky130_fd_sc_hd__mux2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ net555 _01359_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17847_ net469 _01290_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08580_ state vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__buf_4
XFILLER_0_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17778_ net389 _01221_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16729_ clknet_leaf_43_clk _00173_ net658 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09201_ _05207_ _05210_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09132_ sbox1.ah_reg\[0\] _05142_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09063_ _05058_ sbox1.ah\[0\] _05067_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09965_ net42 mix1.data_o\[21\] _05699_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08916_ mix1.data_o\[45\] _04693_ _04695_ mix1.data_o\[37\] vssd1 vssd1 vccd1 vccd1
+ _04940_ sky130_fd_sc_hd__a22o_1
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09896_ addroundkey_data_o\[14\] _05740_ _05697_ vssd1 vssd1 vccd1 vccd1 _05741_
+ sky130_fd_sc_hd__mux2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _04648_ _04860_ _04866_ _04870_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a211o_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08778_ addroundkey_data_o\[123\] mix1.data_o\[123\] _04657_ vssd1 vssd1 vccd1 vccd1
+ _04802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10740_ net126 mix1.data_o\[98\] _06476_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_836 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _06439_ vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12410_ fifo_bank_register.bank\[3\]\[7\] _05284_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13390_ _05451_ fifo_bank_register.bank\[0\]\[86\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ _05487_ fifo_bank_register.bank\[4\]\[103\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07457_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15060_ sub1.data_o\[124\] _03143_ _03331_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__a21oi_4
X_12272_ _05417_ fifo_bank_register.bank\[4\]\[70\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14011_ _02151_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_181_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11223_ _06866_ vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11154_ _06830_ vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__clkbuf_1
XTAP_6131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10105_ sub1.data_o\[35\] _05753_ _05927_ _05928_ _04611_ vssd1 vssd1 vccd1 vccd1
+ _05929_ sky130_fd_sc_hd__a221o_1
XTAP_5430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11085_ _06794_ vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__clkbuf_1
X_15962_ ks1.col\[3\] _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__xor2_4
XTAP_5441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput230 key_i[75] vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
Xinput241 key_i[85] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_218_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17701_ net400 _01144_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14913_ _03160_ _03187_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__xnor2_2
X_10036_ net50 mix1.data_o\[29\] _05817_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__mux2_1
Xinput252 key_i[95] vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__buf_2
XFILLER_0_222_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15893_ _03881_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17632_ net508 _01075_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14844_ sub1.data_o\[118\] _03077_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__a21oi_2
XTAP_4784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17563_ net540 _01006_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
X_14775_ _03051_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__clkbuf_1
X_11987_ _07270_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ net749 _03493_ _04332_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__mux2_1
X_13726_ _08098_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__buf_6
X_10938_ sub1.data_o\[117\] _06679_ _05608_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17494_ net492 _00937_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16445_ net846 _04084_ _04295_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__mux2_1
X_13657_ fifo_bank_register.bank\[1\]\[12\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__a22o_1
X_10869_ net142 ks1.key_reg\[110\] _06579_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12608_ _07598_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__clkbuf_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _04372_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__buf_4
XFILLER_0_183_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13588_ fifo_bank_register.bank\[6\]\[5\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18115_ net442 _01558_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[117\]
+ sky130_fd_sc_hd__dfxtp_1
X_15327_ net768 _03484_ _03549_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12539_ fifo_bank_register.bank\[3\]\[68\] _05413_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18046_ net415 _01489_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15258_ net747 _03510_ _03498_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14209_ fifo_bank_register.bank\[5\]\[72\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[72\]
+ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15189_ _03321_ _03352_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout408 net413 vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__clkbuf_2
Xfanout419 net444 vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_2
XFILLER_0_201_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09750_ _05608_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__buf_4
XFILLER_0_225_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08701_ _04724_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__clkbuf_4
X_09681_ _04649_ _05184_ _05550_ _05551_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__o22a_2
XFILLER_0_94_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_207_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08632_ _04655_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__buf_4
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08563_ _04600_ vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__buf_1
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _04564_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09115_ _05105_ sbox1.inversion_to_invert_var\[0\] sbox1.inversion_to_invert_var\[3\]
+ sbox1.inversion_to_invert_var\[1\] vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09046_ _05058_ _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09948_ mix1.data_o\[19\] _05677_ _05703_ _05704_ sub1.data_o\[19\] vssd1 vssd1 vccd1
+ vccd1 _05788_ sky130_fd_sc_hd__a32o_1
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _05724_ _05725_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__xor2_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ fifo_bank_register.bank\[5\]\[27\] _05327_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07230_ sky130_fd_sc_hd__mux2_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ fifo_bank_register.bank\[2\]\[106\] _05493_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07747_ sky130_fd_sc_hd__mux2_1
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_302 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_174_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _07192_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__clkbuf_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_346 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11772_ fifo_bank_register.bank\[6\]\[90\] _05459_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07157_ sky130_fd_sc_hd__mux2_1
X_14560_ fifo_bank_register.bank\[9\]\[110\] _02874_ _02879_ _02882_ _02885_ vssd1
+ vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__a2111o_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ fifo_bank_register.write_ptr\[2\] _05264_ _05266_ vssd1 vssd1 vccd1 vccd1
+ _08084_ sky130_fd_sc_hd__mux2_1
X_10723_ net253 ks1.key_reg\[96\] _06402_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ fifo_bank_register.bank\[7\]\[103\] _02785_ _02794_ fifo_bank_register.bank\[2\]\[103\]
+ _02823_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ net250 ks1.key_reg\[93\] _03979_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__mux2_1
X_10654_ _06424_ vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__clkbuf_1
X_13442_ _08038_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16161_ addroundkey_round\[2\] _04642_ _04644_ _05542_ vssd1 vssd1 vccd1 vccd1 _04112_
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13373_ _05434_ fifo_bank_register.bank\[0\]\[78\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _08002_ sky130_fd_sc_hd__mux2_1
X_10585_ net110 mix1.data_o\[83\] _06111_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15112_ net750 _03382_ _03171_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12324_ _05470_ fifo_bank_register.bank\[4\]\[95\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16092_ net701 _03901_ _04049_ _04050_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15043_ sub1.data_o\[11\] _03208_ _03059_ _03315_ vssd1 vssd1 vccd1 vccd1 _03316_
+ sky130_fd_sc_hd__a211o_1
X_12255_ _05401_ fifo_bank_register.bank\[4\]\[62\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ _06857_ vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__clkbuf_1
X_12186_ _07375_ vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__clkbuf_1
X_11137_ _06821_ vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16994_ net486 _00437_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11068_ _05299_ fifo_bank_register.bank\[8\]\[14\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06785_ sky130_fd_sc_hd__mux2_1
X_15945_ net219 ks1.key_reg\[65\] _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_190_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ _05851_ vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15876_ _03870_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__clkbuf_1
XTAP_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17615_ net479 _01058_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_14827_ sub1.data_o\[102\] _03055_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a21oi_4
X_18595_ clknet_leaf_69_clk _02024_ net607 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17546_ net522 _00989_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14758_ ks1.col\[31\] _05244_ _04911_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13709_ _02126_ fifo_bank_register.data_out\[18\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17477_ net443 _00920_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
X_14689_ fifo_bank_register.bank\[1\]\[126\] _08111_ _08114_ fifo_bank_register.bank\[8\]\[126\]
+ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16428_ net686 _03914_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16359_ _04255_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18029_ net438 _01472_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09802_ _05655_ _05656_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__xor2_1
XFILLER_0_226_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09733_ _05568_ _04623_ _05593_ _05573_ round\[2\] vssd1 vssd1 vccd1 vccd1 _00151_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09664_ addroundkey_round\[0\] addroundkey_round\[1\] vssd1 vssd1 vccd1 vccd1 _05539_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08615_ _04636_ _04637_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_210_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09595_ net137 vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__buf_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08546_ addroundkey_data_o\[111\] fifo_bank_register.data_out\[111\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_212_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08477_ _04555_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_175_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10370_ addroundkey_data_o\[59\] _06168_ _06169_ vssd1 vssd1 vccd1 vccd1 _06170_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09029_ ks1.key_reg\[18\] _04745_ _04746_ net167 vssd1 vssd1 vccd1 vccd1 _05051_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_104_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ fifo_bank_register.bank\[5\]\[89\] _05457_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1090 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13991_ _02378_ fifo_bank_register.data_out\[48\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15730_ mix1.data_o\[67\] mix1.data_reg\[67\] _03786_ vssd1 vssd1 vccd1 vccd1 _03795_
+ sky130_fd_sc_hd__mux2_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12942_ fifo_bank_register.bank\[1\]\[2\] _05274_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07775_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ mix1.data_o\[34\] net693 _03753_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__mux2_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_110 fifo_bank_register.data_out\[88\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ fifo_bank_register.bank\[2\]\[98\] _05476_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_121 mix1.data_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 sub1.data_o\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ net572 _00843_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_143 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14612_ _02931_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__clkbuf_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ clknet_leaf_30_clk _01810_ net635 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[65\]
+ sky130_fd_sc_hd__dfrtp_4
X_11824_ fifo_bank_register.bank\[6\]\[115\] _05512_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07184_ sky130_fd_sc_hd__mux2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ mix1.data_o\[2\] _03283_ mix1.next_ready_o vssd1 vssd1 vccd1 vccd1 _03722_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_154 net78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_165 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_176 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_187 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ net454 _00774_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_198 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ fifo_bank_register.bank\[1\]\[109\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[109\]
+ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__a22o_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11755_ fifo_bank_register.bank\[6\]\[82\] _05443_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ sub1.data_o\[95\] _06469_ _06318_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__mux2_1
X_17262_ net392 _00705_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14474_ fifo_bank_register.bank\[5\]\[101\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[101\]
+ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11686_ _07111_ vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16213_ net795 _04160_ _04106_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__mux2_1
X_13425_ _08029_ vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__clkbuf_1
X_10637_ _06126_ _06407_ _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__a21o_1
X_17193_ net446 _00636_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16144_ _04868_ _04096_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__xnor2_1
X_10568_ sub1.data_o\[81\] _06341_ _06344_ _06345_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06346_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13356_ _07937_ vssd1 vssd1 vccd1 vccd1 _07993_ sky130_fd_sc_hd__buf_4
XFILLER_0_52_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12307_ _05453_ fifo_bank_register.bank\[4\]\[87\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16075_ net199 ks1.key_reg\[47\] _03982_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__mux2_1
X_13287_ _05348_ fifo_bank_register.bank\[0\]\[37\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07957_ sky130_fd_sc_hd__mux2_1
X_10499_ net229 ks1.key_reg\[74\] _06245_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__mux2_1
X_15026_ sub1.data_o\[2\] _04375_ _04658_ _03298_ vssd1 vssd1 vccd1 vccd1 _03299_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_220_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12238_ _05384_ fifo_bank_register.bank\[4\]\[54\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _05315_ fifo_bank_register.bank\[4\]\[21\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16977_ net503 _00420_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput5 data_i[103] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_4
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15928_ net253 ks1.key_reg\[96\] _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_190_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15859_ _04652_ _03862_ _04673_ _05104_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__o211a_1
XFILLER_0_203_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ _04515_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09380_ _05347_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__clkbuf_1
X_18578_ clknet_leaf_64_clk _02007_ net603 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[105\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08331_ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17529_ net570 _00972_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08262_ _04415_ _04416_ _04417_ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__or4_1
XFILLER_0_131_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_229_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput320 net320 vssd1 vssd1 vccd1 vccd1 data_o[39] sky130_fd_sc_hd__clkbuf_4
Xoutput331 net331 vssd1 vssd1 vccd1 vccd1 data_o[49] sky130_fd_sc_hd__buf_2
Xoutput342 net342 vssd1 vssd1 vccd1 vccd1 data_o[59] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput353 net353 vssd1 vssd1 vccd1 vccd1 data_o[69] sky130_fd_sc_hd__clkbuf_4
Xoutput364 net364 vssd1 vssd1 vccd1 vccd1 data_o[79] sky130_fd_sc_hd__clkbuf_4
Xoutput375 net375 vssd1 vssd1 vccd1 vccd1 data_o[89] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput386 net386 vssd1 vssd1 vccd1 vccd1 data_o[99] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09716_ _05575_ _05577_ _04629_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a21o_1
XFILLER_0_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09647_ net156 vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09578_ fifo_bank_register.bank\[9\]\[100\] _05480_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ addroundkey_data_o\[103\] fifo_bank_register.data_out\[103\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__mux2_2
XFILLER_0_195_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11540_ fifo_bank_register.bank\[7\]\[109\] _05499_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11471_ fifo_bank_register.bank\[7\]\[76\] _05430_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _06998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10422_ net91 mix1.data_o\[66\] _06158_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__mux2_1
X_13210_ _07916_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14190_ _02146_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10353_ _06001_ _06152_ _06153_ _06005_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__a22o_1
X_13141_ _07879_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13072_ _07843_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__clkbuf_1
X_10284_ _06090_ _05972_ sub1.data_o\[52\] _06079_ vssd1 vssd1 vccd1 vccd1 _06091_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12023_ _07289_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__clkbuf_1
X_16900_ net511 _00343_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_1282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17880_ net535 _01323_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16831_ clknet_leaf_74_clk _00275_ net587 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[122\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout580 net596 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__buf_2
XFILLER_0_219_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout591 net595 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_4
X_16762_ clknet_leaf_38_clk _00206_ net668 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[53\]
+ sky130_fd_sc_hd__dfrtp_2
X_13974_ _02363_ fifo_bank_register.data_out\[46\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18501_ clknet_leaf_58_clk _01930_ net618 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_219_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15713_ _03741_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12925_ fifo_bank_register.bank\[2\]\[123\] _05528_ _07628_ vssd1 vssd1 vccd1 vccd1
+ _07765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16693_ clknet_leaf_5_clk _00140_ net592 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18432_ clknet_leaf_24_clk _01862_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[117\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15644_ mix1.data_o\[26\] _03521_ _03742_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__mux2_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _07651_ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__buf_4
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18363_ clknet_leaf_15_clk _01793_ net630 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[48\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ fifo_bank_register.bank\[6\]\[107\] _05495_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07175_ sky130_fd_sc_hd__mux2_1
X_15575_ sub1.data_o\[10\] _03660_ _03710_ sub1.data_o\[74\] vssd1 vssd1 vccd1 vccd1
+ _03713_ sky130_fd_sc_hd__a22o_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ fifo_bank_register.bank\[2\]\[57\] _05390_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ net403 _00757_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ fifo_bank_register.bank\[9\]\[107\] _02793_ _02852_ _02853_ _02854_ vssd1
+ vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a2111o_1
X_18294_ clknet_leaf_45_clk _01725_ net652 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11738_ fifo_bank_register.bank\[6\]\[74\] _05426_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17245_ net487 _00688_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14457_ _02136_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11669_ fifo_bank_register.bank\[6\]\[41\] _05357_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13408_ _08020_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__clkbuf_1
X_17176_ net550 _00619_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14388_ fifo_bank_register.bank\[0\]\[91\] _02732_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02733_ sky130_fd_sc_hd__mux2_2
XFILLER_0_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16127_ ks1.key_reg\[20\] _04081_ _03958_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13339_ _07984_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16058_ net232 ks1.key_reg\[77\] _03918_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15009_ _03266_ _03282_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_138_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08880_ addroundkey_data_o\[8\] mix1.data_o\[8\] _04702_ vssd1 vssd1 vccd1 vccd1
+ _04904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09501_ _05429_ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09432_ fifo_bank_register.bank\[9\]\[53\] _05382_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09363_ net182 vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ addroundkey_data_o\[1\] fifo_bank_register.data_out\[1\] _04468_ vssd1 vssd1
+ vccd1 vccd1 _04470_ sky130_fd_sc_hd__mux2_2
X_09294_ fifo_bank_register.bank\[9\]\[9\] _05288_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_10 _03926_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _04562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08245_ net57 net56 net59 net58 vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__or4_1
XANTENNA_43 _05614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_54 addroundkey_data_o\[119\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_954 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_65 addroundkey_data_o\[34\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_76 addroundkey_data_o\[50\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_87 addroundkey_data_o\[79\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_98 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_219_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10971_ sub1.data_o\[120\] _06709_ _06573_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12710_ fifo_bank_register.bank\[2\]\[20\] _05311_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07653_ sky130_fd_sc_hd__mux2_1
X_13690_ fifo_bank_register.bank\[9\]\[16\] _08190_ _02107_ _02108_ _02109_ vssd1
+ vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12641_ _07615_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15360_ mix1.data_reg\[63\] _03537_ _03145_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12572_ _07579_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14311_ fifo_bank_register.bank\[1\]\[83\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[83\]
+ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11523_ _07025_ vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__clkbuf_1
X_15291_ _03410_ _03535_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_948 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17030_ net514 _00473_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14242_ fifo_bank_register.bank\[7\]\[76\] _02542_ _02551_ fifo_bank_register.bank\[2\]\[76\]
+ _02601_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__a221o_1
XFILLER_0_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11454_ fifo_bank_register.bank\[7\]\[68\] _05413_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10405_ _06200_ vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11385_ fifo_bank_register.bank\[7\]\[35\] _05344_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06953_ sky130_fd_sc_hd__mux2_1
X_14173_ _02540_ fifo_bank_register.data_out\[68\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124_ _07870_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10336_ mix1.data_o\[56\] _06138_ _05993_ _05994_ sub1.data_o\[56\] vssd1 vssd1 vccd1
+ vccd1 _06139_ sky130_fd_sc_hd__a32o_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _06075_ vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__clkbuf_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ net519 _01375_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
X_13055_ _07834_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__clkbuf_1
X_12006_ _07280_ vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__clkbuf_1
X_17863_ net439 _01306_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_10198_ net195 ks1.key_reg\[43\] _05997_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16814_ clknet_leaf_74_clk _00258_ net591 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[105\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_195_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17794_ net514 _01237_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16745_ clknet_leaf_48_clk _00189_ net611 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[36\]
+ sky130_fd_sc_hd__dfrtp_4
X_13957_ fifo_bank_register.bank\[0\]\[44\] _02348_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_979 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12908_ _07756_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16676_ net411 _00124_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13888_ fifo_bank_register.bank\[1\]\[37\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[37\]
+ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15627_ _03740_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18415_ clknet_leaf_13_clk _01845_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[100\]
+ sky130_fd_sc_hd__dfrtp_4
X_12839_ _07720_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__clkbuf_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ clknet_leaf_11_clk _01776_ net623 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15558_ sub1.data_o\[68\] _03691_ _03701_ _03673_ vssd1 vssd1 vccd1 vccd1 _03702_
+ sky130_fd_sc_hd__a22o_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14509_ fifo_bank_register.bank\[1\]\[105\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[105\]
+ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18277_ clknet_leaf_3_clk _01708_ net583 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[43\]
+ sky130_fd_sc_hd__dfrtp_4
X_15489_ _03652_ _04784_ _05196_ _03657_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17228_ net479 _00671_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput30 data_i[126] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__buf_4
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput41 data_i[20] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput52 data_i[30] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_4
Xinput63 data_i[40] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_2
XFILLER_0_124_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput74 data_i[50] vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_4
X_17159_ net518 _00602_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput85 data_i[60] vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput96 data_i[70] vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_2
XFILLER_0_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09981_ _05603_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08932_ ks1.key_reg\[21\] _04730_ _04732_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__or3_1
XFILLER_0_196_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08863_ _04884_ _04885_ _04886_ _04675_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08794_ addroundkey_data_o\[83\] _04677_ _04661_ addroundkey_data_o\[19\] vssd1 vssd1
+ vccd1 vccd1 _04818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ net200 vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__buf_4
XFILLER_0_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _05324_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09277_ _05277_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08228_ net14 net13 net16 net15 vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11170_ _05401_ fifo_bank_register.bank\[8\]\[62\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10121_ net187 ks1.key_reg\[36\] _05920_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__mux2_2
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10052_ addroundkey_data_o\[30\] _05880_ _05872_ vssd1 vssd1 vccd1 vccd1 _05881_
+ sky130_fd_sc_hd__mux2_1
XTAP_5634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14860_ addroundkey_data_o\[29\] _03100_ _05606_ _03135_ vssd1 vssd1 vccd1 vccd1
+ _03136_ sky130_fd_sc_hd__a211o_1
XTAP_5689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ _08181_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__buf_4
XTAP_4977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14791_ _03066_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__buf_4
XTAP_4999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ _04349_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13742_ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__buf_4
X_10954_ _05623_ _06690_ _06694_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_196_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16461_ _04165_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13673_ fifo_bank_register.bank\[1\]\[14\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a22o_1
X_10885_ _06491_ _06629_ _06631_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18200_ clknet_leaf_11_clk _01631_ net622 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15412_ sub1.data_o\[16\] _03606_ _03607_ sub1.next_ready_o vssd1 vssd1 vccd1 vccd1
+ _03608_ sky130_fd_sc_hd__a22o_1
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12624_ _07606_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__clkbuf_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16392_ _04177_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__inv_2
XFILLER_0_182_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18131_ clknet_leaf_22_clk _01574_ net643 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[85\]
+ sky130_fd_sc_hd__dfrtp_4
X_15343_ _03564_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12555_ _07570_ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18062_ net512 _01505_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[64\]
+ sky130_fd_sc_hd__dfxtp_2
X_11506_ _07016_ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__clkbuf_1
X_15274_ _03297_ _03453_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12486_ _07534_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17013_ net396 _00456_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_14225_ fifo_bank_register.bank\[5\]\[74\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[74\]
+ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11437_ _06935_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__buf_4
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14156_ _02525_ fifo_bank_register.data_out\[66\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02526_ sky130_fd_sc_hd__mux2_1
X_11368_ fifo_bank_register.bank\[7\]\[27\] _05327_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13107_ fifo_bank_register.bank\[1\]\[80\] _05438_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07862_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10319_ _06123_ vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14087_ fifo_bank_register.bank\[6\]\[59\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[59\]
+ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__a22o_1
X_11299_ _05530_ fifo_bank_register.bank\[8\]\[124\] _06768_ vssd1 vssd1 vccd1 vccd1
+ _06906_ sky130_fd_sc_hd__mux2_1
X_17915_ net567 _01358_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_13038_ _07825_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17846_ net433 _01289_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14989_ addroundkey_data_o\[122\] _03077_ _03262_ vssd1 vssd1 vccd1 vccd1 _03263_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17777_ net393 _01220_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16728_ clknet_leaf_41_clk _00172_ net659 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16659_ net447 _00107_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09200_ _05208_ _05209_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__xor2_1
XFILLER_0_174_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09131_ _05133_ _05131_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__or2b_1
XFILLER_0_134_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18329_ clknet_leaf_11_clk _01759_ net628 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09062_ sbox1.ah\[0\] sbox1.next_alph\[0\] vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09964_ _05802_ vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08915_ _04928_ _04931_ _04934_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__or4_1
XFILLER_0_228_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09895_ _05738_ _05739_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__xor2_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08846_ _04741_ _04868_ _04869_ _04750_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _04798_ _04738_ _04721_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_174_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10670_ addroundkey_data_o\[90\] _06438_ _06431_ vssd1 vssd1 vccd1 vccd1 _06439_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__buf_4
XFILLER_0_164_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12340_ _07456_ vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12271_ _07364_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__buf_4
XFILLER_0_121_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14010_ fifo_bank_register.bank\[6\]\[50\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[50\]
+ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11222_ _05453_ fifo_bank_register.bank\[8\]\[87\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11153_ _05384_ fifo_bank_register.bank\[8\]\[54\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06830_ sky130_fd_sc_hd__mux2_1
XTAP_6121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_6143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10104_ mix1.data_o\[35\] _05576_ _05916_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__o21a_1
X_11084_ _05315_ fifo_bank_register.bank\[8\]\[21\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06794_ sky130_fd_sc_hd__mux2_1
X_15961_ net256 ks1.key_reg\[99\] _03905_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__mux2_2
XFILLER_0_207_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput220 key_i[66] vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__buf_4
XTAP_5431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput231 key_i[76] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
Xinput242 key_i[86] vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_4
XTAP_5453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14912_ _03183_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__nor2_8
X_10035_ _05865_ vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__clkbuf_1
X_17700_ net447 _01143_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput253 key_i[96] vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__buf_4
XTAP_4730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15892_ sub1.data_o\[98\] _03880_ _03876_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__mux2_1
XTAP_5475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14843_ sub1.data_o\[22\] _03100_ _03058_ _03118_ vssd1 vssd1 vccd1 vccd1 _03119_
+ sky130_fd_sc_hd__a211o_1
X_17631_ net508 _01074_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17562_ net537 _01005_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
X_14774_ ks1.col\[23\] _05244_ _00007_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11986_ fifo_bank_register.bank\[5\]\[63\] _05403_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07270_ sky130_fd_sc_hd__mux2_1
X_16513_ _04340_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13725_ _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ net20 mix1.data_o\[117\] _05602_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__mux2_1
X_17493_ net503 _00936_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ _04302_ vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ fifo_bank_register.bank\[6\]\[12\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__a22o_1
X_10868_ _06583_ _06615_ _06616_ _06587_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ fifo_bank_register.bank\[3\]\[100\] _05480_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16375_ _04263_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13587_ fifo_bank_register.bank\[7\]\[5\] _08078_ _08093_ fifo_bank_register.bank\[2\]\[5\]
+ _08152_ vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10799_ sub1.data_o\[103\] _06554_ _06478_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__mux2_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18114_ net457 _01557_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[116\]
+ sky130_fd_sc_hd__dfxtp_1
X_15326_ _03555_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12538_ _07561_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18045_ net395 _01488_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15257_ _03196_ _03509_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__xnor2_4
X_12469_ _07525_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14208_ _02572_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15188_ _03386_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ fifo_bank_register.bank\[0\]\[64\] _02510_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout409 net413 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__buf_2
XFILLER_0_123_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08700_ _04644_ _04722_ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a21oi_1
X_09680_ _05154_ _05243_ _05060_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_1208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08631_ _04654_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__clkbuf_4
X_17829_ net402 _01272_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
X_08562_ addroundkey_data_o\[119\] fifo_bank_register.data_out\[119\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__mux2_2
XFILLER_0_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08493_ addroundkey_data_o\[86\] fifo_bank_register.data_out\[86\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__mux2_2
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09114_ _05105_ sbox1.inversion_to_invert_var\[0\] _05115_ vssd1 vssd1 vccd1 vccd1
+ _05125_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09045_ _05060_ _05062_ _05063_ _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__a31o_4
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09947_ sub1.data_o\[19\] _05786_ _05701_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ net161 ks1.key_reg\[12\] _05708_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__mux2_1
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ addroundkey_data_o\[110\] mix1.data_o\[110\] _04665_ vssd1 vssd1 vccd1 vccd1
+ _04853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ fifo_bank_register.bank\[6\]\[123\] _05528_ _07055_ vssd1 vssd1 vccd1 vccd1
+ _07192_ sky130_fd_sc_hd__mux2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_314 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_325 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_336 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_347 _06705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _07078_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__buf_4
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _08083_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__clkbuf_1
X_10722_ _06381_ _06479_ _06484_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_165_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14490_ fifo_bank_register.bank\[5\]\[103\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[103\]
+ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_165_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13441_ _05501_ fifo_bank_register.bank\[0\]\[110\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08038_ sky130_fd_sc_hd__mux2_1
X_10653_ addroundkey_data_o\[88\] _06423_ _06327_ vssd1 vssd1 vccd1 vccd1 _06424_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16160_ _04108_ _04109_ _04110_ _04723_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__a211o_2
XFILLER_0_36_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13372_ _08001_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10584_ _06360_ vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15111_ _03372_ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12323_ _07447_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__clkbuf_1
X_16091_ _04915_ _04048_ _03914_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15042_ sub1.data_o\[75\] _03064_ _03084_ sub1.data_o\[43\] vssd1 vssd1 vccd1 vccd1
+ _03315_ sky130_fd_sc_hd__a22o_1
X_12254_ _07411_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11205_ _05436_ fifo_bank_register.bank\[8\]\[79\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12185_ _05331_ fifo_bank_register.bank\[4\]\[29\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11136_ _05367_ fifo_bank_register.bank\[8\]\[46\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06821_ sky130_fd_sc_hd__mux2_1
X_16993_ net486 _00436_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ _06784_ vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__clkbuf_1
X_15944_ _03905_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__buf_4
XTAP_5261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10018_ addroundkey_data_o\[26\] _05850_ _05793_ vssd1 vssd1 vccd1 vccd1 _05851_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15875_ sub1.data_o\[92\] _05218_ _04888_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__mux2_1
XTAP_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14826_ sub1.data_o\[6\] _03100_ _03058_ _03101_ vssd1 vssd1 vccd1 vccd1 _03102_
+ sky130_fd_sc_hd__a211o_1
XTAP_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17614_ net480 _01057_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18594_ clknet_leaf_69_clk _02023_ net608 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14757_ _03042_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__clkbuf_1
X_17545_ net515 _00988_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11969_ fifo_bank_register.bank\[5\]\[55\] _05386_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13708_ fifo_bank_register.bank\[0\]\[18\] _02125_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17476_ net495 _00919_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14688_ fifo_bank_register.bank\[6\]\[126\] _08104_ _08107_ fifo_bank_register.bank\[4\]\[126\]
+ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13639_ _08114_ vssd1 vssd1 vccd1 vccd1 _08200_ sky130_fd_sc_hd__clkbuf_4
X_16427_ _04215_ _04012_ _04293_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16358_ net817 _04030_ _04252_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15309_ _03546_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16289_ _04218_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18028_ net438 _01471_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[30\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09801_ net202 ks1.key_reg\[4\] _05625_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09732_ _05586_ _05587_ _05589_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__o31a_1
XFILLER_0_198_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09663_ addroundkey_round\[0\] _04637_ _04723_ _05538_ vssd1 vssd1 vccd1 vccd1 _00136_
+ sky130_fd_sc_hd__a211o_1
X_08614_ _04638_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09594_ _05492_ vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ _04591_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08476_ addroundkey_data_o\[78\] fifo_bank_register.data_out\[78\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ net180 ks1.key_reg\[2\] _04725_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13990_ fifo_bank_register.bank\[0\]\[48\] _02377_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12941_ _07774_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__clkbuf_1
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15660_ _03758_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _07737_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_100 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_111 fifo_bank_register.data_out\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_122 mix1.data_o\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14611_ _02930_ fifo_bank_register.data_out\[116\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02931_ sky130_fd_sc_hd__mux2_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_133 sub1.data_o\[47\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ _07183_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__clkbuf_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _03721_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_144 net28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_166 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ net447 _00773_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ fifo_bank_register.bank\[6\]\[109\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[109\]
+ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__a22o_1
XANTENNA_177 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_188 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11754_ _07147_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_199 net131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10705_ net123 mix1.data_o\[95\] _06316_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__mux2_1
X_17261_ net414 _00704_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14473_ _02808_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11685_ fifo_bank_register.bank\[6\]\[49\] _05373_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16212_ _04831_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__xnor2_1
X_13424_ _05485_ fifo_bank_register.bank\[0\]\[102\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10636_ _06395_ _06342_ sub1.data_o\[87\] _06384_ vssd1 vssd1 vccd1 vccd1 _06408_
+ sky130_fd_sc_hd__a31o_1
X_17192_ net447 _00635_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16143_ _04094_ _04095_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13355_ _07992_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__clkbuf_1
X_10567_ mix1.data_o\[81\] _06129_ _06093_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__o21a_1
XFILLER_0_183_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12306_ _07438_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16074_ net699 ks1.next_ready_o _04033_ _04034_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__o22a_1
X_13286_ _07956_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10498_ _06250_ _06281_ _06282_ _06254_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__a22o_1
X_15025_ sub1.data_o\[66\] _03062_ _03091_ sub1.data_o\[34\] vssd1 vssd1 vccd1 vccd1
+ _03298_ sky130_fd_sc_hd__a22o_1
X_12237_ _07402_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12168_ _07366_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11119_ _05350_ fifo_bank_register.bank\[8\]\[38\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06812_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16976_ net500 _00419_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_12099_ fifo_bank_register.bank\[5\]\[117\] _05516_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 data_i[104] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__buf_4
X_15927_ _04742_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__buf_4
XFILLER_0_223_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15858_ sub1.state\[4\] _03861_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14809_ addroundkey_data_o\[24\] _04376_ _03084_ addroundkey_data_o\[56\] vssd1 vssd1
+ vccd1 vccd1 _03085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18577_ clknet_leaf_75_clk _02006_ net587 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[104\]
+ sky130_fd_sc_hd__dfrtp_1
X_15789_ mix1.data_o\[95\] net725 _03819_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08330_ _04466_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__buf_6
X_17528_ net556 _00971_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08261_ net39 net38 net42 net41 vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17459_ net459 _00902_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput310 net310 vssd1 vssd1 vccd1 vccd1 data_o[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput321 net321 vssd1 vssd1 vccd1 vccd1 data_o[3] sky130_fd_sc_hd__clkbuf_4
Xoutput332 net332 vssd1 vssd1 vccd1 vccd1 data_o[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput343 net343 vssd1 vssd1 vccd1 vccd1 data_o[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput354 net354 vssd1 vssd1 vccd1 vccd1 data_o[6] sky130_fd_sc_hd__clkbuf_4
Xoutput365 net365 vssd1 vssd1 vccd1 vccd1 data_o[7] sky130_fd_sc_hd__clkbuf_4
Xoutput376 net376 vssd1 vssd1 vccd1 vccd1 data_o[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput387 net387 vssd1 vssd1 vccd1 vccd1 data_o[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09715_ _04613_ _05576_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__nand2_1
XFILLER_0_198_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09646_ _05527_ vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _05312_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__buf_4
XFILLER_0_179_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08528_ _04582_ vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08459_ _04546_ vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_2
XFILLER_0_108_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_3__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11470_ _06997_ vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10421_ _06214_ vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ fifo_bank_register.bank\[1\]\[96\] _05472_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07879_ sky130_fd_sc_hd__mux2_1
X_10352_ mix1.data_o\[58\] _06138_ _05993_ _05994_ sub1.data_o\[58\] vssd1 vssd1 vccd1
+ vccd1 _06153_ sky130_fd_sc_hd__a32o_1
XFILLER_0_103_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13071_ fifo_bank_register.bank\[1\]\[63\] _05403_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07843_ sky130_fd_sc_hd__mux2_1
X_10283_ _04624_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12022_ fifo_bank_register.bank\[5\]\[80\] _05438_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16830_ clknet_leaf_73_clk _00274_ net593 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[121\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_228_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout570 net576 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__buf_2
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_4
Xfanout592 net595 vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_2
X_16761_ clknet_leaf_68_clk _00205_ net609 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[52\]
+ sky130_fd_sc_hd__dfrtp_4
X_13973_ fifo_bank_register.bank\[0\]\[46\] _02362_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18500_ clknet_leaf_55_clk _01929_ net614 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_214_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15712_ _03785_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__clkbuf_1
X_12924_ _07764_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__clkbuf_1
X_16692_ clknet_leaf_50_clk _00139_ net616 vssd1 vssd1 vccd1 vccd1 addroundkey_round\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_220_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18431_ clknet_leaf_24_clk _01861_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[116\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_158_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15643_ _03749_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _07728_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__clkbuf_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11806_ _07174_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__clkbuf_1
X_18362_ clknet_leaf_0_clk _01792_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[47\]
+ sky130_fd_sc_hd__dfrtp_4
X_15574_ _03700_ _03709_ _05554_ _03712_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a31o_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _07692_ vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17313_ net401 _00756_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
X_14525_ fifo_bank_register.bank\[1\]\[107\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[107\]
+ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__a22o_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _07138_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__clkbuf_1
X_18293_ clknet_leaf_47_clk _01724_ net652 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[59\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_166_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17244_ net488 _00687_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14456_ _02792_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__clkbuf_1
X_11668_ _07102_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_226_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13407_ _05468_ fifo_bank_register.bank\[0\]\[94\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ _06392_ vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__clkbuf_1
X_17175_ net564 _00618_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14387_ fifo_bank_register.bank\[9\]\[91\] _02712_ _02729_ _02730_ _02731_ vssd1
+ vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a2111o_1
X_11599_ _07065_ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16126_ _04744_ _04080_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__xnor2_1
X_13338_ _05399_ fifo_bank_register.bank\[0\]\[61\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16057_ net197 ks1.key_reg\[45\] _03982_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13269_ _07947_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15008_ _03273_ _03281_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__xor2_4
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16959_ net490 _00402_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09500_ fifo_bank_register.bank\[9\]\[75\] _05428_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ net206 vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__clkbuf_4
X_18629_ clknet_leaf_23_clk _02058_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[122\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_172_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09362_ _05335_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08313_ _04469_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_1
XFILLER_0_129_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09293_ net257 vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__buf_2
XANTENNA_11 _04391_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_191_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_22 _04570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 _04601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ net53 net52 net55 net54 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__or4_1
XFILLER_0_145_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_44 _05614_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_55 addroundkey_data_o\[121\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_66 addroundkey_data_o\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_77 addroundkey_data_o\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_88 fifo_bank_register.data_out\[114\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_99 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10970_ net24 mix1.data_o\[120\] _06571_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09629_ net149 vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__buf_2
XFILLER_0_211_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12640_ fifo_bank_register.bank\[3\]\[116\] _05514_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12571_ fifo_bank_register.bank\[3\]\[83\] _05445_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14310_ fifo_bank_register.bank\[6\]\[83\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[83\]
+ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
X_11522_ fifo_bank_register.bank\[7\]\[100\] _05480_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07025_ sky130_fd_sc_hd__mux2_1
X_15290_ _03187_ _03418_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ fifo_bank_register.bank\[5\]\[76\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[76\]
+ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_184_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11453_ _06988_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10404_ addroundkey_data_o\[63\] _06199_ _06169_ vssd1 vssd1 vccd1 vccd1 _06200_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14172_ fifo_bank_register.bank\[0\]\[68\] _02539_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02540_ sky130_fd_sc_hd__mux2_1
X_11384_ _06952_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13123_ fifo_bank_register.bank\[1\]\[88\] _05455_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07870_ sky130_fd_sc_hd__mux2_1
X_10335_ _05585_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ net516 _01374_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
X_13054_ fifo_bank_register.bank\[1\]\[55\] _05386_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10266_ addroundkey_data_o\[50\] _06074_ _06064_ vssd1 vssd1 vccd1 vccd1 _06075_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ fifo_bank_register.bank\[5\]\[72\] _05422_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07280_ sky130_fd_sc_hd__mux2_1
X_17862_ net421 _01305_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10197_ _06001_ _06011_ _06012_ _06005_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__a22o_1
XFILLER_0_219_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16813_ clknet_leaf_74_clk _00257_ net591 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[104\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17793_ net572 _01236_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16744_ clknet_leaf_45_clk _00188_ net653 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[35\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_205_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13956_ fifo_bank_register.bank\[9\]\[44\] _02307_ _02345_ _02346_ _02347_ vssd1
+ vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_159_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12907_ fifo_bank_register.bank\[2\]\[114\] _05510_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13887_ fifo_bank_register.bank\[6\]\[37\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[37\]
+ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a22o_1
X_16675_ net470 _00123_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_201_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18414_ clknet_leaf_13_clk _01844_ net628 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[99\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15626_ mix1.data_o\[18\] _03493_ _03730_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__mux2_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ fifo_bank_register.bank\[2\]\[81\] _05441_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07720_ sky130_fd_sc_hd__mux2_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18345_ clknet_leaf_11_clk _01775_ net631 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15557_ sub1.data_o\[100\] sub1.data_o\[36\] _03671_ vssd1 vssd1 vccd1 vccd1 _03701_
+ sky130_fd_sc_hd__mux2_1
X_12769_ _07683_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__clkbuf_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clknet_3_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14508_ fifo_bank_register.bank\[6\]\[105\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[105\]
+ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__a22o_1
X_18276_ clknet_leaf_2_clk _01707_ net583 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[42\]
+ sky130_fd_sc_hd__dfrtp_4
X_15488_ sub1.data_o\[107\] _03600_ _03653_ sub1.data_o\[43\] vssd1 vssd1 vccd1 vccd1
+ _03657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput20 data_i[117] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_4
X_17227_ net476 _00670_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput31 data_i[127] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_4
X_14439_ _02777_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 data_i[21] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_4
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput53 data_i[31] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_163_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput64 data_i[41] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_4
XFILLER_0_130_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput75 data_i[51] vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_8
X_17158_ net514 _00601_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput86 data_i[61] vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_4
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput97 data_i[71] vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__buf_4
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16109_ ks1.key_reg\[18\] _04065_ _03958_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09980_ _05816_ vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__clkbuf_1
X_17089_ net440 _00532_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08931_ _04653_ _04924_ _04939_ _04954_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__a211o_2
XFILLER_0_228_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08862_ addroundkey_data_o\[24\] mix1.data_o\[24\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08793_ _04807_ _04810_ _04813_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__or4_1
XFILLER_0_93_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09414_ _05370_ vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09345_ fifo_bank_register.bank\[9\]\[25\] _05323_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09276_ fifo_bank_register.bank\[9\]\[3\] _05276_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08227_ net5 net4 net7 net6 vssd1 vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1053 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10120_ _05899_ _05937_ _05942_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_219_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10051_ _05878_ _05879_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13810_ _02217_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__clkbuf_1
XTAP_4978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__buf_4
XTAP_4989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ _08119_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__clkbuf_8
X_10953_ sub1.data_o\[118\] _05613_ _06692_ _06693_ _04610_ vssd1 vssd1 vccd1 vccd1
+ _06694_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13672_ fifo_bank_register.bank\[6\]\[14\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a22o_1
X_16460_ _04373_ _04155_ _04311_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_211_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10884_ _06630_ _06514_ sub1.data_o\[112\] _05675_ vssd1 vssd1 vccd1 vccd1 _06631_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15411_ sub1.data_o\[112\] sub1.data_o\[48\] _05598_ vssd1 vssd1 vccd1 vccd1 _03607_
+ sky130_fd_sc_hd__mux2_1
X_12623_ fifo_bank_register.bank\[3\]\[108\] _05497_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16391_ _04273_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__clkbuf_1
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_186_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15342_ net710 _03507_ _03560_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__mux2_1
X_18130_ clknet_leaf_28_clk _01573_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[84\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12554_ fifo_bank_register.bank\[3\]\[75\] _05428_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11505_ fifo_bank_register.bank\[7\]\[92\] _05464_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07016_ sky130_fd_sc_hd__mux2_1
X_15273_ _03522_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__clkbuf_1
X_18061_ net575 _01504_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12485_ fifo_bank_register.bank\[3\]\[42\] _05359_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17012_ net392 _00455_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_14224_ _02586_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11436_ _06979_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14155_ fifo_bank_register.bank\[0\]\[66\] _02524_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02525_ sky130_fd_sc_hd__mux2_1
X_11367_ _06943_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _07794_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ addroundkey_data_o\[54\] _06122_ _06064_ vssd1 vssd1 vccd1 vccd1 _06123_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14086_ fifo_bank_register.bank\[7\]\[59\] _02461_ _02389_ fifo_bank_register.bank\[2\]\[59\]
+ _02462_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a221o_1
X_11298_ _06905_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__clkbuf_1
X_17914_ net567 _01357_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_13037_ fifo_bank_register.bank\[1\]\[47\] _05369_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07825_ sky130_fd_sc_hd__mux2_1
X_10249_ mix1.data_o\[49\] _05952_ _05916_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17845_ net411 _01288_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17776_ net394 _01219_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_14988_ addroundkey_data_o\[26\] _04375_ _04900_ _03261_ vssd1 vssd1 vccd1 vccd1
+ _03262_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16727_ clknet_leaf_40_clk _00171_ net659 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_152_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13939_ fifo_bank_register.bank\[1\]\[42\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[42\]
+ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16658_ net449 _00106_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15609_ _03731_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16589_ net499 _00037_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_14_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09130_ sbox1.ah_reg\[2\] _05111_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__nand2_1
X_18328_ clknet_leaf_9_clk _01758_ net631 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ _04971_ _05016_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18259_ clknet_leaf_43_clk _01690_ net655 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_142_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09963_ addroundkey_data_o\[20\] _05801_ _05793_ vssd1 vssd1 vccd1 vccd1 _05802_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08914_ _04935_ _04936_ _04937_ _04689_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__a22o_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ net163 ks1.key_reg\[14\] _05708_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__mux2_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ net181 ks1.key_reg\[30\] _04725_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ ks1.key_reg\[3\] _04726_ _04799_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_212_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09328_ _05268_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__buf_6
XFILLER_0_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ fifo_bank_register.write_ptr\[3\] _05253_ _05252_ vssd1 vssd1 vccd1 vccd1
+ _05263_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _07419_ vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ _06865_ vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11152_ _06829_ vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__clkbuf_1
XTAP_6111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ _05575_ _05925_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__a21o_1
XFILLER_0_222_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11083_ _06793_ vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__clkbuf_1
X_15960_ net691 _03901_ _03931_ _03932_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a22o_1
Xinput210 key_i[57] vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_8
XTAP_5421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput221 key_i[67] vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_4
XTAP_5443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14911_ addroundkey_data_o\[119\] _03077_ _03185_ vssd1 vssd1 vccd1 vccd1 _03186_
+ sky130_fd_sc_hd__a21oi_2
X_10034_ addroundkey_data_o\[28\] _05864_ _05793_ vssd1 vssd1 vccd1 vccd1 _05865_
+ sky130_fd_sc_hd__mux2_1
Xinput232 key_i[77] vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
XTAP_5454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput243 key_i[87] vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput254 key_i[97] vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_4
XTAP_5465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15891_ _05559_ sub1.data_o\[66\] _05200_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__mux2_1
XTAP_5476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ net485 _01073_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14842_ sub1.data_o\[86\] _03062_ _03091_ sub1.data_o\[54\] vssd1 vssd1 vccd1 vccd1
+ _03118_ sky130_fd_sc_hd__a22o_1
XTAP_4753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17561_ net538 _01004_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11985_ _07269_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__clkbuf_1
X_14773_ _03050_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16512_ net738 _03491_ _04332_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__mux2_1
X_10936_ _06678_ vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__clkbuf_1
X_13724_ _08095_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__buf_6
X_17492_ net503 _00935_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_168_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_168_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16443_ net842 _04076_ _04295_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ mix1.data_o\[110\] _06463_ _06575_ _06576_ sub1.data_o\[110\] vssd1 vssd1
+ vccd1 vccd1 _06616_ sky130_fd_sc_hd__a32o_1
X_13655_ fifo_bank_register.bank\[7\]\[12\] _08182_ _08191_ fifo_bank_register.bank\[2\]\[12\]
+ _02078_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12606_ _07508_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__buf_4
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ fifo_bank_register.bank\[5\]\[5\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[5\]
+ vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16374_ net805 _04094_ _04252_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10798_ net5 mix1.data_o\[103\] _06476_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__mux2_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18113_ net471 _01556_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[115\]
+ sky130_fd_sc_hd__dfxtp_4
X_15325_ net730 _03477_ _03549_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__mux2_1
X_12537_ fifo_bank_register.bank\[3\]\[67\] _05411_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ net390 _01487_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15256_ _03168_ _03400_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__xor2_2
XFILLER_0_124_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12468_ fifo_bank_register.bank\[3\]\[34\] _05342_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14207_ _02571_ fifo_bank_register.data_out\[71\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02572_ sky130_fd_sc_hd__mux2_1
X_11419_ fifo_bank_register.bank\[7\]\[51\] _05378_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06971_ sky130_fd_sc_hd__mux2_1
X_15187_ _03421_ _03449_ _03450_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__o21a_1
XFILLER_0_160_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12399_ _07488_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14138_ fifo_bank_register.bank\[9\]\[64\] _02469_ _02507_ _02508_ _02509_ vssd1
+ vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14069_ fifo_bank_register.bank\[6\]\[57\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[57\]
+ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__a22o_1
XFILLER_0_225_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_clk clknet_3_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_225_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08630_ _04617_ _04616_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_206_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17828_ net454 _01271_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08561_ _04599_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__buf_2
XFILLER_0_222_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17759_ net488 _01202_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08492_ _04563_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09113_ sbox1.inversion_to_invert_var\[1\] _05105_ vssd1 vssd1 vccd1 vccd1 _05124_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09044_ _05060_ _05054_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09946_ net39 mix1.data_o\[19\] _05699_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__mux2_1
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _05712_ _05722_ _05723_ _05716_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__a22o_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ mix1.data_o\[102\] _04650_ _04701_ _04851_ vssd1 vssd1 vccd1 vccd1 _04852_
+ sky130_fd_sc_hd__o211a_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _04777_ _04779_ _04782_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__a21o_1
XANTENNA_304 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_315 net224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_326 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_337 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_348 addroundkey_data_o\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11770_ _07155_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__clkbuf_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ sub1.data_o\[96\] _06341_ _06481_ _06482_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06484_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ _07937_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__buf_4
XFILLER_0_193_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ _06421_ _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__xor2_1
XFILLER_0_193_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13371_ _05432_ fifo_bank_register.bank\[0\]\[77\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _08001_ sky130_fd_sc_hd__mux2_1
X_10583_ addroundkey_data_o\[82\] _06359_ _06327_ vssd1 vssd1 vccd1 vccd1 _06360_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15110_ _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__xor2_2
X_12322_ _05468_ fifo_bank_register.bank\[4\]\[94\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16090_ _04915_ _04048_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__or2_1
XFILLER_0_224_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15041_ _03310_ _03313_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__nor2_8
XFILLER_0_146_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12253_ _05399_ fifo_bank_register.bank\[4\]\[61\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07411_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11204_ _06856_ vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12184_ _07374_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11135_ _06820_ vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16992_ net508 _00435_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11066_ _05297_ fifo_bank_register.bank\[8\]\[13\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06784_ sky130_fd_sc_hd__mux2_1
X_15943_ ks1.col\[1\] _03916_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__xor2_4
XFILLER_0_223_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10017_ _05848_ _05849_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__xor2_1
XTAP_5284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _03869_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__clkbuf_1
XTAP_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17613_ net477 _01056_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14825_ sub1.data_o\[70\] _03062_ _03091_ sub1.data_o\[38\] vssd1 vssd1 vccd1 vccd1
+ _03101_ sky130_fd_sc_hd__a22o_1
XTAP_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18593_ clknet_leaf_65_clk _02022_ net604 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ net522 _00987_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ ks1.col\[30\] _05235_ _04911_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11968_ _07260_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13707_ fifo_bank_register.bank\[9\]\[18\] _08190_ _02122_ _02123_ _02124_ vssd1
+ vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_188_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10919_ mix1.data_o\[115\] _04626_ _05617_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__o21a_1
X_17475_ net495 _00918_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
X_11899_ _07224_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14687_ fifo_bank_register.bank\[7\]\[126\] _08077_ _08092_ fifo_bank_register.bank\[2\]\[126\]
+ _02996_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16426_ net678 _03914_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_172_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13638_ _08111_ vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16357_ _04254_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_229_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13569_ _08137_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15308_ net762 _03392_ _03539_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16288_ net818 _04217_ _04206_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18027_ net480 _01470_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_15239_ _03290_ _03374_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_164_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_199_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09800_ _05629_ _05653_ _05654_ _05633_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09731_ _05590_ _05591_ _05586_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_201_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09662_ addroundkey_round\[0\] _04644_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08613_ addroundkey_start_i _04615_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__nand2_2
XFILLER_0_59_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09593_ fifo_bank_register.bank\[9\]\[105\] _05491_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08544_ addroundkey_data_o\[110\] fifo_bank_register.data_out\[110\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__mux2_4
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ _04554_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__buf_1
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09027_ _04645_ _05046_ _05048_ _04755_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__o22a_1
XFILLER_0_182_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09929_ sub1.data_o\[17\] _05753_ _05769_ _05770_ _04611_ vssd1 vssd1 vccd1 vccd1
+ _05771_ sky130_fd_sc_hd__a221o_1
XFILLER_0_226_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12940_ fifo_bank_register.bank\[1\]\[1\] _05272_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07774_ sky130_fd_sc_hd__mux2_1
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12871_ fifo_bank_register.bank\[2\]\[97\] _05474_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07737_ sky130_fd_sc_hd__mux2_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_101 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_112 mix1.data_o\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 mix1.data_o\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ fifo_bank_register.bank\[0\]\[116\] _02929_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02930_ sky130_fd_sc_hd__mux2_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_134 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ fifo_bank_register.bank\[6\]\[114\] _05510_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07183_ sky130_fd_sc_hd__mux2_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ mix1.data_o\[1\] _03236_ mix1.next_ready_o vssd1 vssd1 vccd1 vccd1 _03721_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ fifo_bank_register.bank\[7\]\[109\] _02866_ _02794_ fifo_bank_register.bank\[2\]\[109\]
+ _02867_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__a221o_1
XANTENNA_178 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ fifo_bank_register.bank\[6\]\[81\] _05441_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07147_ sky130_fd_sc_hd__mux2_1
XANTENNA_189 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _06468_ vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17260_ net416 _00703_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11684_ _07110_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__clkbuf_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ _02807_ fifo_bank_register.data_out\[100\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16211_ _04157_ _04158_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_180_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10635_ sub1.data_o\[87\] _06406_ _06113_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13423_ _08028_ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17191_ net454 _00634_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ _05415_ fifo_bank_register.bank\[0\]\[69\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07992_ sky130_fd_sc_hd__mux2_1
X_16142_ net207 ks1.key_reg\[54\] _03982_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__mux2_1
X_10566_ _06126_ _06340_ _06343_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12305_ _05451_ fifo_bank_register.bank\[4\]\[86\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13285_ _05346_ fifo_bank_register.bank\[0\]\[36\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07956_ sky130_fd_sc_hd__mux2_1
X_16073_ _04862_ _04032_ _04371_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__a21o_1
X_10497_ mix1.data_o\[74\] _06217_ _06241_ _06242_ sub1.data_o\[74\] vssd1 vssd1 vccd1
+ vccd1 _06282_ sky130_fd_sc_hd__a32o_1
X_15024_ _03293_ _03296_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__nor2_4
X_12236_ _05382_ fifo_bank_register.bank\[4\]\[53\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12167_ _05311_ fifo_bank_register.bank\[4\]\[20\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07366_ sky130_fd_sc_hd__mux2_1
X_11118_ _06811_ vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16975_ net480 _00418_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_12098_ _07328_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11049_ _05280_ fifo_bank_register.bank\[8\]\[5\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06775_ sky130_fd_sc_hd__mux2_1
X_15926_ _04371_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 data_i[105] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_4
XTAP_5092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _04362_ _04363_ _04364_ _04365_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__or4_1
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14808_ _03066_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__buf_4
X_18576_ clknet_leaf_80_clk _02005_ net580 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[103\]
+ sky130_fd_sc_hd__dfrtp_1
X_15788_ _03825_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__clkbuf_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17527_ net405 _00970_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14739_ _03033_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08260_ net35 net34 net37 net36 vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__or4_1
XFILLER_0_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17458_ net452 _00901_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16409_ _04284_ vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17389_ net415 _00832_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput300 net300 vssd1 vssd1 vccd1 vccd1 data_o[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput311 net311 vssd1 vssd1 vccd1 vccd1 data_o[30] sky130_fd_sc_hd__buf_2
XFILLER_0_11_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput322 net322 vssd1 vssd1 vccd1 vccd1 data_o[40] sky130_fd_sc_hd__clkbuf_4
Xoutput333 net333 vssd1 vssd1 vccd1 vccd1 data_o[50] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput344 net344 vssd1 vssd1 vccd1 vccd1 data_o[60] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_199_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput355 net355 vssd1 vssd1 vccd1 vccd1 data_o[70] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput366 net366 vssd1 vssd1 vccd1 vccd1 data_o[80] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1098 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput377 net377 vssd1 vssd1 vccd1 vccd1 data_o[90] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput388 net388 vssd1 vssd1 vccd1 vccd1 ready_o sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_226_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09714_ _04626_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_184_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09645_ fifo_bank_register.bank\[9\]\[122\] _05526_ _05269_ vssd1 vssd1 vccd1 vccd1
+ _05527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ net131 vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__buf_2
XFILLER_0_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08527_ addroundkey_data_o\[102\] fifo_bank_register.data_out\[102\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__mux2_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08458_ addroundkey_data_o\[69\] fifo_bank_register.data_out\[69\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08389_ _04509_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10420_ addroundkey_data_o\[65\] _06213_ _06169_ vssd1 vssd1 vccd1 vccd1 _06214_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10351_ sub1.data_o\[58\] _06151_ _05991_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13070_ _07842_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__clkbuf_1
X_10282_ sub1.data_o\[52\] _06088_ _05936_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12021_ _07221_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__buf_4
XFILLER_0_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout560 net561 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__buf_2
XFILLER_0_219_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout571 net576 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_2
X_16760_ clknet_leaf_39_clk _00204_ net663 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[51\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout582 net585 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_2
X_13972_ fifo_bank_register.bank\[9\]\[46\] _02307_ _02359_ _02360_ _02361_ vssd1
+ vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a2111o_1
Xfanout593 net595 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_219_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15711_ mix1.data_o\[58\] net798 _03775_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__mux2_1
X_12923_ fifo_bank_register.bank\[2\]\[122\] _05526_ _07628_ vssd1 vssd1 vccd1 vccd1
+ _07764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16691_ clknet_leaf_50_clk _00138_ net616 vssd1 vssd1 vccd1 vccd1 addroundkey_round\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18430_ clknet_leaf_23_clk _01860_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[115\]
+ sky130_fd_sc_hd__dfrtp_2
X_15642_ mix1.data_o\[25\] _03516_ _03742_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12854_ fifo_bank_register.bank\[2\]\[89\] _05457_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07728_ sky130_fd_sc_hd__mux2_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_189_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18361_ clknet_leaf_84_clk _01791_ net582 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[46\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ fifo_bank_register.bank\[6\]\[106\] _05493_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15573_ sub1.data_o\[9\] _03660_ _03710_ sub1.data_o\[73\] vssd1 vssd1 vccd1 vccd1
+ _03712_ sky130_fd_sc_hd__a22o_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ fifo_bank_register.bank\[2\]\[56\] _05388_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07692_ sky130_fd_sc_hd__mux2_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ net409 _00755_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14524_ fifo_bank_register.bank\[6\]\[107\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[107\]
+ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a22o_1
X_18292_ clknet_leaf_46_clk _01723_ net651 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[58\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11736_ fifo_bank_register.bank\[6\]\[73\] _05424_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07138_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17243_ net487 _00686_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14455_ _02791_ fifo_bank_register.data_out\[99\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02792_ sky130_fd_sc_hd__mux2_1
X_11667_ fifo_bank_register.bank\[6\]\[40\] _05354_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13406_ _08019_ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__clkbuf_1
X_10618_ addroundkey_data_o\[85\] _06391_ _06327_ vssd1 vssd1 vccd1 vccd1 _06392_
+ sky130_fd_sc_hd__mux2_1
X_17174_ net565 _00617_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11598_ fifo_bank_register.bank\[6\]\[8\] _05286_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07065_ sky130_fd_sc_hd__mux2_1
X_14386_ fifo_bank_register.bank\[1\]\[91\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[91\]
+ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16125_ _04078_ _04079_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__xor2_2
X_10549_ _06328_ vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13337_ _07983_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16056_ _04018_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13268_ _05329_ fifo_bank_register.bank\[0\]\[28\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15007_ _03207_ _03280_ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_161_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12219_ _05365_ fifo_bank_register.bank\[4\]\[45\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13199_ _07909_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16958_ net442 _00401_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15909_ _04369_ _04943_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__nor2_2
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16889_ net572 _00332_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09430_ _05381_ vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__clkbuf_1
X_18628_ clknet_leaf_25_clk _02057_ net648 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[121\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ fifo_bank_register.bank\[9\]\[30\] _05333_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18559_ clknet_leaf_76_clk _01988_ net590 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[86\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08312_ addroundkey_data_o\[0\] fifo_bank_register.data_out\[0\] _04468_ vssd1 vssd1
+ vccd1 vccd1 _04469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09292_ _05287_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _04435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _04571_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ net44 net43 net46 net45 vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__or4_1
XANTENNA_34 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_45 _06051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 addroundkey_data_o\[121\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 addroundkey_data_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_78 addroundkey_data_o\[64\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_89 fifo_bank_register.data_out\[115\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_160_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09628_ _05515_ vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09559_ fifo_bank_register.bank\[9\]\[94\] _05468_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12570_ _07578_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11521_ _06935_ vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__buf_4
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11452_ fifo_bank_register.bank\[7\]\[67\] _05411_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06988_ sky130_fd_sc_hd__mux2_1
X_14240_ _02600_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10403_ _06197_ _06198_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14171_ fifo_bank_register.bank\[9\]\[68\] _02469_ _02536_ _02537_ _02538_ vssd1
+ vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_46_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11383_ fifo_bank_register.bank\[7\]\[34\] _05342_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10334_ sub1.data_o\[56\] _06136_ _05991_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__mux2_1
X_13122_ _07869_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__clkbuf_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17930_ net511 _01373_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
X_13053_ _07833_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__clkbuf_1
X_10265_ _06072_ _06073_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_218_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12004_ _07279_ vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__clkbuf_1
X_17861_ net471 _01304_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
X_10196_ mix1.data_o\[43\] _05876_ _05993_ _05994_ sub1.data_o\[43\] vssd1 vssd1 vccd1
+ vccd1 _06012_ sky130_fd_sc_hd__a32o_1
XFILLER_0_187_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16812_ clknet_leaf_75_clk _00256_ net586 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[103\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17792_ net558 _01235_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout390 net391 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__buf_1
XFILLER_0_75_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16743_ clknet_leaf_48_clk _00187_ net611 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13955_ fifo_bank_register.bank\[1\]\[44\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[44\]
+ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__a22o_1
XFILLER_0_221_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12906_ _07755_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16674_ net456 _00122_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
X_13886_ fifo_bank_register.bank\[7\]\[37\] _02218_ _02227_ fifo_bank_register.bank\[2\]\[37\]
+ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a221o_1
X_18413_ clknet_leaf_16_clk _01843_ net630 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[98\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_159_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15625_ _03739_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _07719_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18344_ clknet_leaf_11_clk _01774_ net623 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ _05103_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__buf_4
XFILLER_0_139_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12768_ fifo_bank_register.bank\[2\]\[48\] _05371_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07683_ sky130_fd_sc_hd__mux2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14507_ fifo_bank_register.bank\[7\]\[105\] _02785_ _02794_ fifo_bank_register.bank\[2\]\[105\]
+ _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18275_ clknet_leaf_3_clk _01706_ net583 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[41\]
+ sky130_fd_sc_hd__dfrtp_4
X_11719_ fifo_bank_register.bank\[6\]\[65\] _05407_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07129_ sky130_fd_sc_hd__mux2_1
X_15487_ _03652_ _04784_ _05560_ _03656_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12699_ _07646_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17226_ net476 _00669_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput10 data_i[108] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__buf_2
X_14438_ _02775_ fifo_bank_register.data_out\[97\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02777_ sky130_fd_sc_hd__mux2_1
Xinput21 data_i[118] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput32 data_i[12] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__buf_4
XFILLER_0_226_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput43 data_i[22] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_2
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput54 data_i[32] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17157_ net523 _00600_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput65 data_i[42] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__buf_4
XFILLER_0_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14369_ _02142_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__clkbuf_4
Xinput76 data_i[52] vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_4
Xinput87 data_i[62] vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_4
Xinput98 data_i[72] vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__clkbuf_4
X_16108_ _05052_ _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_229_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17088_ net493 _00531_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08930_ _04942_ _04945_ _04950_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16039_ net195 ks1.key_reg\[43\] _03910_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08861_ addroundkey_data_o\[48\] mix1.data_o\[48\] _04666_ vssd1 vssd1 vccd1 vccd1
+ _04885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08792_ _04670_ _04814_ _04815_ _04713_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a22o_1
XFILLER_0_224_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09413_ fifo_bank_register.bank\[9\]\[47\] _05369_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09344_ net175 vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__buf_2
XFILLER_0_59_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09275_ net191 vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_173_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08226_ net9 net8 net11 net10 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10050_ net181 ks1.key_reg\[30\] _05825_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__mux2_2
XTAP_5614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_199_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13740_ fifo_bank_register.bank\[9\]\[20\] _02137_ _02145_ _02150_ _02155_ vssd1
+ vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_74_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10952_ mix1.data_o\[118\] _04626_ _05617_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13671_ fifo_bank_register.bank\[7\]\[14\] _08182_ _08191_ fifo_bank_register.bank\[2\]\[14\]
+ _02092_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__a221o_1
X_10883_ _04624_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15410_ _04369_ _04949_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__nor2_2
XFILLER_0_13_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12622_ _07605_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__clkbuf_1
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16390_ ks1.key_reg\[92\] _04272_ _04264_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__mux2_1
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15341_ _03563_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12553_ _07569_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18060_ net523 _01503_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_11504_ _07015_ vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15272_ net752 _03521_ _03498_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ _07533_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17011_ net405 _00454_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14223_ _02585_ fifo_bank_register.data_out\[73\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11435_ fifo_bank_register.bank\[7\]\[59\] _05394_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366_ fifo_bank_register.bank\[7\]\[26\] _05325_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06943_ sky130_fd_sc_hd__mux2_1
X_14154_ fifo_bank_register.bank\[9\]\[66\] _02469_ _02521_ _02522_ _02523_ vssd1
+ vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_162_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ _06120_ _06121_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13105_ _07860_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11297_ _05528_ fifo_bank_register.bank\[8\]\[123\] _06768_ vssd1 vssd1 vccd1 vccd1
+ _06905_ sky130_fd_sc_hd__mux2_1
X_14085_ fifo_bank_register.bank\[5\]\[59\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[59\]
+ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a22o_1
X_10248_ _05949_ _06056_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a21o_1
X_17913_ net575 _01356_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_13036_ _07824_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17844_ net432 _01287_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
X_10179_ _05707_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17775_ net398 _01218_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_191_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14987_ addroundkey_data_o\[90\] _03062_ _03091_ addroundkey_data_o\[58\] vssd1 vssd1
+ vccd1 vccd1 _03261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16726_ clknet_leaf_41_clk _00170_ net658 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13938_ fifo_bank_register.bank\[6\]\[42\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[42\]
+ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16657_ net454 _00105_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
X_13869_ fifo_bank_register.bank\[5\]\[35\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[35\]
+ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15608_ mix1.data_o\[9\] _03424_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16588_ net486 _00036_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18327_ clknet_leaf_11_clk _01757_ net631 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15539_ sub1.data_o\[62\] _05235_ _04884_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ sbox1.ah\[2\] _05071_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__nand2_1
X_18258_ clknet_leaf_47_clk _01689_ net652 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_182_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_170_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17209_ net470 _00652_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18189_ clknet_leaf_24_clk _01620_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09962_ _05799_ _05800_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__xor2_1
XFILLER_0_200_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08913_ addroundkey_data_o\[5\] mix1.data_o\[5\] _04657_ vssd1 vssd1 vccd1 vccd1
+ _04937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09893_ _05712_ _05736_ _05737_ _05716_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__a22o_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ ks1.key_reg\[22\] _04725_ _04867_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_176_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08775_ ks1.key_reg\[3\] _04730_ _04732_ net191 vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__o31a_1
XFILLER_0_174_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09327_ net170 vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_193_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ fifo_bank_register.read_ptr\[2\] vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__buf_2
XFILLER_0_209_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08209_ _04368_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09189_ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11220_ _05451_ fifo_bank_register.bank\[8\]\[86\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11151_ _05382_ fifo_bank_register.bank\[8\]\[53\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06829_ sky130_fd_sc_hd__mux2_1
XTAP_6101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10102_ _05913_ _05754_ sub1.data_o\[35\] _05902_ vssd1 vssd1 vccd1 vccd1 _05926_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _05311_ fifo_bank_register.bank\[8\]\[20\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput200 key_i[48] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_4
XTAP_5411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput211 key_i[58] vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_4
XTAP_5433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910_ addroundkey_data_o\[23\] _04375_ _04900_ _03184_ vssd1 vssd1 vccd1 vccd1
+ _03185_ sky130_fd_sc_hd__a211o_1
X_10033_ _05862_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__xor2_1
Xinput222 key_i[68] vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__buf_4
XTAP_5444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput233 key_i[78] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_4
XTAP_5455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15890_ _03879_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__clkbuf_1
Xinput244 key_i[88] vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__buf_4
XTAP_4721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput255 key_i[98] vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__buf_4
XTAP_5466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _03099_ _03116_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_76_1136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ net538 _01003_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14772_ ks1.col\[22\] _05235_ _00007_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__mux2_1
X_11984_ fifo_bank_register.bank\[5\]\[62\] _05401_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16511_ _04339_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__clkbuf_1
X_13723_ _02138_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10935_ addroundkey_data_o\[116\] _06677_ _06612_ vssd1 vssd1 vccd1 vccd1 _06678_
+ sky130_fd_sc_hd__mux2_1
X_17491_ net507 _00934_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16442_ _04301_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__clkbuf_1
X_13654_ fifo_bank_register.bank\[5\]\[12\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10866_ sub1.data_o\[110\] _06614_ _06573_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12605_ _07596_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__clkbuf_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _04262_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__clkbuf_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _08151_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10797_ _06553_ vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__clkbuf_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18112_ net454 _01555_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[114\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _03554_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__clkbuf_1
X_12536_ _07560_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_998 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18043_ net406 _01486_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[45\]
+ sky130_fd_sc_hd__dfxtp_1
X_15255_ _03508_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ _07524_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14206_ fifo_bank_register.bank\[0\]\[71\] _02570_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11418_ _06970_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__clkbuf_1
X_15186_ _03421_ _03449_ _05198_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12398_ fifo_bank_register.bank\[3\]\[1\] _05272_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14137_ fifo_bank_register.bank\[1\]\[64\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[64\]
+ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__a22o_1
X_11349_ _06933_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14068_ fifo_bank_register.bank\[7\]\[57\] _02380_ _02389_ fifo_bank_register.bank\[2\]\[57\]
+ _02446_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__a221o_1
XFILLER_0_207_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13019_ _07815_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17827_ net404 _01270_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08560_ addroundkey_data_o\[118\] fifo_bank_register.data_out\[118\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__mux2_1
X_17758_ net482 _01201_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08491_ addroundkey_data_o\[85\] fifo_bank_register.data_out\[85\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__mux2_1
X_16709_ clknet_leaf_50_clk _00153_ net616 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17689_ net539 _01132_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09112_ _05112_ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09043_ _05010_ _05009_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09945_ _05785_ vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ mix1.data_o\[12\] _05677_ _05703_ _05704_ sub1.data_o\[12\] vssd1 vssd1 vccd1
+ vccd1 _05723_ sky130_fd_sc_hd__a32o_1
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08827_ addroundkey_data_o\[102\] _04778_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__or2_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _04689_ _04780_ _04716_ _04781_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a22o_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_305 net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_327 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08689_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_349 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _04610_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__clkbuf_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10651_ net244 ks1.key_reg\[88\] _06324_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10582_ _06357_ _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__xnor2_1
X_13370_ _08000_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ _07446_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15040_ addroundkey_data_o\[123\] _03057_ _03312_ vssd1 vssd1 vccd1 vccd1 _03313_
+ sky130_fd_sc_hd__a21oi_2
X_12252_ _07410_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11203_ _05434_ fifo_bank_register.bank\[8\]\[78\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06856_ sky130_fd_sc_hd__mux2_1
X_12183_ _05329_ fifo_bank_register.bank\[4\]\[28\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11134_ _05365_ fifo_bank_register.bank\[8\]\[45\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06820_ sky130_fd_sc_hd__mux2_1
X_16991_ net508 _00434_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_11065_ _06783_ vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__clkbuf_1
X_15942_ net254 ks1.key_reg\[97\] _03902_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__mux2_2
XTAP_5230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ net176 ks1.key_reg\[26\] _05825_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__mux2_2
XTAP_5274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15873_ sub1.data_o\[91\] _05195_ _04888_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__mux2_1
XTAP_5285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14824_ _04375_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__buf_4
XTAP_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17612_ net479 _01055_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18592_ clknet_leaf_77_clk _02021_ net589 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[119\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17543_ net521 _00986_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _03041_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__clkbuf_1
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ fifo_bank_register.bank\[5\]\[54\] _05384_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13706_ fifo_bank_register.bank\[1\]\[18\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__a22o_1
X_10918_ _05574_ _06660_ _06661_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__a21o_1
X_17474_ net495 _00917_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14686_ fifo_bank_register.bank\[5\]\[126\] _08096_ _08099_ fifo_bank_register.bank\[3\]\[126\]
+ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11898_ fifo_bank_register.bank\[5\]\[21\] _05315_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16425_ _04292_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__clkbuf_1
X_13637_ fifo_bank_register.bank\[6\]\[10\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__a22o_1
XFILLER_0_229_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10849_ sub1.data_o\[108\] _06599_ _06573_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16356_ ks1.key_reg\[77\] _04023_ _04252_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13568_ _08136_ fifo_bank_register.data_out\[2\] _08064_ vssd1 vssd1 vccd1 vccd1
+ _08137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15307_ _03545_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12519_ _07551_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__clkbuf_1
X_16287_ _04024_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13499_ fifo_bank_register.read_ptr\[3\] _08074_ vssd1 vssd1 vccd1 vccd1 _08076_
+ sky130_fd_sc_hd__nor2b_1
XFILLER_0_180_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18026_ net485 _01469_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_15238_ _03314_ _03453_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__xor2_2
XFILLER_0_152_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15169_ _03431_ _03434_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09730_ round\[1\] _04613_ round\[2\] vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09661_ _05537_ vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08612_ addroundkey_start_i ks1.ready_o vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_222_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ net136 vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__buf_2
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08543_ _04590_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08474_ addroundkey_data_o\[77\] fifo_bank_register.data_out\[77\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ ks1.key_reg\[10\] _04735_ _05047_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09928_ mix1.data_o\[17\] _05576_ _05758_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__o21a_1
XFILLER_0_204_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09859_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__buf_4
XFILLER_0_226_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12870_ _07736_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__clkbuf_1
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_102 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_113 mix1.data_o\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ _07182_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__clkbuf_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 mix1.data_o\[24\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_157 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_212_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ fifo_bank_register.bank\[5\]\[109\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[109\]
+ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__a22o_1
XANTENNA_168 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ _07146_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__clkbuf_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ addroundkey_data_o\[94\] _06467_ _06431_ vssd1 vssd1 vccd1 vccd1 _06468_
+ sky130_fd_sc_hd__mux2_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ fifo_bank_register.bank\[0\]\[100\] _02805_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11683_ fifo_bank_register.bank\[6\]\[48\] _05371_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07110_ sky130_fd_sc_hd__mux2_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16210_ net212 ks1.key_reg\[59\] _03907_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13422_ _05483_ fifo_bank_register.bank\[0\]\[101\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08028_ sky130_fd_sc_hd__mux2_1
X_10634_ net114 mix1.data_o\[87\] _06111_ vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__mux2_1
X_17190_ net448 _00633_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16141_ _04092_ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__xor2_2
X_13353_ _07991_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__clkbuf_1
X_10565_ _06090_ _06342_ sub1.data_o\[81\] _06079_ vssd1 vssd1 vccd1 vccd1 _06343_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _07437_ vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16072_ _04862_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13284_ _07955_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__clkbuf_1
X_10496_ sub1.data_o\[74\] _06280_ _06239_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15023_ addroundkey_data_o\[115\] _03079_ _03295_ vssd1 vssd1 vccd1 vccd1 _03296_
+ sky130_fd_sc_hd__a21oi_2
X_12235_ _07401_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12166_ _07364_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__buf_4
X_11117_ _05348_ fifo_bank_register.bank\[8\]\[37\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06811_ sky130_fd_sc_hd__mux2_1
X_16974_ net480 _00417_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
X_12097_ fifo_bank_register.bank\[5\]\[116\] _05514_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15925_ _03717_ _04943_ _05245_ _03900_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a31o_1
X_11048_ _06774_ vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 data_i[106] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_4
XTAP_5082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ _03860_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__clkbuf_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14807_ sub1.data_o\[120\] _03079_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_204_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15787_ mix1.data_o\[94\] net716 _03819_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__mux2_1
X_18575_ clknet_leaf_75_clk _02004_ net587 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ fifo_bank_register.bank\[1\]\[29\] _05331_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07805_ sky130_fd_sc_hd__mux2_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_157_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17526_ net392 _00969_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_14738_ ks1.col\[5\] _05225_ _04916_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17457_ net451 _00900_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14669_ _02981_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16408_ net799 _03934_ _04281_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__mux2_1
X_17388_ net428 _00831_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16339_ net823 _03953_ _04240_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput301 net301 vssd1 vssd1 vccd1 vccd1 data_o[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput312 net312 vssd1 vssd1 vccd1 vccd1 data_o[31] sky130_fd_sc_hd__buf_2
XFILLER_0_207_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_199_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput323 net323 vssd1 vssd1 vccd1 vccd1 data_o[41] sky130_fd_sc_hd__clkbuf_4
X_18009_ net535 _01452_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput334 net334 vssd1 vssd1 vccd1 vccd1 data_o[51] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput345 net345 vssd1 vssd1 vccd1 vccd1 data_o[61] sky130_fd_sc_hd__buf_2
XFILLER_0_11_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput356 net356 vssd1 vssd1 vccd1 vccd1 data_o[71] sky130_fd_sc_hd__clkbuf_4
Xoutput367 net367 vssd1 vssd1 vccd1 vccd1 data_o[81] sky130_fd_sc_hd__buf_2
XFILLER_0_199_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput378 net378 vssd1 vssd1 vccd1 vccd1 data_o[91] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09713_ _05574_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09644_ net155 vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_184_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09575_ _05479_ vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08526_ _04581_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08457_ _04478_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__buf_8
XFILLER_0_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08388_ addroundkey_data_o\[36\] fifo_bank_register.data_out\[36\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__mux2_2
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10350_ net82 mix1.data_o\[58\] _05989_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09009_ mix1.data_o\[42\] _04692_ _04694_ mix1.data_o\[34\] vssd1 vssd1 vccd1 vccd1
+ _05031_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10281_ net76 mix1.data_o\[52\] _05934_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12020_ _07287_ vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout550 net551 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__clkbuf_2
Xfanout561 net564 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout572 net576 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__buf_2
Xfanout583 net584 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_4
X_13971_ fifo_bank_register.bank\[1\]\[46\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[46\]
+ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout594 net595 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__clkbuf_2
X_15710_ _03784_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__clkbuf_1
X_12922_ _07763_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16690_ clknet_leaf_54_clk _00137_ net616 vssd1 vssd1 vccd1 vccd1 addroundkey_round\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15641_ _03748_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12853_ _07727_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__clkbuf_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18360_ clknet_leaf_1_clk _01790_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[45\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _07173_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__clkbuf_1
X_15572_ _03700_ _03709_ _05548_ _03711_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__a31o_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _07691_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ net536 _00754_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ fifo_bank_register.bank\[7\]\[107\] _02785_ _02794_ fifo_bank_register.bank\[2\]\[107\]
+ _02851_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a221o_1
X_18291_ clknet_leaf_71_clk _01722_ net652 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[57\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _07137_ vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17242_ net487 _00685_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14454_ fifo_bank_register.bank\[0\]\[99\] _02790_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11666_ _07078_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__buf_4
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13405_ _05466_ fifo_bank_register.bank\[0\]\[93\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10617_ _06389_ _06390_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__xnor2_1
X_17173_ net553 _00616_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14385_ fifo_bank_register.bank\[6\]\[91\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[91\]
+ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11597_ _07064_ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16124_ net205 ks1.key_reg\[52\] _03937_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13336_ _05396_ fifo_bank_register.bank\[0\]\[60\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07983_ sky130_fd_sc_hd__mux2_1
X_10548_ addroundkey_data_o\[79\] _06326_ _06327_ vssd1 vssd1 vccd1 vccd1 _06328_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16055_ ks1.key_reg\[12\] _04017_ _03958_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__mux2_1
X_13267_ _07946_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__clkbuf_1
X_10479_ net98 mix1.data_o\[72\] _06237_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15006_ _03276_ _03279_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__nor2_8
X_12218_ _07392_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13198_ fifo_bank_register.bank\[1\]\[124\] _05530_ _07771_ vssd1 vssd1 vccd1 vccd1
+ _07909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12149_ _05295_ fifo_bank_register.bank\[4\]\[12\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16957_ net469 _00400_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15908_ _03891_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16888_ net558 _00331_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_177_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18627_ clknet_leaf_23_clk _02056_ net645 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_188_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15839_ mix1.data_o\[119\] net790 _03729_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09360_ _05312_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__buf_4
XFILLER_0_133_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18558_ clknet_leaf_65_clk _01987_ net589 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[85\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08311_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__buf_12
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17509_ net424 _00952_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09291_ fifo_bank_register.bank\[9\]\[8\] _05286_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18489_ clknet_leaf_59_clk _01918_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_13 _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ net48 net47 net50 net49 vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__or4_1
XANTENNA_24 _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 _05043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 _06336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_57 addroundkey_data_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_68 addroundkey_data_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_79 addroundkey_data_o\[67\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ fifo_bank_register.bank\[9\]\[116\] _05514_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09558_ net251 vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_211_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08509_ _04572_ vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09489_ _05421_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11520_ _07023_ vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ _06987_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10402_ net217 ks1.key_reg\[63\] _06166_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__mux2_2
X_14170_ fifo_bank_register.bank\[1\]\[68\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[68\]
+ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__a22o_1
X_11382_ _06951_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ fifo_bank_register.bank\[1\]\[87\] _05453_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07869_ sky130_fd_sc_hd__mux2_1
X_10333_ net80 mix1.data_o\[56\] _05989_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13052_ fifo_bank_register.bank\[1\]\[54\] _05384_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07833_ sky130_fd_sc_hd__mux2_1
X_10264_ net203 ks1.key_reg\[50\] _05920_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__mux2_2
X_12003_ fifo_bank_register.bank\[5\]\[71\] _05420_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10195_ sub1.data_o\[43\] _06010_ _05991_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__mux2_1
X_17860_ net531 _01303_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16811_ clknet_leaf_74_clk _00255_ net591 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[102\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_218_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17791_ net550 _01234_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout391 net444 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_219_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16742_ clknet_leaf_47_clk _00186_ net611 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[33\]
+ sky130_fd_sc_hd__dfrtp_4
X_13954_ fifo_bank_register.bank\[6\]\[44\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[44\]
+ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12905_ fifo_bank_register.bank\[2\]\[113\] _05508_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07755_ sky130_fd_sc_hd__mux2_1
X_16673_ net469 _00121_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13885_ fifo_bank_register.bank\[5\]\[37\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[37\]
+ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__a22o_1
XFILLER_0_213_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18412_ clknet_leaf_14_clk _01842_ net630 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[97\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_186_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15624_ mix1.data_o\[17\] _03491_ _03730_ vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__mux2_1
X_12836_ fifo_bank_register.bank\[2\]\[80\] _05438_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07719_ sky130_fd_sc_hd__mux2_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18343_ clknet_leaf_38_clk _01773_ net668 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_189_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15555_ _03668_ _04935_ _05196_ _03699_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__a31o_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _07682_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__clkbuf_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14506_ fifo_bank_register.bank\[5\]\[105\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[105\]
+ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18274_ clknet_leaf_3_clk _01705_ net583 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[40\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11718_ _07128_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__clkbuf_1
X_15486_ sub1.data_o\[106\] _03600_ _03653_ sub1.data_o\[42\] vssd1 vssd1 vccd1 vccd1
+ _03656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12698_ fifo_bank_register.bank\[2\]\[15\] _05301_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17225_ net475 _00668_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14437_ _08063_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__buf_4
XFILLER_0_226_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput11 data_i[109] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_4
X_11649_ _07092_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput22 data_i[119] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_4
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput33 data_i[13] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_2
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput44 data_i[23] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17156_ net523 _00599_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14368_ _02140_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__clkbuf_4
Xinput55 data_i[33] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_4
Xinput66 data_i[43] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_4
Xinput77 data_i[53] vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_4
X_16107_ _04062_ _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__xor2_2
X_13319_ _05380_ fifo_bank_register.bank\[0\]\[52\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07974_ sky130_fd_sc_hd__mux2_1
Xinput88 data_i[63] vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput99 data_i[73] vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__buf_4
X_17087_ net491 _00530_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
X_14299_ _02653_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16038_ net708 ks1.next_ready_o _04001_ _04002_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__o22a_1
XFILLER_0_228_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08860_ _04670_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08791_ addroundkey_data_o\[67\] mix1.data_o\[67\] _04805_ vssd1 vssd1 vccd1 vccd1
+ _04815_ sky130_fd_sc_hd__mux2_1
X_17989_ net443 _01432_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09412_ net199 vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09343_ _05322_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09274_ _05275_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ net31 _04381_ net30 net594 vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__or4b_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08989_ _04872_ _05010_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__nor2_1
XTAP_4925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10951_ _05574_ _06690_ _06691_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13670_ fifo_bank_register.bank\[5\]\[14\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__a22o_1
X_10882_ sub1.data_o\[112\] _06628_ _06478_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ fifo_bank_register.bank\[3\]\[107\] _05495_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ net740 _03505_ _03560_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12552_ fifo_bank_register.bank\[3\]\[74\] _05426_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11503_ fifo_bank_register.bank\[7\]\[91\] _05462_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07015_ sky130_fd_sc_hd__mux2_1
X_15271_ _03431_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_19_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12483_ fifo_bank_register.bank\[3\]\[41\] _05357_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17010_ net392 _00453_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14222_ fifo_bank_register.bank\[0\]\[73\] _02584_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02585_ sky130_fd_sc_hd__mux2_1
X_11434_ _06978_ vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14153_ fifo_bank_register.bank\[1\]\[66\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[66\]
+ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11365_ _06942_ vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13104_ fifo_bank_register.bank\[1\]\[79\] _05436_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07860_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10316_ net207 ks1.key_reg\[54\] _06097_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__mux2_1
X_14084_ _08181_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11296_ _06904_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13035_ fifo_bank_register.bank\[1\]\[46\] _05367_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07824_ sky130_fd_sc_hd__mux2_1
X_17912_ net557 _01355_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
X_10247_ _05913_ _05972_ sub1.data_o\[49\] _05902_ vssd1 vssd1 vccd1 vccd1 _06057_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17843_ net458 _01286_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
X_10178_ _05829_ _05992_ _05995_ _05833_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17774_ net395 _01217_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14986_ sub1.data_o\[122\] _03077_ _03259_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_191_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16725_ clknet_leaf_41_clk _00169_ net658 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_159_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13937_ fifo_bank_register.bank\[7\]\[42\] _02299_ _02308_ fifo_bank_register.bank\[2\]\[42\]
+ _02330_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a221o_1
XFILLER_0_187_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13868_ _02269_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__clkbuf_1
X_16656_ net403 _00104_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_201_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15607_ _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__clkbuf_4
X_12819_ fifo_bank_register.bank\[2\]\[72\] _05422_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16587_ net486 _00035_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_13799_ fifo_bank_register.bank\[0\]\[27\] _02207_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18326_ clknet_leaf_11_clk _01756_ net631 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15538_ _03688_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__clkbuf_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18257_ clknet_leaf_21_clk _01688_ net646 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_15469_ sub1.data_o\[36\] _03644_ _03636_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17208_ net456 _00651_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18188_ clknet_leaf_18_clk _01619_ net638 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[82\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17139_ net406 _00582_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ net170 ks1.key_reg\[20\] _05708_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08912_ addroundkey_data_o\[61\] mix1.data_o\[61\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09892_ mix1.data_o\[14\] _05677_ _05703_ _05704_ sub1.data_o\[14\] vssd1 vssd1 vccd1
+ vccd1 _05737_ sky130_fd_sc_hd__a32o_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ ks1.key_reg\[22\] _04729_ _04731_ net172 vssd1 vssd1 vccd1 vccd1 _04867_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_97_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_225_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08774_ ks1.key_reg\[11\] _04735_ _04797_ net152 vssd1 vssd1 vccd1 vccd1 _04798_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_224_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09326_ _05310_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09257_ fifo_bank_register.read_ptr\[1\] _05260_ vssd1 vssd1 vccd1 vccd1 _05261_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08208_ _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09188_ _05198_ _04367_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__nor2_1
XFILLER_0_181_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11150_ _06828_ vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__clkbuf_1
XTAP_6102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10101_ sub1.data_o\[35\] _05924_ _05751_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__mux2_1
XTAP_6124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11081_ _06791_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__buf_4
XTAP_5401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput201 key_i[49] vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_8
XTAP_5412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput212 key_i[59] vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_4
X_10032_ net178 ks1.key_reg\[28\] _05825_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__mux2_2
XTAP_5434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput223 key_i[69] vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_4
XTAP_5445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput234 key_i[79] vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput245 key_i[89] vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__buf_4
Xinput256 key_i[99] vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__buf_4
XTAP_5467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14840_ _03107_ _03115_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__xor2_2
XTAP_5489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ _03049_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_216_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11983_ _07268_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__clkbuf_1
XTAP_4799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16510_ net771 _03487_ _04332_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__mux2_1
X_13722_ _08091_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__buf_6
X_10934_ _06675_ _06676_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_169_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17490_ net500 _00933_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13653_ _02077_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__clkbuf_1
X_16441_ net793 _04068_ _04295_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10865_ net13 mix1.data_o\[110\] _06571_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12604_ fifo_bank_register.bank\[3\]\[99\] _05478_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07596_ sky130_fd_sc_hd__mux2_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16372_ net800 _04086_ _04252_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13584_ _08150_ fifo_bank_register.data_out\[4\] _08064_ vssd1 vssd1 vccd1 vccd1
+ _08151_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10796_ addroundkey_data_o\[102\] _06552_ _06522_ vssd1 vssd1 vccd1 vccd1 _06553_
+ sky130_fd_sc_hd__mux2_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ net718 _03467_ _03549_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__mux2_1
X_18111_ net470 _01554_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12535_ fifo_bank_register.bank\[3\]\[66\] _05409_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_227_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15254_ net792 _03507_ _03498_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18042_ net389 _01485_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ fifo_bank_register.bank\[3\]\[33\] _05340_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14205_ fifo_bank_register.bank\[9\]\[71\] _02550_ _02567_ _02568_ _02569_ vssd1
+ vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_227_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11417_ fifo_bank_register.bank\[7\]\[50\] _05375_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06970_ sky130_fd_sc_hd__mux2_1
X_15185_ _03281_ _03448_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_160_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12397_ _07487_ vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14136_ fifo_bank_register.bank\[6\]\[64\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[64\]
+ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11348_ fifo_bank_register.bank\[7\]\[18\] _05307_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14067_ fifo_bank_register.bank\[5\]\[57\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[57\]
+ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a22o_1
X_11279_ _05510_ fifo_bank_register.bank\[8\]\[114\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13018_ fifo_bank_register.bank\[1\]\[38\] _05350_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17826_ net410 _01269_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17757_ net483 _01200_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14969_ addroundkey_data_o\[15\] _04376_ _05606_ _03242_ vssd1 vssd1 vccd1 vccd1
+ _03243_ sky130_fd_sc_hd__a211o_1
XFILLER_0_222_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16708_ clknet_leaf_44_clk next_addroundkey_start_i net658 vssd1 vssd1 vccd1 vccd1
+ addroundkey_start_i sky130_fd_sc_hd__dfrtp_4
XFILLER_0_159_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08490_ _04562_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17688_ net539 _01131_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16639_ net555 _00087_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_169_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09111_ _05120_ _05121_ sbox1.alph\[3\] vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18309_ clknet_leaf_2_clk _01740_ net624 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[75\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09042_ _05010_ _05009_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09944_ addroundkey_data_o\[18\] _05784_ _05697_ vssd1 vssd1 vccd1 vccd1 _05785_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09875_ sub1.data_o\[12\] _05721_ _05701_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__mux2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _04848_ _04849_ _04650_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__mux2_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08757_ addroundkey_data_o\[89\] mix1.data_o\[89\] _04662_ vssd1 vssd1 vccd1 vccd1
+ _04781_ sky130_fd_sc_hd__mux2_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_306 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_317 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_328 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08688_ sub1.state\[3\] sub1.state\[2\] _04687_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__and3b_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10650_ _06416_ _06418_ _06419_ _06420_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09309_ net163 vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__buf_2
XFILLER_0_180_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10581_ net238 ks1.key_reg\[82\] _06097_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__mux2_4
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _05466_ fifo_bank_register.bank\[4\]\[93\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12251_ _05396_ fifo_bank_register.bank\[4\]\[60\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11202_ _06855_ vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__clkbuf_1
X_12182_ _07373_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11133_ _06819_ vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16990_ net482 _00433_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11064_ _05295_ fifo_bank_register.bank\[8\]\[12\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06783_ sky130_fd_sc_hd__mux2_1
X_15941_ net704 _03901_ _03913_ _03915_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__a22o_1
XTAP_5231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10015_ _05829_ _05846_ _05847_ _05833_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__a22o_1
XTAP_5264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15872_ _03868_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__clkbuf_1
XTAP_5286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17611_ net476 _01054_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_162_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14823_ _03095_ _03098_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__nor2_8
XTAP_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18591_ clknet_leaf_75_clk _02020_ net587 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ net512 _00985_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14754_ ks1.col\[29\] _05225_ _04911_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11966_ _07259_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__clkbuf_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10917_ _06630_ _06514_ sub1.data_o\[115\] _05675_ vssd1 vssd1 vccd1 vccd1 _06661_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ fifo_bank_register.bank\[6\]\[18\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__a22o_1
X_17473_ net439 _00916_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
X_14685_ _02995_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11897_ _07223_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13636_ _08107_ vssd1 vssd1 vccd1 vccd1 _08197_ sky130_fd_sc_hd__clkbuf_4
X_16424_ net797 _04006_ _04281_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__mux2_1
X_10848_ net10 mix1.data_o\[108\] _06571_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13567_ fifo_bank_register.bank\[0\]\[2\] _08135_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08136_ sky130_fd_sc_hd__mux2_1
X_16355_ _04253_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__clkbuf_1
X_10779_ _06491_ _06535_ _06536_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15306_ net789 _03382_ _03539_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__mux2_1
X_12518_ fifo_bank_register.bank\[3\]\[58\] _05392_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07551_ sky130_fd_sc_hd__mux2_1
X_16286_ _04215_ _04016_ _04216_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13498_ _08067_ _08074_ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18025_ net426 _01468_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[27\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_112_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15237_ _03494_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12449_ fifo_bank_register.bank\[3\]\[25\] _05323_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15168_ _03432_ _03433_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14119_ fifo_bank_register.bank\[7\]\[62\] _02461_ _02470_ fifo_bank_register.bank\[2\]\[62\]
+ _02492_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15099_ addroundkey_data_o\[100\] _03143_ _03369_ vssd1 vssd1 vccd1 vccd1 _03370_
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_157_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09660_ fifo_bank_register.bank\[9\]\[127\] _05536_ _05269_ vssd1 vssd1 vccd1 vccd1
+ _05537_ sky130_fd_sc_hd__mux2_1
X_08611_ _04632_ _04633_ _04634_ _04635_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__or4_2
X_17809_ net552 _01252_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09591_ _05490_ vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_206_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ addroundkey_data_o\[109\] fifo_bank_register.data_out\[109\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__mux2_2
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08473_ _04553_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_198_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09025_ ks1.key_reg\[10\] _04745_ _04746_ net141 vssd1 vssd1 vccd1 vccd1 _05047_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_182_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09927_ _05575_ _05767_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a21o_1
XFILLER_0_217_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09858_ _04638_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _04741_ _04796_ _04801_ _04832_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__o211a_1
XFILLER_0_198_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09789_ net62 mix1.data_o\[3\] _05604_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__mux2_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11820_ fifo_bank_register.bank\[6\]\[113\] _05508_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07182_ sky130_fd_sc_hd__mux2_1
XANTENNA_103 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_114 mix1.data_o\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 mix1.data_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_136 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ fifo_bank_register.bank\[6\]\[80\] _05438_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07146_ sky130_fd_sc_hd__mux2_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_169 net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _06465_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__xor2_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _02157_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11682_ _07109_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13421_ _08027_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__clkbuf_1
X_10633_ _06405_ vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16140_ net242 ks1.key_reg\[86\] _03906_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13352_ _05413_ fifo_bank_register.bank\[0\]\[68\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ sub1.ready_o vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12303_ _05449_ fifo_bank_register.bank\[4\]\[85\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16071_ _04030_ _04031_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__xor2_4
XFILLER_0_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13283_ _05344_ fifo_bank_register.bank\[0\]\[35\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07955_ sky130_fd_sc_hd__mux2_1
X_10495_ net100 mix1.data_o\[74\] _06237_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15022_ addroundkey_data_o\[19\] _03208_ _03086_ _03294_ vssd1 vssd1 vccd1 vccd1
+ _03295_ sky130_fd_sc_hd__a211o_1
X_12234_ _05380_ fifo_bank_register.bank\[4\]\[52\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12165_ _07340_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__buf_6
X_11116_ _06810_ vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16973_ net479 _00416_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12096_ _07327_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__clkbuf_1
XTAP_5050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15924_ sub1.data_o\[47\] _03576_ _03892_ sub1.data_o\[111\] vssd1 vssd1 vccd1 vccd1
+ _03900_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11047_ _05278_ fifo_bank_register.bank\[8\]\[4\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06774_ sky130_fd_sc_hd__mux2_1
XTAP_5061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput9 data_i[107] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_4
XTAP_5083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ mix1.data_o\[127\] net706 _03729_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__mux2_1
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ sub1.data_o\[88\] _03072_ _03080_ _03081_ vssd1 vssd1 vccd1 vccd1 _03082_
+ sky130_fd_sc_hd__a211o_1
X_18574_ clknet_leaf_81_clk _02003_ net578 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15786_ _03824_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__clkbuf_1
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _07804_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__clkbuf_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ net394 _00968_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_14737_ _03032_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__clkbuf_1
X_11949_ _07250_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17456_ net465 _00899_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
X_14668_ _02980_ fifo_bank_register.data_out\[123\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _02981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16407_ _04283_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13619_ _08076_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__buf_6
XFILLER_0_166_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17387_ net417 _00830_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14599_ fifo_bank_register.bank\[6\]\[115\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[115\]
+ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16338_ _04244_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16269_ _04207_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput302 net302 vssd1 vssd1 vccd1 vccd1 data_o[22] sky130_fd_sc_hd__buf_2
X_18008_ net493 _01451_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[10\]
+ sky130_fd_sc_hd__dfxtp_1
Xoutput313 net313 vssd1 vssd1 vccd1 vccd1 data_o[32] sky130_fd_sc_hd__clkbuf_4
Xoutput324 net324 vssd1 vssd1 vccd1 vccd1 data_o[42] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput335 net335 vssd1 vssd1 vccd1 vccd1 data_o[52] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput346 net346 vssd1 vssd1 vccd1 vccd1 data_o[62] sky130_fd_sc_hd__buf_2
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput357 net357 vssd1 vssd1 vccd1 vccd1 data_o[72] sky130_fd_sc_hd__buf_2
Xoutput368 net368 vssd1 vssd1 vccd1 vccd1 data_o[82] sky130_fd_sc_hd__buf_2
XFILLER_0_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput379 net379 vssd1 vssd1 vccd1 vccd1 data_o[92] sky130_fd_sc_hd__buf_2
XFILLER_0_199_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09712_ _04625_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_208_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09643_ _05525_ vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09574_ fifo_bank_register.bank\[9\]\[99\] _05478_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08525_ addroundkey_data_o\[101\] fifo_bank_register.data_out\[101\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_62_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08456_ _04544_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08387_ _04508_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09008_ _05020_ _05023_ _05026_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__or4_1
X_10280_ _06087_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout540 net542 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__clkbuf_2
Xfanout551 net577 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__buf_2
Xfanout562 net564 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_2
XFILLER_0_217_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13970_ fifo_bank_register.bank\[6\]\[46\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[46\]
+ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a22o_1
Xfanout573 net576 vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__clkbuf_2
Xfanout584 net585 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
Xfanout595 net596 vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__clkbuf_4
X_12921_ fifo_bank_register.bank\[2\]\[121\] _05524_ _07628_ vssd1 vssd1 vccd1 vccd1
+ _07763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ mix1.data_o\[24\] _03514_ _03742_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ fifo_bank_register.bank\[2\]\[88\] _05455_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07727_ sky130_fd_sc_hd__mux2_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ fifo_bank_register.bank\[6\]\[105\] _05491_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07173_ sky130_fd_sc_hd__mux2_1
X_15571_ sub1.data_o\[8\] _03660_ _03710_ sub1.data_o\[72\] vssd1 vssd1 vccd1 vccd1
+ _03711_ sky130_fd_sc_hd__a22o_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ fifo_bank_register.bank\[2\]\[55\] _05386_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_clk clknet_3_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17310_ net541 _00753_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ fifo_bank_register.bank\[6\]\[72\] _05422_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07137_ sky130_fd_sc_hd__mux2_1
X_14522_ fifo_bank_register.bank\[5\]\[107\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[107\]
+ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a22o_1
X_18290_ clknet_leaf_46_clk _01721_ net652 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[56\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17241_ net502 _00684_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11665_ _07100_ vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__clkbuf_1
X_14453_ fifo_bank_register.bank\[9\]\[99\] _02712_ _02787_ _02788_ _02789_ vssd1
+ vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_86_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13404_ _08018_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__clkbuf_1
X_10616_ net241 ks1.key_reg\[85\] _06097_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__mux2_4
XFILLER_0_148_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14384_ fifo_bank_register.bank\[7\]\[91\] _02704_ _02713_ fifo_bank_register.bank\[2\]\[91\]
+ _02728_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a221o_1
X_17172_ net525 _00615_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11596_ fifo_bank_register.bank\[6\]\[7\] _05284_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13335_ _07937_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16123_ _04076_ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__xor2_4
X_10547_ _05792_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__buf_6
XFILLER_0_84_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13266_ _05327_ fifo_bank_register.bank\[0\]\[27\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16054_ _04736_ _04016_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_161_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10478_ _06265_ vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15005_ addroundkey_data_o\[97\] _03056_ _03278_ vssd1 vssd1 vccd1 vccd1 _03279_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12217_ _05363_ fifo_bank_register.bank\[4\]\[44\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13197_ _07908_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12148_ _07355_ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16956_ net457 _00399_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
X_12079_ _07318_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15907_ sub1.data_o\[103\] _03890_ _03876_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16887_ net405 _00330_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_18626_ clknet_leaf_24_clk _02055_ net645 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[119\]
+ sky130_fd_sc_hd__dfrtp_1
X_15838_ _03851_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18557_ clknet_leaf_78_clk _01986_ net589 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[84\]
+ sky130_fd_sc_hd__dfrtp_1
X_15769_ _03815_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08310_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__buf_8
X_17508_ net418 _00951_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09290_ net246 vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__clkbuf_4
X_18488_ clknet_leaf_56_clk _01917_ net614 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _04394_ _04395_ _04396_ _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__or4_1
XFILLER_0_145_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_14 _04487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ net548 _00882_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_25 _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_184_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_36 _05244_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 _06348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_58 addroundkey_data_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_69 addroundkey_data_o\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09626_ net148 vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__buf_2
XFILLER_0_223_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09557_ _05467_ vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08508_ addroundkey_data_o\[93\] fifo_bank_register.data_out\[93\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__mux2_4
XFILLER_0_210_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09488_ fifo_bank_register.bank\[9\]\[71\] _05420_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08439_ addroundkey_data_o\[60\] fifo_bank_register.data_out\[60\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ fifo_bank_register.bank\[7\]\[66\] _05409_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ _06171_ _06195_ _06196_ _06175_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11381_ fifo_bank_register.bank\[7\]\[33\] _05340_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _07868_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__clkbuf_1
X_10332_ _06135_ vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13051_ _07832_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__clkbuf_1
X_10263_ _05899_ _06067_ _06071_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12002_ _07278_ vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10194_ net66 mix1.data_o\[43\] _05989_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16810_ clknet_leaf_81_clk _00254_ net586 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[101\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_205_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17790_ net571 _01233_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16741_ clknet_leaf_47_clk _00185_ net651 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[32\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout392 net397 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_2
XFILLER_0_219_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13953_ fifo_bank_register.bank\[7\]\[44\] _02299_ _02308_ fifo_bank_register.bank\[2\]\[44\]
+ _02344_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a221o_1
XFILLER_0_221_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12904_ _07754_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16672_ net433 _00120_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ _02283_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__clkbuf_1
X_18411_ clknet_leaf_13_clk _01841_ net628 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[96\]
+ sky130_fd_sc_hd__dfrtp_4
X_15623_ _03738_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__clkbuf_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _07651_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_186_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18342_ clknet_leaf_38_clk _01772_ net668 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15554_ sub1.data_o\[67\] _03691_ _03698_ _03673_ vssd1 vssd1 vccd1 vccd1 _03699_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ fifo_bank_register.bank\[2\]\[47\] _05369_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14505_ _02836_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18273_ clknet_leaf_34_clk _01704_ net662 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ fifo_bank_register.bank\[6\]\[64\] _05405_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_189_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15485_ _03652_ _04784_ _05554_ _03655_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__a31o_1
X_12697_ _07645_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17224_ net476 _00667_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11648_ fifo_bank_register.bank\[6\]\[31\] _05336_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14436_ fifo_bank_register.bank\[0\]\[97\] _02774_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02775_ sky130_fd_sc_hd__mux2_1
Xinput12 data_i[10] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__buf_2
XFILLER_0_142_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput23 data_i[11] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput34 data_i[14] vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput45 data_i[24] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__buf_2
XFILLER_0_123_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17155_ net527 _00598_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11579_ _05249_ _05250_ _06910_ net597 vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__and4b_1
X_14367_ _02138_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__clkbuf_4
Xinput56 data_i[34] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput67 data_i[44] vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_4
Xinput78 data_i[54] vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__buf_4
X_16106_ net203 ks1.key_reg\[50\] _03937_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__mux2_1
X_13318_ _07973_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__clkbuf_1
Xinput89 data_i[64] vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__buf_4
XFILLER_0_204_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14298_ _02652_ fifo_bank_register.data_out\[81\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17086_ net441 _00529_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16037_ _05048_ _04000_ _04371_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13249_ _07936_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08790_ addroundkey_data_o\[51\] mix1.data_o\[51\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _04814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17988_ net531 _01431_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16939_ net450 _00382_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ _05368_ vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__clkbuf_1
X_18609_ clknet_leaf_13_clk _02038_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[102\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_177_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09342_ fifo_bank_register.bank\[9\]\[24\] _05321_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09273_ fifo_bank_register.bank\[9\]\[2\] _05274_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_173_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ net27 net26 net29 net28 vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08988_ _04872_ _05010_ _04649_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__a21o_1
XTAP_4926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10950_ _06630_ sub1.ready_o sub1.data_o\[118\] _05675_ vssd1 vssd1 vccd1 vccd1 _06691_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ fifo_bank_register.bank\[9\]\[110\] _05501_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10881_ net15 mix1.data_o\[112\] _06476_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12620_ _07604_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12551_ _07568_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__clkbuf_1
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11502_ _07014_ vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15270_ _03442_ _03519_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__xnor2_2
X_12482_ _07532_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14221_ fifo_bank_register.bank\[9\]\[73\] _02550_ _02581_ _02582_ _02583_ vssd1
+ vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a2111o_1
X_11433_ fifo_bank_register.bank\[7\]\[58\] _05392_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14152_ fifo_bank_register.bank\[6\]\[66\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[66\]
+ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11364_ fifo_bank_register.bank\[7\]\[25\] _05323_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10315_ _06076_ _06114_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_123_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13103_ _07859_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14083_ _02460_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__clkbuf_1
X_11295_ _05526_ fifo_bank_register.bank\[8\]\[122\] _06768_ vssd1 vssd1 vccd1 vccd1
+ _06904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13034_ _07823_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__clkbuf_1
X_17911_ net408 _01354_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
X_10246_ sub1.data_o\[49\] _06055_ _05936_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17842_ net453 _01285_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10177_ mix1.data_o\[41\] _05876_ _05993_ _05994_ sub1.data_o\[41\] vssd1 vssd1 vccd1
+ vccd1 _05995_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17773_ net415 _01216_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_14985_ sub1.data_o\[26\] _04375_ _04658_ _03258_ vssd1 vssd1 vccd1 vccd1 _03259_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_57_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16724_ clknet_leaf_42_clk _00168_ net659 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13936_ fifo_bank_register.bank\[5\]\[42\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[42\]
+ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_199_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16655_ net402 _00103_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13867_ _02268_ fifo_bank_register.data_out\[34\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15606_ _04379_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__buf_6
XFILLER_0_215_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12818_ _07709_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__clkbuf_1
X_16586_ net510 _00034_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ fifo_bank_register.bank\[9\]\[27\] _02137_ _02204_ _02205_ _02206_ vssd1
+ vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_56_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18325_ clknet_leaf_11_clk _01755_ net628 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_210_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15537_ sub1.data_o\[61\] _05227_ _04884_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__mux2_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ fifo_bank_register.bank\[2\]\[39\] _05352_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18256_ clknet_leaf_22_clk _01687_ net646 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15468_ sub1.data_o\[68\] _05218_ _03633_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17207_ net469 _00650_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14419_ fifo_bank_register.bank\[9\]\[95\] _02712_ _02757_ _02758_ _02759_ vssd1
+ vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__a2111o_1
X_18187_ clknet_leaf_18_clk _01618_ net638 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_181_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15399_ _03019_ _03593_ _05196_ _03599_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17138_ net389 _00581_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09960_ _05712_ _05796_ _05798_ _05716_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17069_ net458 _00512_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08911_ _04684_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__clkbuf_4
X_09891_ sub1.data_o\[14\] _05735_ _05701_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__mux2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _04862_ _04755_ _04863_ _04865_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_176_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08773_ ks1.key_reg\[11\] _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09325_ fifo_bank_register.bank\[9\]\[19\] _05309_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ fifo_bank_register.write_ptr\[3\] _05255_ _05253_ vssd1 vssd1 vccd1 vccd1
+ _05260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08207_ sub1.state\[4\] _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09187_ _04617_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10100_ net57 mix1.data_o\[35\] _05749_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ _06767_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__buf_8
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _05829_ _05860_ _05861_ _05833_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__a22o_1
Xinput202 key_i[4] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_4
XTAP_5424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput213 key_i[5] vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_4
XTAP_5435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput224 key_i[6] vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_4
XTAP_5446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput235 key_i[7] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__buf_4
XTAP_5457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput246 key_i[8] vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__buf_4
XFILLER_0_227_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput257 key_i[9] vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_216_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14770_ ks1.col\[21\] _05225_ _00007_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__mux2_1
XTAP_4789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ fifo_bank_register.bank\[5\]\[61\] _05399_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13721_ _02136_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__buf_4
XFILLER_0_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10933_ net148 ks1.key_reg\[116\] _04639_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__mux2_2
XFILLER_0_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ _04300_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__clkbuf_1
X_10864_ _06613_ vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__clkbuf_1
X_13652_ _02076_ fifo_bank_register.data_out\[11\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _02077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12603_ _07595_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__clkbuf_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16371_ _04261_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ fifo_bank_register.bank\[0\]\[4\] _08149_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08150_ sky130_fd_sc_hd__mux2_1
X_10795_ _06550_ _06551_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__xnor2_1
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18110_ net470 _01553_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _03553_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12534_ _07559_ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18041_ net407 _01484_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[43\]
+ sky130_fd_sc_hd__dfxtp_2
X_15253_ _03117_ _03391_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_163_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12465_ _07523_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_227_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14204_ fifo_bank_register.bank\[1\]\[71\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[71\]
+ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a22o_1
XFILLER_0_223_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11416_ _06935_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__buf_4
X_15184_ _03233_ _03265_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__xor2_1
X_12396_ fifo_bank_register.bank\[3\]\[0\] _05248_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14135_ fifo_bank_register.bank\[7\]\[64\] _02461_ _02470_ fifo_bank_register.bank\[2\]\[64\]
+ _02506_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__a221o_1
X_11347_ _06932_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14066_ _02445_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__clkbuf_1
X_11278_ _06895_ vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10229_ _06001_ _06039_ _06040_ _06005_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13017_ _07814_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17825_ net401 _01268_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1 first_round_reg vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17756_ net501 _01199_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14968_ addroundkey_data_o\[79\] _03108_ _03092_ addroundkey_data_o\[47\] vssd1 vssd1
+ vccd1 vccd1 _03242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16707_ clknet_leaf_44_clk next_addroundkey_ready_o net658 vssd1 vssd1 vccd1 vccd1
+ addroundkey_ready_o sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13919_ fifo_bank_register.bank\[6\]\[40\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[40\]
+ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17687_ net540 _01130_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
X_14899_ sub1.data_o\[30\] _04376_ _03081_ _03173_ vssd1 vssd1 vccd1 vccd1 _03174_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_187_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16638_ net525 _00086_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16569_ net478 _00017_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09110_ _05109_ _05110_ _05118_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__and3_1
X_18308_ clknet_leaf_2_clk _01739_ net624 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[74\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_169_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09041_ _04833_ _05059_ _05060_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__mux2_1
X_18239_ clknet_leaf_32_clk _01670_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ _05782_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09874_ net32 mix1.data_o\[12\] _05699_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__mux2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08825_ addroundkey_data_o\[46\] _04692_ _04694_ addroundkey_data_o\[38\] vssd1 vssd1
+ vccd1 vccd1 _04849_ sky130_fd_sc_hd__a22o_1
XFILLER_0_225_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08756_ addroundkey_data_o\[1\] mix1.data_o\[1\] _04662_ vssd1 vssd1 vccd1 vccd1
+ _04780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_307 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_318 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_329 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _04706_ _04707_ _04708_ _04710_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__a22o_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_166_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09308_ _05298_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__clkbuf_1
X_10580_ _06076_ _06352_ _06356_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ sub1.data_o\[23\] _05200_ _05203_ sub1.data_o\[87\] vssd1 vssd1 vccd1 vccd1
+ _05246_ sky130_fd_sc_hd__a22o_1
XFILLER_0_173_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _07364_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__buf_4
XFILLER_0_224_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11201_ _05432_ fifo_bank_register.bank\[8\]\[77\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06855_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _05327_ fifo_bank_register.bank\[4\]\[27\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11132_ _05363_ fifo_bank_register.bank\[8\]\[44\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ _06782_ vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__clkbuf_1
X_15940_ _04920_ _03912_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__a21oi_1
XTAP_5221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ mix1.data_o\[26\] _05797_ _05821_ _05822_ sub1.data_o\[26\] vssd1 vssd1 vccd1
+ vccd1 _05847_ sky130_fd_sc_hd__a32o_1
XFILLER_0_200_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ sub1.data_o\[90\] _05559_ _04888_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__mux2_1
XTAP_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17610_ net475 _01053_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14822_ addroundkey_data_o\[109\] _03078_ _03097_ vssd1 vssd1 vccd1 vccd1 _03098_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_204_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18590_ clknet_leaf_76_clk _02019_ net588 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ net522 _00984_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _03040_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ fifo_bank_register.bank\[5\]\[53\] _05382_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07259_ sky130_fd_sc_hd__mux2_1
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13704_ fifo_bank_register.bank\[7\]\[18\] _08182_ _08191_ fifo_bank_register.bank\[2\]\[18\]
+ _02121_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__a221o_1
X_10916_ sub1.data_o\[115\] _06659_ _05608_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__mux2_1
X_17472_ net490 _00915_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14684_ _02994_ fifo_bank_register.data_out\[125\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _02995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11896_ fifo_bank_register.bank\[5\]\[20\] _05311_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16423_ _04291_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _08104_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__clkbuf_4
X_10847_ _06598_ vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__clkbuf_1
X_16354_ net796 _04014_ _04252_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ fifo_bank_register.bank\[9\]\[2\] _08090_ _08132_ _08133_ _08134_ vssd1 vssd1
+ vccd1 vccd1 _08135_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10778_ _06395_ _06514_ sub1.data_o\[101\] _06384_ vssd1 vssd1 vccd1 vccd1 _06536_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15305_ _03544_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12517_ _07550_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__clkbuf_1
X_16285_ net679 _04136_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_180_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13497_ fifo_bank_register.read_ptr\[0\] fifo_bank_register.read_ptr\[1\] _05262_
+ vssd1 vssd1 vccd1 vccd1 _08074_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18024_ net510 _01467_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[26\]
+ sky130_fd_sc_hd__dfxtp_1
X_15236_ net748 _03493_ _03425_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12448_ _07514_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15167_ _03273_ _03305_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__xor2_1
XFILLER_0_160_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12379_ _07476_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14118_ fifo_bank_register.bank\[5\]\[62\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[62\]
+ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ addroundkey_data_o\[4\] _04379_ _05607_ _03368_ vssd1 vssd1 vccd1 vccd1 _03369_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14049_ _02430_ fifo_bank_register.data_out\[54\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08610_ round\[2\] addroundkey_round\[2\] vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__xor2_1
X_17808_ net546 _01251_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09590_ fifo_bank_register.bank\[9\]\[104\] _05489_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17739_ net473 _01182_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_08541_ _04466_ vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__buf_8
XFILLER_0_49_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08472_ addroundkey_data_o\[76\] fifo_bank_register.data_out\[76\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09024_ ks1.key_reg\[26\] _04735_ _05045_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09926_ _05201_ _05754_ sub1.data_o\[17\] _05585_ vssd1 vssd1 vccd1 vccd1 _05768_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09857_ _05629_ _05702_ _05705_ _05633_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__a22o_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _04648_ _04830_ _04831_ _04750_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_38_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09788_ _05644_ vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08739_ addroundkey_data_o\[121\] _04658_ _04762_ _04653_ vssd1 vssd1 vccd1 vccd1
+ _04763_ sky130_fd_sc_hd__o211a_1
XANTENNA_104 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_115 mix1.data_o\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 mix1.data_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_148 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11750_ _07078_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__buf_4
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ net251 ks1.key_reg\[94\] _06324_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__mux2_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ fifo_bank_register.bank\[6\]\[47\] _05369_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13420_ _05480_ fifo_bank_register.bank\[0\]\[100\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08027_ sky130_fd_sc_hd__mux2_1
X_10632_ addroundkey_data_o\[86\] _06404_ _06327_ vssd1 vssd1 vccd1 vccd1 _06405_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10563_ _05613_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13351_ _07990_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12302_ _07436_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16070_ net198 ks1.key_reg\[46\] _03910_ vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__mux2_2
XFILLER_0_134_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13282_ _07954_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__clkbuf_1
X_10494_ _06279_ vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__clkbuf_1
X_15021_ addroundkey_data_o\[83\] _03209_ _03084_ addroundkey_data_o\[51\] vssd1 vssd1
+ vccd1 vccd1 _03294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12233_ _07400_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ _07363_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11115_ _05346_ fifo_bank_register.bank\[8\]\[36\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16972_ net479 _00415_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_12095_ fifo_bank_register.bank\[5\]\[115\] _05512_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_194_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15923_ _03717_ _04943_ _05236_ _03899_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__a31o_1
X_11046_ _06773_ vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__clkbuf_1
XTAP_5040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _03859_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__clkbuf_1
XTAP_5095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _03058_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__buf_4
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18573_ clknet_leaf_81_clk _02002_ net578 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[100\]
+ sky130_fd_sc_hd__dfrtp_1
X_15785_ mix1.data_o\[93\] net773 _03819_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__mux2_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12997_ fifo_bank_register.bank\[1\]\[28\] _05329_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17524_ net391 _00967_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ ks1.col\[4\] _05217_ _04916_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__mux2_1
X_11948_ fifo_bank_register.bank\[5\]\[45\] _05365_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ net467 _00898_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14667_ fifo_bank_register.bank\[0\]\[123\] _02979_ _08120_ vssd1 vssd1 vccd1 vccd1
+ _02980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11879_ _07213_ vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16406_ net828 _03926_ _04281_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13618_ _08180_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__clkbuf_1
X_17386_ net422 _00829_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ fifo_bank_register.bank\[7\]\[115\] _02866_ _02875_ fifo_bank_register.bank\[2\]\[115\]
+ _02918_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a221o_1
XFILLER_0_229_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16337_ net847 _03945_ _04240_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13549_ _08119_ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__buf_4
XFILLER_0_125_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_207_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16268_ net825 _03947_ _04206_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18007_ net426 _01450_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15219_ _03466_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__or2_1
XFILLER_0_164_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput303 net303 vssd1 vssd1 vccd1 vccd1 data_o[23] sky130_fd_sc_hd__clkbuf_4
Xoutput314 net314 vssd1 vssd1 vccd1 vccd1 data_o[33] sky130_fd_sc_hd__buf_2
X_16199_ _04146_ _04147_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__xor2_2
Xoutput325 net325 vssd1 vssd1 vccd1 vccd1 data_o[43] sky130_fd_sc_hd__clkbuf_4
Xoutput336 net336 vssd1 vssd1 vccd1 vccd1 data_o[53] sky130_fd_sc_hd__clkbuf_4
Xoutput347 net347 vssd1 vssd1 vccd1 vccd1 data_o[63] sky130_fd_sc_hd__buf_2
Xoutput358 net358 vssd1 vssd1 vccd1 vccd1 data_o[73] sky130_fd_sc_hd__buf_2
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput369 net369 vssd1 vssd1 vccd1 vccd1 data_o[83] sky130_fd_sc_hd__buf_2
XFILLER_0_142_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09711_ _04619_ _05571_ _05572_ _05573_ _04613_ vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__a32o_1
XFILLER_0_208_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09642_ fifo_bank_register.bank\[9\]\[121\] _05524_ _05269_ vssd1 vssd1 vccd1 vccd1
+ _05525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09573_ net256 vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__buf_2
XFILLER_0_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08524_ _04580_ vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__buf_1
XFILLER_0_171_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08455_ addroundkey_data_o\[68\] fifo_bank_register.data_out\[68\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08386_ addroundkey_data_o\[35\] fifo_bank_register.data_out\[35\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__mux2_2
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09007_ _04684_ _05027_ _05028_ _04689_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout530 fifo_bank_register.clk vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__clkbuf_4
Xfanout541 net542 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_2
X_09909_ sub1.data_o\[16\] _05750_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__mux2_1
Xfanout552 net554 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__buf_2
Xfanout563 net564 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__clkbuf_2
Xfanout574 net576 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__buf_2
Xfanout585 net596 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12920_ _07762_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__clkbuf_1
Xfanout596 net259 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _07726_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__clkbuf_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _07172_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15570_ _04369_ _03709_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__nor2_2
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12782_ _07690_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__clkbuf_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _02850_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__clkbuf_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _07136_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__clkbuf_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ net503 _00683_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ fifo_bank_register.bank\[1\]\[99\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[99\]
+ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__a22o_1
X_11664_ fifo_bank_register.bank\[6\]\[39\] _05352_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13403_ _05464_ fifo_bank_register.bank\[0\]\[92\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08018_ sky130_fd_sc_hd__mux2_1
X_10615_ _06381_ _06383_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17171_ net554 _00614_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
X_14383_ fifo_bank_register.bank\[5\]\[91\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[91\]
+ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__a22o_1
X_11595_ _07063_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16122_ net240 ks1.key_reg\[84\] _03906_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux2_2
X_13334_ _07981_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__clkbuf_1
X_10546_ _06323_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__xor2_1
XFILLER_0_165_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ _04014_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _07945_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10477_ addroundkey_data_o\[71\] _06264_ _06248_ vssd1 vssd1 vccd1 vccd1 _06265_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15004_ addroundkey_data_o\[1\] _03208_ _03086_ _03277_ vssd1 vssd1 vccd1 vccd1 _03278_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12216_ _07391_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13196_ fifo_bank_register.bank\[1\]\[123\] _05528_ _07771_ vssd1 vssd1 vccd1 vccd1
+ _07908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12147_ _05293_ fifo_bank_register.bank\[4\]\[11\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07355_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16955_ net432 _00398_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
X_12078_ fifo_bank_register.bank\[5\]\[107\] _05495_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15906_ _05244_ sub1.data_o\[71\] _05199_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__mux2_1
X_11029_ _05615_ _06759_ _06760_ _05567_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16886_ net393 _00329_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18625_ clknet_leaf_23_clk _02054_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[118\]
+ sky130_fd_sc_hd__dfrtp_1
X_15837_ mix1.data_o\[118\] net779 _03841_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15768_ mix1.data_o\[85\] net775 _03808_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18556_ clknet_leaf_77_clk _01985_ net590 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[83\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14719_ sub1.data_o\[53\] sub1.data_o\[117\] _05598_ vssd1 vssd1 vccd1 vccd1 _03022_
+ sky130_fd_sc_hd__mux2_1
X_17507_ net499 _00950_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18487_ clknet_leaf_54_clk _01916_ net615 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_15699_ mix1.data_o\[52\] net764 _03775_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08240_ net75 net74 net77 net76 vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17438_ net565 _00881_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_200_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_15 _04492_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_48 _06358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17369_ net505 _00812_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_172_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_59 addroundkey_data_o\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09625_ _05513_ vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ fifo_bank_register.bank\[9\]\[93\] _05466_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08507_ _04571_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09487_ net226 vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__buf_2
XFILLER_0_109_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08438_ _04535_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08369_ addroundkey_data_o\[27\] fifo_bank_register.data_out\[27\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__mux2_4
XFILLER_0_191_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10400_ mix1.data_o\[63\] _06138_ _06162_ _06163_ sub1.data_o\[63\] vssd1 vssd1 vccd1
+ vccd1 _06196_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11380_ _06950_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10331_ addroundkey_data_o\[55\] _06134_ _06064_ vssd1 vssd1 vccd1 vccd1 _06135_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ sub1.data_o\[50\] _05971_ _06069_ _06070_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _06071_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13050_ fifo_bank_register.bank\[1\]\[53\] _05382_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12001_ fifo_bank_register.bank\[5\]\[70\] _05417_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10193_ _06009_ vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16740_ clknet_leaf_47_clk _00184_ net651 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[31\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13952_ fifo_bank_register.bank\[5\]\[44\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[44\]
+ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__a22o_1
Xfanout393 net397 vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_2
XFILLER_0_199_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12903_ fifo_bank_register.bank\[2\]\[112\] _05506_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07754_ sky130_fd_sc_hd__mux2_1
X_16671_ net413 _00119_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13883_ _02282_ fifo_bank_register.data_out\[36\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15622_ mix1.data_o\[16\] _03487_ _03730_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18410_ clknet_leaf_0_clk _01840_ net622 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[95\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_159_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _07717_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18341_ clknet_leaf_37_clk _01771_ net668 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_9_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15553_ sub1.data_o\[99\] sub1.data_o\[35\] _03671_ vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _07681_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__clkbuf_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _02835_ fifo_bank_register.data_out\[104\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02836_ sky130_fd_sc_hd__mux2_1
X_18272_ clknet_leaf_34_clk _01703_ net662 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[38\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _07127_ vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__clkbuf_1
X_15484_ sub1.data_o\[105\] _03600_ _03653_ sub1.data_o\[41\] vssd1 vssd1 vccd1 vccd1
+ _03655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12696_ fifo_bank_register.bank\[2\]\[14\] _05299_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17223_ net492 _00666_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14435_ fifo_bank_register.bank\[9\]\[97\] _02712_ _02771_ _02772_ _02773_ vssd1
+ vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11647_ _07091_ vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 data_i[110] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__buf_4
XFILLER_0_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput24 data_i[120] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_4
X_17154_ net515 _00597_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 data_i[15] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_4
X_14366_ _02136_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput46 data_i[25] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_4
X_11578_ _07053_ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__clkbuf_1
Xinput57 data_i[35] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__buf_2
Xinput68 data_i[45] vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_4
XFILLER_0_141_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16105_ _04060_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__xor2_4
X_13317_ _05378_ fifo_bank_register.bank\[0\]\[51\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput79 data_i[55] vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__buf_4
X_10529_ sub1.data_o\[78\] _06309_ _06239_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17085_ net430 _00528_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14297_ fifo_bank_register.bank\[0\]\[81\] _02651_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16036_ _05048_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__nor2_1
X_13248_ _05309_ fifo_bank_register.bank\[0\]\[19\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _07899_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17987_ net531 _01430_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_165_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16938_ net452 _00381_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ net437 _00312_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09410_ fifo_bank_register.bank\[9\]\[46\] _05367_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05368_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18608_ clknet_leaf_13_clk _02037_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[101\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09341_ net174 vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__clkbuf_4
X_18539_ clknet_leaf_60_clk _01968_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[66\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09272_ net180 vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__buf_2
XFILLER_0_34_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08223_ net22 net21 net25 net24 vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ _04794_ _04752_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__xor2_1
XFILLER_0_199_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09608_ _05312_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__buf_4
XFILLER_0_218_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10880_ _06627_ vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ net244 vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__buf_2
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ fifo_bank_register.bank\[3\]\[73\] _05424_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07568_ sky130_fd_sc_hd__mux2_1
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11501_ fifo_bank_register.bank\[7\]\[90\] _05459_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12481_ fifo_bank_register.bank\[3\]\[40\] _05354_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14220_ fifo_bank_register.bank\[1\]\[73\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[73\]
+ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__a22o_1
X_11432_ _06977_ vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14151_ fifo_bank_register.bank\[7\]\[66\] _02461_ _02470_ fifo_bank_register.bank\[2\]\[66\]
+ _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__a221o_1
X_11363_ _06941_ vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ fifo_bank_register.bank\[1\]\[78\] _05434_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07859_ sky130_fd_sc_hd__mux2_1
X_10314_ sub1.data_o\[54\] _05971_ _06116_ _06117_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06119_ sky130_fd_sc_hd__a221o_1
X_14082_ _02459_ fifo_bank_register.data_out\[58\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11294_ _06903_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17910_ net396 _01353_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
X_13033_ fifo_bank_register.bank\[1\]\[45\] _05365_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07823_ sky130_fd_sc_hd__mux2_1
X_10245_ net72 mix1.data_o\[49\] _05934_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10176_ _05620_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__buf_2
XFILLER_0_121_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17841_ net451 _01284_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
X_14984_ sub1.data_o\[90\] _03061_ _03065_ sub1.data_o\[58\] vssd1 vssd1 vccd1 vccd1
+ _03258_ sky130_fd_sc_hd__a22o_1
X_17772_ net416 _01215_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16723_ clknet_leaf_43_clk _00167_ net655 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_13935_ _02329_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16654_ net455 _00102_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13866_ fifo_bank_register.bank\[0\]\[34\] _02267_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15605_ _03728_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12817_ fifo_bank_register.bank\[2\]\[71\] _05420_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16585_ net508 _00033_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13797_ fifo_bank_register.bank\[1\]\[27\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__a22o_1
XFILLER_0_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18324_ clknet_leaf_9_clk _01754_ net631 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_15536_ _03687_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _07672_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18255_ clknet_leaf_22_clk _01686_ net646 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15467_ _03643_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12679_ fifo_bank_register.bank\[2\]\[6\] _05282_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ net433 _00649_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
X_14418_ fifo_bank_register.bank\[1\]\[95\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[95\]
+ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__a22o_1
X_18186_ clknet_leaf_18_clk _01617_ net638 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[80\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15398_ sub1.data_o\[75\] _03594_ _03595_ sub1.data_o\[11\] vssd1 vssd1 vccd1 vccd1
+ _03599_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17137_ net393 _00580_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14349_ fifo_bank_register.bank\[5\]\[88\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[88\]
+ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17068_ net464 _00511_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08910_ _04888_ _04932_ _04933_ _04891_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16019_ ks1.key_reg\[8\] _03985_ _03958_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09890_ net34 mix1.data_o\[14\] _05699_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__mux2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ ks1.key_reg\[6\] _04725_ _04864_ net224 vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__a22o_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ ks1.key_reg\[19\] _04742_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_224_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ net168 vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__buf_2
XFILLER_0_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09255_ fifo_bank_register.read_ptr\[3\] _05256_ _05258_ vssd1 vssd1 vccd1 vccd1
+ _05259_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08206_ _04362_ _04363_ _04364_ _04365_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__nor4_1
XFILLER_0_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09186_ _04369_ _04946_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nor2_2
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ mix1.data_o\[28\] _05797_ _05821_ _05822_ sub1.data_o\[28\] vssd1 vssd1 vccd1
+ vccd1 _05861_ sky130_fd_sc_hd__a32o_1
XTAP_5414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput203 key_i[50] vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput214 key_i[60] vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput225 key_i[70] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_4
Xinput236 key_i[80] vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__clkbuf_8
XTAP_5447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput247 key_i[90] vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_4
XTAP_4713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput258 load_i vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__buf_6
XFILLER_0_76_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ _07267_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__clkbuf_1
X_13720_ _08088_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10932_ _05623_ _06670_ _06674_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ fifo_bank_register.bank\[0\]\[11\] _02075_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10863_ addroundkey_data_o\[109\] _06611_ _06612_ vssd1 vssd1 vccd1 vccd1 _06613_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12602_ fifo_bank_register.bank\[3\]\[98\] _05476_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07595_ sky130_fd_sc_hd__mux2_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16370_ net803 _04078_ _04252_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ fifo_bank_register.bank\[9\]\[4\] _08090_ _08146_ _08147_ _08148_ vssd1 vssd1
+ vccd1 vccd1 _08149_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_186_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10794_ net133 ks1.key_reg\[102\] _06402_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__mux2_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ net767 _03456_ _03549_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ fifo_bank_register.bank\[3\]\[65\] _05407_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ net399 _01483_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[42\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_227_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15252_ _03506_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12464_ fifo_bank_register.bank\[3\]\[32\] _05338_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14203_ fifo_bank_register.bank\[6\]\[71\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[71\]
+ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11415_ _06968_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__clkbuf_1
X_15183_ _03447_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12395_ _07485_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ fifo_bank_register.bank\[5\]\[64\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[64\]
+ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11346_ fifo_bank_register.bank\[7\]\[17\] _05305_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14065_ _02444_ fifo_bank_register.data_out\[56\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02445_ sky130_fd_sc_hd__mux2_1
X_11277_ _05508_ fifo_bank_register.bank\[8\]\[113\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13016_ fifo_bank_register.bank\[1\]\[37\] _05348_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10228_ mix1.data_o\[47\] _05876_ _05993_ _05994_ sub1.data_o\[47\] vssd1 vssd1 vccd1
+ vccd1 _06040_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17824_ net409 _01267_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
Xhold2 ks1.key_reg\[61\] vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ _05977_ _05978_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_206_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14967_ sub1.data_o\[111\] _03078_ _03240_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a21oi_2
X_17755_ net482 _01198_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16706_ clknet_leaf_40_clk _00152_ net669 vssd1 vssd1 vccd1 vccd1 round\[3\] sky130_fd_sc_hd__dfrtp_4
X_13918_ _02148_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__clkbuf_4
X_14898_ sub1.data_o\[94\] _03063_ _03092_ sub1.data_o\[62\] vssd1 vssd1 vccd1 vccd1
+ _03173_ sky130_fd_sc_hd__a22o_1
X_17686_ net541 _01129_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
X_13849_ fifo_bank_register.bank\[9\]\[32\] _02226_ _02250_ _02251_ _02252_ vssd1
+ vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a2111o_1
X_16637_ net554 _00085_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16568_ net478 _00016_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18307_ clknet_leaf_1_clk _01738_ net624 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[73\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15519_ sub1.data_o\[53\] _03663_ _03677_ _03673_ vssd1 vssd1 vccd1 vccd1 _03678_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16499_ _04333_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09040_ _04874_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__buf_4
X_18238_ clknet_leaf_32_clk _01669_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18169_ clknet_leaf_77_clk _01600_ net589 vssd1 vssd1 vccd1 vccd1 ks1.col\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09942_ net167 ks1.key_reg\[18\] _05762_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__mux2_2
XFILLER_0_229_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09873_ _05720_ vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__clkbuf_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ mix1.data_o\[46\] _04692_ _04694_ mix1.data_o\[38\] vssd1 vssd1 vccd1 vccd1
+ _04848_ sky130_fd_sc_hd__a22o_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ addroundkey_data_o\[41\] mix1.data_o\[41\] _04778_ vssd1 vssd1 vccd1 vccd1
+ _04779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08686_ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__buf_2
XANTENNA_319 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09307_ fifo_bank_register.bank\[9\]\[13\] _05297_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09238_ _05244_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__buf_6
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09169_ _05178_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11200_ _06854_ vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ _07372_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11131_ _06818_ vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ _05293_ fifo_bank_register.bank\[8\]\[11\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06782_ sky130_fd_sc_hd__mux2_1
XTAP_5211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10013_ sub1.data_o\[26\] _05845_ _05819_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15870_ _03867_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__clkbuf_1
XTAP_5255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14821_ addroundkey_data_o\[13\] _04376_ _05606_ _03096_ vssd1 vssd1 vccd1 vccd1
+ _03097_ sky130_fd_sc_hd__a211o_1
XTAP_5299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ ks1.col\[28\] _05217_ _04911_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__mux2_1
X_17540_ net521 _00983_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _07258_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ fifo_bank_register.bank\[5\]\[18\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[18\]
+ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a22o_1
X_10915_ net18 mix1.data_o\[115\] _05602_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__mux2_1
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17471_ net440 _00914_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
X_14683_ fifo_bank_register.bank\[0\]\[125\] _02993_ _08120_ vssd1 vssd1 vccd1 vccd1
+ _02994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11895_ _07221_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_169_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13634_ fifo_bank_register.bank\[7\]\[10\] _08182_ _08191_ fifo_bank_register.bank\[2\]\[10\]
+ _08194_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__a221o_1
X_16422_ ks1.key_reg\[106\] _03998_ _04281_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__mux2_1
X_10846_ addroundkey_data_o\[107\] _06597_ _06522_ vssd1 vssd1 vccd1 vccd1 _06598_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16353_ _04372_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__buf_4
X_13565_ fifo_bank_register.bank\[1\]\[2\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _08134_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10777_ sub1.data_o\[101\] _06534_ _06478_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15304_ net700 _03363_ _03539_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__mux2_1
X_12516_ fifo_bank_register.bank\[3\]\[57\] _05390_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16284_ _04371_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__buf_4
XFILLER_0_212_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13496_ _08067_ _08073_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__xnor2_1
X_15235_ _03266_ _03326_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__xor2_2
XFILLER_0_180_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18023_ net513 _01466_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_12447_ fifo_bank_register.bank\[3\]\[24\] _05321_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15166_ _03225_ _03280_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__xor2_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12378_ _05524_ fifo_bank_register.bank\[4\]\[121\] _07341_ vssd1 vssd1 vccd1 vccd1
+ _07476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14117_ _02491_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__clkbuf_1
X_11329_ fifo_bank_register.bank\[7\]\[9\] _05288_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06923_ sky130_fd_sc_hd__mux2_1
X_15097_ addroundkey_data_o\[68\] _03072_ _03068_ addroundkey_data_o\[36\] vssd1 vssd1
+ vccd1 vccd1 _03368_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14048_ fifo_bank_register.bank\[0\]\[54\] _02429_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_206_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17807_ net552 _01250_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15999_ net702 _03901_ _03966_ _03967_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08540_ _04588_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17738_ net474 _01181_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08471_ _04552_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17669_ net524 _01112_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09023_ ks1.key_reg\[26\] _04745_ _04746_ net176 vssd1 vssd1 vccd1 vccd1 _05045_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09925_ sub1.data_o\[17\] _05766_ _05751_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09856_ mix1.data_o\[10\] _05677_ _05703_ _05704_ sub1.data_o\[10\] vssd1 vssd1 vccd1
+ vccd1 _05705_ sky130_fd_sc_hd__a32o_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08807_ net177 ks1.key_reg\[27\] _04726_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ addroundkey_data_o\[2\] _05643_ next_addroundkey_ready_o vssd1 vssd1 vccd1
+ vccd1 _05644_ sky130_fd_sc_hd__mux2_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08738_ mix1.data_o\[121\] _04698_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__or2_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_116 mix1.data_o\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_127 mix1.data_o\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_149 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08669_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__clkbuf_4
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _06416_ _06462_ _06464_ _06420_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__a22o_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _07108_ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__clkbuf_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_924 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ _06401_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13350_ _05411_ fifo_bank_register.bank\[0\]\[67\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07990_ sky130_fd_sc_hd__mux2_1
X_10562_ sub1.data_o\[81\] _06339_ _06113_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12301_ _05447_ fifo_bank_register.bank\[4\]\[84\] _07431_ vssd1 vssd1 vccd1 vccd1
+ _07436_ sky130_fd_sc_hd__mux2_1
X_13281_ _05342_ fifo_bank_register.bank\[0\]\[34\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10493_ addroundkey_data_o\[73\] _06278_ _06248_ vssd1 vssd1 vccd1 vccd1 _06279_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15020_ sub1.data_o\[115\] _03079_ _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12232_ _05378_ fifo_bank_register.bank\[4\]\[51\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12163_ _05309_ fifo_bank_register.bank\[4\]\[19\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11114_ _06809_ vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__clkbuf_1
X_16971_ net476 _00414_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_12094_ _07326_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15922_ sub1.data_o\[46\] _03576_ _03892_ sub1.data_o\[110\] vssd1 vssd1 vccd1 vccd1
+ _03899_ sky130_fd_sc_hd__a22o_1
X_11045_ _05276_ fifo_bank_register.bank\[8\]\[3\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15853_ mix1.data_o\[126\] net765 _03729_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__mux2_1
XTAP_5096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14804_ sub1.data_o\[24\] _04376_ _03067_ sub1.data_o\[56\] vssd1 vssd1 vccd1 vccd1
+ _03080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18572_ clknet_leaf_82_clk _02001_ net587 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[99\]
+ sky130_fd_sc_hd__dfrtp_1
X_15784_ _03823_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__clkbuf_1
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _07803_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__clkbuf_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ net394 _00966_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11947_ _07249_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14735_ _03031_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__clkbuf_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14666_ fifo_bank_register.bank\[9\]\[123\] _08089_ _02976_ _02977_ _02978_ vssd1
+ vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a2111o_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ net462 _00897_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_196_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11878_ fifo_bank_register.bank\[5\]\[12\] _05295_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13617_ _08179_ fifo_bank_register.data_out\[8\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _08180_ sky130_fd_sc_hd__mux2_1
X_16405_ _04282_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__clkbuf_1
X_10829_ _06582_ vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17385_ net428 _00828_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_14597_ fifo_bank_register.bank\[5\]\[115\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[115\]
+ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a22o_1
XFILLER_0_223_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13548_ _08087_ _08113_ _08118_ vssd1 vssd1 vccd1 vccd1 _08119_ sky130_fd_sc_hd__or3_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16336_ _04243_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16267_ _03957_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13479_ _08056_ fifo_bank_register.write_ptr\[3\] vssd1 vssd1 vccd1 vccd1 _08058_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_207_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15218_ _03099_ _03344_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__xor2_4
X_18006_ net426 _01449_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput304 net304 vssd1 vssd1 vccd1 vccd1 data_o[24] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16198_ net211 ks1.key_reg\[58\] _03937_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput315 net315 vssd1 vssd1 vccd1 vccd1 data_o[34] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput326 net326 vssd1 vssd1 vccd1 vccd1 data_o[44] sky130_fd_sc_hd__clkbuf_4
Xoutput337 net337 vssd1 vssd1 vccd1 vccd1 data_o[54] sky130_fd_sc_hd__clkbuf_4
X_15149_ _03107_ _03195_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput348 net348 vssd1 vssd1 vccd1 vccd1 data_o[64] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput359 net359 vssd1 vssd1 vccd1 vccd1 data_o[74] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09710_ _05568_ net258 vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__nor2_1
X_09641_ net154 vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__buf_4
XFILLER_0_207_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09572_ _05477_ vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08523_ addroundkey_data_o\[100\] fifo_bank_register.data_out\[100\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__mux2_2
XFILLER_0_195_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ _04543_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08385_ _04507_ vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_163_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09006_ addroundkey_data_o\[2\] mix1.data_o\[2\] _04805_ vssd1 vssd1 vccd1 vccd1
+ _05028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout520 net530 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_2
Xfanout531 net537 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__buf_2
XFILLER_0_217_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout542 net577 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_2
X_09908_ _05607_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__buf_4
Xfanout553 net554 vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout564 net569 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__clkbuf_2
Xfanout575 net576 vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__buf_1
Xfanout586 net588 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__clkbuf_4
X_09839_ _05689_ vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__clkbuf_1
Xfanout597 net602 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_2
XFILLER_0_77_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ fifo_bank_register.bank\[2\]\[87\] _05453_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ fifo_bank_register.bank\[6\]\[104\] _05489_ _07167_ vssd1 vssd1 vccd1 vccd1
+ _07172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12781_ fifo_bank_register.bank\[2\]\[54\] _05384_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07690_ sky130_fd_sc_hd__mux2_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _02849_ fifo_bank_register.data_out\[106\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02850_ sky130_fd_sc_hd__mux2_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ fifo_bank_register.bank\[6\]\[71\] _05420_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14451_ fifo_bank_register.bank\[6\]\[99\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[99\]
+ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ _07099_ vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__clkbuf_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13402_ _08017_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10614_ sub1.data_o\[85\] _06341_ _06386_ _06387_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17170_ net545 _00613_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14382_ _02727_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__clkbuf_1
X_11594_ fifo_bank_register.bank\[6\]\[6\] _05282_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16121_ ks1.col\[20\] _04075_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__xor2_4
XFILLER_0_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13333_ _05394_ fifo_bank_register.bank\[0\]\[59\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07981_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ net234 ks1.key_reg\[79\] _06324_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__mux2_2
XFILLER_0_165_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ net196 ks1.key_reg\[44\] _03907_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_228_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13264_ _05325_ fifo_bank_register.bank\[0\]\[26\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10476_ _06262_ _06263_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__xor2_1
X_15003_ addroundkey_data_o\[65\] _03209_ _03067_ addroundkey_data_o\[33\] vssd1 vssd1
+ vccd1 vccd1 _03277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12215_ _05361_ fifo_bank_register.bank\[4\]\[43\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13195_ _07907_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12146_ _07354_ vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16954_ net456 _00397_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
X_12077_ _07317_ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15905_ _03889_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__clkbuf_1
X_11028_ mix1.data_o\[127\] _05676_ _05758_ _05620_ sub1.data_o\[127\] vssd1 vssd1
+ vccd1 vccd1 _06760_ sky130_fd_sc_hd__a32o_1
XFILLER_0_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16885_ net394 _00328_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18624_ clknet_leaf_24_clk _02053_ net645 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[117\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_205_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15836_ _03850_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__clkbuf_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18555_ clknet_leaf_77_clk _01984_ net590 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[82\]
+ sky130_fd_sc_hd__dfrtp_1
X_15767_ _03814_ vssd1 vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12979_ _07770_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__buf_8
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17506_ net487 _00949_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
X_14718_ _03019_ _04927_ _05219_ _03021_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18486_ clknet_leaf_58_clk _01915_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_15698_ _03778_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17437_ net560 _00880_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14649_ fifo_bank_register.bank\[1\]\[121\] _08111_ _08114_ fifo_bank_register.bank\[8\]\[121\]
+ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_16 _04499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_27 _04577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _05547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 _06368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ net533 _00811_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16319_ net676 _04136_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17299_ net544 _00742_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ fifo_bank_register.bank\[9\]\[115\] _05512_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ net250 vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__buf_2
XFILLER_0_195_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08506_ addroundkey_data_o\[92\] fifo_bank_register.data_out\[92\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__mux2_8
XFILLER_0_210_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09486_ _05419_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08437_ addroundkey_data_o\[59\] fifo_bank_register.data_out\[59\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__mux2_2
XFILLER_0_93_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08368_ _04498_ vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08299_ net190 net192 net193 net189 vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10330_ _06132_ _06133_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ mix1.data_o\[50\] _05952_ _05916_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12000_ _07221_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_218_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10192_ addroundkey_data_o\[42\] _06008_ _05980_ vssd1 vssd1 vccd1 vccd1 _06009_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13951_ _02343_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_199_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout394 net397 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_2
X_12902_ _07753_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__clkbuf_1
X_13882_ fifo_bank_register.bank\[0\]\[36\] _02281_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02282_ sky130_fd_sc_hd__mux2_1
X_16670_ net471 _00118_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15621_ _03737_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12833_ fifo_bank_register.bank\[2\]\[79\] _05436_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07717_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ clknet_leaf_35_clk _01770_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_185_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15552_ _03668_ _04935_ _05560_ _03697_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a31o_1
X_12764_ fifo_bank_register.bank\[2\]\[46\] _05367_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07681_ sky130_fd_sc_hd__mux2_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ fifo_bank_register.bank\[6\]\[63\] _05403_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14503_ fifo_bank_register.bank\[0\]\[104\] _02834_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02835_ sky130_fd_sc_hd__mux2_1
X_18271_ clknet_leaf_32_clk _01702_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[37\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15483_ _03652_ _04784_ _05548_ _03654_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__a31o_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ _07644_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_182_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17222_ net475 _00665_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11646_ fifo_bank_register.bank\[6\]\[30\] _05333_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07091_ sky130_fd_sc_hd__mux2_1
X_14434_ fifo_bank_register.bank\[1\]\[97\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[97\]
+ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 data_i[111] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__buf_2
Xinput25 data_i[121] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_4
X_14365_ _02711_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__clkbuf_1
X_17153_ net573 _00596_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput36 data_i[16] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11577_ fifo_bank_register.bank\[7\]\[127\] _05536_ _06912_ vssd1 vssd1 vccd1 vccd1
+ _07053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput47 data_i[26] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput58 data_i[36] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_2
X_13316_ _07972_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__clkbuf_1
X_16104_ net238 ks1.key_reg\[82\] _03906_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__mux2_2
XFILLER_0_150_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10528_ net104 mix1.data_o\[78\] _06237_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__mux2_1
Xinput69 data_i[46] vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_4
X_17084_ net412 _00527_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
X_14296_ fifo_bank_register.bank\[9\]\[81\] _02631_ _02648_ _02649_ _02650_ vssd1
+ vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_220_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ _07935_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__clkbuf_1
X_16035_ _03995_ _03999_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10459_ addroundkey_data_o\[69\] _06247_ _06248_ vssd1 vssd1 vccd1 vccd1 _06249_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13178_ fifo_bank_register.bank\[1\]\[114\] _05510_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07899_ sky130_fd_sc_hd__mux2_1
X_12129_ _07345_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17986_ net531 _01429_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
X_16937_ net445 _00380_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16868_ net430 _00311_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18607_ clknet_leaf_14_clk _02036_ net629 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[100\]
+ sky130_fd_sc_hd__dfrtp_1
X_15819_ mix1.data_o\[109\] net787 _03841_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16799_ clknet_leaf_63_clk _00243_ net598 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[90\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_220_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09340_ _05320_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18538_ clknet_leaf_60_clk _01967_ net601 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[65\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ _05273_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__clkbuf_1
X_18469_ clknet_leaf_4_clk _01899_ net592 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[109\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08222_ _04379_ vssd1 vssd1 vccd1 vccd1 mix1.next_ready_o sky130_fd_sc_hd__buf_4
XFILLER_0_28_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08986_ _04648_ _04998_ _05003_ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a211o_2
XFILLER_0_220_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09607_ net142 vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09538_ _05454_ vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ fifo_bank_register.bank\[9\]\[65\] _05407_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05408_ sky130_fd_sc_hd__mux2_1
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ _06935_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12480_ _07508_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__buf_4
XFILLER_0_164_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11431_ fifo_bank_register.bank\[7\]\[57\] _05390_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14150_ fifo_bank_register.bank\[5\]\[66\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[66\]
+ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__a22o_1
X_11362_ fifo_bank_register.bank\[7\]\[24\] _05321_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13101_ _07858_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10313_ _04610_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14081_ fifo_bank_register.bank\[0\]\[58\] _02458_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02459_ sky130_fd_sc_hd__mux2_1
X_11293_ _05524_ fifo_bank_register.bank\[8\]\[121\] _06768_ vssd1 vssd1 vccd1 vccd1
+ _06903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _07822_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__clkbuf_1
X_10244_ _06054_ vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17840_ net465 _01283_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10175_ _05757_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__buf_2
XFILLER_0_218_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17771_ net417 _01214_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_14983_ _03253_ _03256_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__nor2_4
X_16722_ clknet_leaf_42_clk _00166_ net659 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_13934_ _02328_ fifo_bank_register.data_out\[41\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16653_ net402 _00101_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_13865_ fifo_bank_register.bank\[9\]\[34\] _02226_ _02264_ _02265_ _02266_ vssd1
+ vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a2111o_1
X_15604_ mix1.data_o\[8\] _03411_ mix1.next_ready_o vssd1 vssd1 vccd1 vccd1 _03728_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12816_ _07708_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__clkbuf_1
X_16584_ net482 _00032_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_13796_ fifo_bank_register.bank\[6\]\[27\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18323_ clknet_leaf_9_clk _01753_ net631 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15535_ sub1.data_o\[60\] _05218_ _04884_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__mux2_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ fifo_bank_register.bank\[2\]\[38\] _05350_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18254_ clknet_leaf_21_clk _01685_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_15466_ sub1.data_o\[35\] _03642_ _03636_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__mux2_1
X_12678_ _07635_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17205_ net411 _00648_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11629_ fifo_bank_register.bank\[6\]\[22\] _05317_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07082_ sky130_fd_sc_hd__mux2_1
X_14417_ fifo_bank_register.bank\[6\]\[95\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[95\]
+ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18185_ clknet_leaf_14_clk _01616_ net629 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[79\]
+ sky130_fd_sc_hd__dfrtp_1
X_15397_ _03019_ _03593_ _05560_ _03598_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17136_ net406 _00579_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14348_ _02696_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14279_ fifo_bank_register.bank\[5\]\[80\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[80\]
+ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a22o_1
X_17067_ net446 _00510_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16018_ _04913_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__xnor2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08840_ ks1.key_reg\[6\] _04729_ _04731_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__or3_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08771_ ks1.key_reg\[19\] _04730_ _04732_ net168 vssd1 vssd1 vccd1 vccd1 _04795_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_178_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ net451 _01412_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_215_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09323_ _05308_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ fifo_bank_register.read_ptr\[0\] _05249_ vssd1 vssd1 vccd1 vccd1 _05258_
+ sky130_fd_sc_hd__xor2_2
XFILLER_0_29_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ sub1.state\[2\] vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_161_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09185_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput204 key_i[51] vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_4
XTAP_5415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput215 key_i[61] vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_4
XFILLER_0_216_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput226 key_i[71] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_8
Xinput237 key_i[81] vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__buf_4
XTAP_5448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput248 key_i[91] vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_215_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08969_ _04706_ _04991_ _04992_ _04710_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a22o_1
Xinput259 reset vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_216_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ fifo_bank_register.bank\[5\]\[60\] _05396_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07267_ sky130_fd_sc_hd__mux2_1
XTAP_4769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ sub1.data_o\[116\] _06513_ _06672_ _06673_ _04610_ vssd1 vssd1 vccd1 vccd1
+ _06674_ sky130_fd_sc_hd__a221o_1
XFILLER_0_211_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10862_ _05792_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__buf_4
X_13650_ fifo_bank_register.bank\[9\]\[11\] _08190_ _02072_ _02073_ _02074_ vssd1
+ vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_168_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12601_ _07594_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13581_ fifo_bank_register.bank\[1\]\[4\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _06381_ _06545_ _06549_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__o21ai_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15320_ _03552_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ _07558_ vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15251_ net775 _03505_ _03498_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12463_ _07522_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11414_ fifo_bank_register.bank\[7\]\[49\] _05373_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14202_ fifo_bank_register.bank\[7\]\[71\] _02542_ _02551_ fifo_bank_register.bank\[2\]\[71\]
+ _02566_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__a221o_1
X_15182_ net760 _03446_ _03425_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ _07484_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__buf_4
XFILLER_0_62_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14133_ _02505_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11345_ _06931_ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14064_ fifo_bank_register.bank\[0\]\[56\] _02443_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02444_ sky130_fd_sc_hd__mux2_1
X_11276_ _06894_ vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13015_ _07813_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10227_ sub1.data_o\[47\] _06038_ _05991_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17823_ net547 _01266_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10158_ net190 ks1.key_reg\[39\] _05920_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__mux2_1
XTAP_5960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 ks1.key_reg\[57\] vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17754_ net501 _01197_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10089_ _05913_ _05754_ sub1.data_o\[34\] _05902_ vssd1 vssd1 vccd1 vccd1 _05914_
+ sky130_fd_sc_hd__a31o_1
X_14966_ sub1.data_o\[15\] _04376_ _03058_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ clknet_leaf_40_clk _00151_ net669 vssd1 vssd1 vccd1 vccd1 round\[2\] sky130_fd_sc_hd__dfrtp_4
X_13917_ _02146_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17685_ net547 _01128_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
X_14897_ _03172_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16636_ net545 _00084_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
X_13848_ fifo_bank_register.bank\[1\]\[32\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[32\]
+ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16567_ net477 _00015_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13779_ fifo_bank_register.bank\[7\]\[25\] _02128_ _02139_ fifo_bank_register.bank\[2\]\[25\]
+ _02189_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18306_ clknet_leaf_1_clk _01737_ net624 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[72\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15518_ sub1.data_o\[21\] sub1.data_o\[85\] _03671_ vssd1 vssd1 vccd1 vccd1 _03677_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16498_ net751 _03435_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_969 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18237_ clknet_leaf_26_clk _01668_ net642 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_15449_ sub1.data_o\[30\] _05235_ _04879_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18168_ clknet_leaf_4_clk _01599_ net591 vssd1 vssd1 vccd1 vccd1 ks1.col\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17119_ net508 _00562_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18099_ net450 _01542_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09941_ _05568_ _05777_ _05781_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09872_ addroundkey_data_o\[11\] _05719_ _05697_ vssd1 vssd1 vccd1 vccd1 _05720_
+ sky130_fd_sc_hd__mux2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _04837_ _04840_ _04843_ _04846_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__or4_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _04662_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__buf_4
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _04362_ _04673_ _04364_ _04365_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__and4_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_309 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_178_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09306_ net162 vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__buf_2
XFILLER_0_113_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09237_ _05241_ _05243_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__xor2_4
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _05177_ _05157_ _05176_ _05119_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ _05107_ _05108_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__or2_2
XFILLER_0_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11130_ _05361_ fifo_bank_register.bank\[8\]\[43\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11061_ _06781_ vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__clkbuf_1
XTAP_5201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ net47 mix1.data_o\[26\] _05817_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14820_ addroundkey_data_o\[77\] _03063_ _03092_ addroundkey_data_o\[45\] vssd1 vssd1
+ vccd1 vccd1 _03096_ sky130_fd_sc_hd__a22o_1
XTAP_5289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14751_ _03039_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11963_ fifo_bank_register.bank\[5\]\[52\] _05380_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07258_ sky130_fd_sc_hd__mux2_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_83_clk clknet_3_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_212_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _02120_ vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__clkbuf_1
X_10914_ _06658_ vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17470_ net442 _00913_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11894_ _07197_ vssd1 vssd1 vccd1 vccd1 _07221_ sky130_fd_sc_hd__buf_8
X_14682_ fifo_bank_register.bank\[9\]\[125\] _08089_ _02990_ _02991_ _02992_ vssd1
+ vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_184_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16421_ _04215_ _03989_ _04290_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_211_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13633_ fifo_bank_register.bank\[5\]\[10\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[10\]
+ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__a22o_1
X_10845_ _06595_ _06596_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__xor2_1
XFILLER_0_183_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16352_ ks1.next_ready_o _04007_ _04251_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a21oi_1
X_10776_ net3 mix1.data_o\[101\] _06476_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__mux2_1
X_13564_ fifo_bank_register.bank\[6\]\[2\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _08133_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15303_ _03543_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12515_ _07549_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13495_ fifo_bank_register.read_ptr\[0\] _08068_ _08072_ vssd1 vssd1 vccd1 vccd1
+ _08073_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16283_ _04214_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__clkbuf_1
X_18022_ net482 _01465_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ _03492_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ _07513_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15165_ _03420_ _03429_ _03430_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a21o_4
XFILLER_0_26_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12377_ _07475_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11328_ _06922_ vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__clkbuf_1
X_14116_ _02490_ fifo_bank_register.data_out\[61\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02491_ sky130_fd_sc_hd__mux2_1
X_15096_ sub1.data_o\[100\] _03057_ _03366_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_227_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14047_ fifo_bank_register.bank\[9\]\[54\] _02388_ _02426_ _02427_ _02428_ vssd1
+ vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__a2111o_1
X_11259_ _06885_ vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17806_ net552 _01249_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15998_ _04865_ _03965_ _03914_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_222_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17737_ net473 _01180_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_14949_ addroundkey_data_o\[105\] _03078_ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_222_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08470_ addroundkey_data_o\[75\] fifo_bank_register.data_out\[75\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__mux2_2
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17668_ net523 _01111_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16619_ net572 _00067_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17599_ net439 _01042_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09022_ _04648_ _05043_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09924_ net37 mix1.data_o\[17\] _05749_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09855_ _05620_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__clkbuf_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _04653_ _04802_ _04817_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__a211o_2
XFILLER_0_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09786_ _05641_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ ks1.key_reg\[25\] _04726_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_217_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_106 fifo_bank_register.data_out\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_117 mix1.data_o\[112\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 mix1.data_o\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08668_ _04363_ sub1.state\[2\] sub1.state\[3\] _04362_ vssd1 vssd1 vccd1 vccd1 _04692_
+ sky130_fd_sc_hd__and4bb_2
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _04617_ mix1.ready_o vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__nand2_4
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10630_ net242 ks1.key_reg\[86\] _06402_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10561_ net108 mix1.data_o\[81\] _06111_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12300_ _07435_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13280_ _07953_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10492_ _06276_ _06277_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__xor2_1
XFILLER_0_224_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ _07399_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12162_ _07362_ vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11113_ _05344_ fifo_bank_register.bank\[8\]\[35\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16970_ net476 _00413_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_12093_ fifo_bank_register.bank\[5\]\[114\] _05510_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15921_ _03717_ _04943_ _05228_ _03898_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a31o_1
X_11044_ _06772_ vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15852_ _03858_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__clkbuf_1
XTAP_5075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__buf_4
XFILLER_0_160_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18571_ clknet_leaf_81_clk _02000_ net586 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[98\]
+ sky130_fd_sc_hd__dfrtp_1
X_15783_ mix1.data_o\[92\] net782 _03819_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_1
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ fifo_bank_register.bank\[1\]\[27\] _05327_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07803_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_56_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ net391 _00965_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14734_ ks1.col\[3\] _05172_ _04916_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__mux2_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ fifo_bank_register.bank\[5\]\[44\] _05363_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ net467 _00896_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14665_ fifo_bank_register.bank\[1\]\[123\] _08111_ _08114_ fifo_bank_register.bank\[8\]\[123\]
+ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__a22o_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _07212_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__clkbuf_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16404_ net827 _03917_ _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13616_ fifo_bank_register.bank\[0\]\[8\] _08178_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08179_ sky130_fd_sc_hd__mux2_1
X_17384_ net430 _00827_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_10828_ addroundkey_data_o\[105\] _06581_ _06522_ vssd1 vssd1 vccd1 vccd1 _06582_
+ sky130_fd_sc_hd__mux2_1
X_14596_ _02917_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16335_ net836 _03936_ _04240_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13547_ _08056_ _08070_ vssd1 vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_171_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10759_ _06381_ _06512_ _06518_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_54_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16266_ _04205_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13478_ _08056_ fifo_bank_register.write_ptr\[3\] vssd1 vssd1 vccd1 vccd1 _08057_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_113_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_207_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18005_ net425 _01448_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15217_ _03478_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12429_ fifo_bank_register.bank\[3\]\[16\] _05303_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput305 net305 vssd1 vssd1 vccd1 vccd1 data_o[25] sky130_fd_sc_hd__buf_2
X_16197_ _04144_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__xor2_2
Xoutput316 net316 vssd1 vssd1 vccd1 vccd1 data_o[35] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput327 net327 vssd1 vssd1 vccd1 vccd1 data_o[45] sky130_fd_sc_hd__clkbuf_4
Xoutput338 net338 vssd1 vssd1 vccd1 vccd1 data_o[55] sky130_fd_sc_hd__clkbuf_4
X_15148_ _03413_ _03414_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__xnor2_4
Xoutput349 net349 vssd1 vssd1 vccd1 vccd1 data_o[65] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15079_ addroundkey_data_o\[99\] _03079_ _03350_ vssd1 vssd1 vccd1 vccd1 _03351_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09640_ _05523_ vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09571_ fifo_bank_register.bank\[9\]\[98\] _05476_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_47_clk clknet_3_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_223_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08522_ _04579_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_222_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08453_ addroundkey_data_o\[67\] fifo_bank_register.data_out\[67\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08384_ addroundkey_data_o\[34\] fifo_bank_register.data_out\[34\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09005_ addroundkey_data_o\[58\] mix1.data_o\[58\] _04665_ vssd1 vssd1 vccd1 vccd1
+ _05027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout510 net511 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout521 net529 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_2
X_09907_ net36 mix1.data_o\[16\] _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__mux2_1
Xfanout532 net537 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_217_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout543 net551 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__buf_2
Xfanout554 net559 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__buf_2
Xfanout565 net569 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_2
Xfanout576 net577 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__clkbuf_2
X_09838_ addroundkey_data_o\[8\] _05688_ next_addroundkey_ready_o vssd1 vssd1 vccd1
+ vccd1 _05689_ sky130_fd_sc_hd__mux2_1
Xfanout587 net588 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout598 net601 vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09769_ addroundkey_data_o\[0\] _05627_ next_addroundkey_ready_o vssd1 vssd1 vccd1
+ vccd1 _05628_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_198_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _07171_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _07689_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__clkbuf_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _07135_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__clkbuf_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ fifo_bank_register.bank\[7\]\[99\] _02785_ _02713_ fifo_bank_register.bank\[2\]\[99\]
+ _02786_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11662_ fifo_bank_register.bank\[6\]\[38\] _05350_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07099_ sky130_fd_sc_hd__mux2_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13401_ _05462_ fifo_bank_register.bank\[0\]\[91\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08017_ sky130_fd_sc_hd__mux2_1
X_10613_ mix1.data_o\[85\] _06129_ _06093_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__o21a_1
X_11593_ _07062_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14381_ _02726_ fifo_bank_register.data_out\[90\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16120_ net148 ks1.key_reg\[116\] _03976_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__mux2_2
X_13332_ _07980_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__clkbuf_1
X_10544_ _05707_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__buf_4
XFILLER_0_162_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16051_ _04012_ _04013_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13263_ _07944_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__clkbuf_1
X_10475_ net226 ks1.key_reg\[71\] _06245_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15002_ sub1.data_o\[97\] _03056_ _03275_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_110_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12214_ _07390_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__clkbuf_1
X_13194_ fifo_bank_register.bank\[1\]\[122\] _05526_ _07771_ vssd1 vssd1 vccd1 vccd1
+ _07907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _05290_ fifo_bank_register.bank\[4\]\[10\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16953_ net469 _00396_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
X_12076_ fifo_bank_register.bank\[5\]\[106\] _05493_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_159_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15904_ sub1.data_o\[102\] _03888_ _03876_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__mux2_1
X_11027_ sub1.data_o\[127\] _06758_ _05609_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_159_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16884_ net394 _00327_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18623_ clknet_leaf_23_clk _02052_ net644 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15835_ mix1.data_o\[117\] net776 _03841_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18554_ clknet_leaf_77_clk _01983_ net589 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[81\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15766_ mix1.data_o\[84\] net783 _03808_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__mux2_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12978_ _07793_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__clkbuf_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ net488 _00948_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_14717_ sub1.data_o\[84\] _03010_ _03020_ sub1.next_ready_o vssd1 vssd1 vccd1 vccd1
+ _03021_ sky130_fd_sc_hd__a22o_1
X_11929_ fifo_bank_register.bank\[5\]\[36\] _05346_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07240_ sky130_fd_sc_hd__mux2_1
X_18485_ clknet_leaf_57_clk _01914_ net602 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_15697_ mix1.data_o\[51\] net763 _03775_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17436_ net560 _00879_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
X_14648_ fifo_bank_register.bank\[6\]\[121\] _08104_ _08107_ fifo_bank_register.bank\[4\]\[121\]
+ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__a22o_1
XFILLER_0_172_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _04508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _04591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_39 _05553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ net532 _00810_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14579_ _02902_ fifo_bank_register.data_out\[112\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02903_ sky130_fd_sc_hd__mux2_1
X_16318_ ks1.next_ready_o _04159_ _04233_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_207_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17298_ net543 _00741_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16249_ ks1.col\[31\] _04192_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_207_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_215_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09623_ net147 vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__buf_2
XFILLER_0_218_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09554_ _05465_ vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08505_ _04570_ vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__clkbuf_1
X_09485_ fifo_bank_register.bank\[9\]\[70\] _05417_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08436_ _04478_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__buf_8
XFILLER_0_148_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08367_ addroundkey_data_o\[26\] fifo_bank_register.data_out\[26\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__mux2_2
XFILLER_0_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08298_ net195 net194 net197 net196 vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_225_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ _05949_ _06067_ _06068_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10191_ _06006_ _06007_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13950_ _02342_ fifo_bank_register.data_out\[43\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout395 net397 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__buf_2
XFILLER_0_199_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12901_ fifo_bank_register.bank\[2\]\[111\] _05504_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07753_ sky130_fd_sc_hd__mux2_1
X_13881_ fifo_bank_register.bank\[9\]\[36\] _02226_ _02278_ _02279_ _02280_ vssd1
+ vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15620_ mix1.data_o\[15\] _03484_ _03730_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__mux2_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12832_ _07716_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15551_ sub1.data_o\[66\] _03691_ _03696_ _03673_ vssd1 vssd1 vccd1 vccd1 _03697_
+ sky130_fd_sc_hd__a22o_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _07680_ vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ fifo_bank_register.bank\[9\]\[104\] _02793_ _02831_ _02832_ _02833_ vssd1
+ vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_210_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18270_ clknet_leaf_33_clk _01701_ net653 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[36\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _07126_ vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15482_ sub1.data_o\[104\] _03600_ _03653_ sub1.data_o\[40\] vssd1 vssd1 vccd1 vccd1
+ _03654_ sky130_fd_sc_hd__a22o_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ fifo_bank_register.bank\[2\]\[13\] _05297_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_204_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ net441 _00664_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14433_ fifo_bank_register.bank\[6\]\[97\] _02718_ _02719_ fifo_bank_register.bank\[4\]\[97\]
+ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11645_ _07078_ vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__buf_4
XFILLER_0_182_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17152_ net558 _00595_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
Xinput15 data_i[112] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14364_ _02710_ fifo_bank_register.data_out\[89\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02711_ sky130_fd_sc_hd__mux2_1
X_11576_ _07052_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__clkbuf_1
Xinput26 data_i[122] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_2
XFILLER_0_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput37 data_i[17] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_4
Xinput48 data_i[27] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_2
XFILLER_0_135_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16103_ ks1.col\[18\] _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__xor2_4
Xinput59 data_i[37] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_8
X_13315_ _05375_ fifo_bank_register.bank\[0\]\[50\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17083_ net434 _00526_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
X_10527_ _06308_ vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_161_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14295_ fifo_bank_register.bank\[1\]\[81\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[81\]
+ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16034_ _03996_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__xor2_2
X_13246_ _05307_ fifo_bank_register.bank\[0\]\[18\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07935_ sky130_fd_sc_hd__mux2_1
X_10458_ _05792_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__buf_4
XFILLER_0_204_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10389_ _06186_ vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__clkbuf_1
X_13177_ _07898_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12128_ _05274_ fifo_bank_register.bank\[4\]\[2\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07345_ sky130_fd_sc_hd__mux2_1
X_17985_ net437 _01428_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
X_16936_ net448 _00379_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
X_12059_ fifo_bank_register.bank\[5\]\[98\] _05476_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16867_ net499 _00310_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15818_ _03741_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_172_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18606_ clknet_leaf_14_clk _02035_ net630 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[99\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_205_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16798_ clknet_leaf_79_clk _00242_ net579 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[89\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_172_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18537_ clknet_leaf_60_clk _01966_ net601 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[64\]
+ sky130_fd_sc_hd__dfrtp_1
X_15749_ mix1.data_o\[76\] net777 _03797_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09270_ fifo_bank_register.bank\[9\]\[1\] _05272_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18468_ clknet_leaf_3_clk _01898_ net584 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[108\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08221_ _04378_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__clkbuf_4
X_17419_ net518 _00862_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18399_ clknet_leaf_24_clk _01829_ net646 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[84\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08985_ _04755_ _05005_ _05007_ _00007_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09606_ _05500_ vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09537_ fifo_bank_register.bank\[9\]\[87\] _05453_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09468_ net219 vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__buf_2
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08419_ _04525_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_175_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09399_ _05360_ vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_163_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ _06976_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ _06940_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10312_ mix1.data_o\[54\] _05952_ _06093_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13100_ fifo_bank_register.bank\[1\]\[77\] _05432_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11292_ _06902_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__clkbuf_1
X_14080_ fifo_bank_register.bank\[9\]\[58\] _02388_ _02455_ _02456_ _02457_ vssd1
+ vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13031_ fifo_bank_register.bank\[1\]\[44\] _05363_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07822_ sky130_fd_sc_hd__mux2_1
X_10243_ addroundkey_data_o\[48\] _06053_ _05980_ vssd1 vssd1 vccd1 vccd1 _06054_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10174_ sub1.data_o\[41\] _05990_ _05991_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_219_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17770_ net422 _01213_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_14982_ addroundkey_data_o\[106\] _03056_ _03255_ vssd1 vssd1 vccd1 vccd1 _03256_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_206_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16721_ clknet_leaf_52_clk _00165_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_13933_ fifo_bank_register.bank\[0\]\[41\] _02327_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16652_ net410 _00100_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13864_ fifo_bank_register.bank\[1\]\[34\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[34\]
+ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a22o_1
X_15603_ _03727_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__clkbuf_1
X_12815_ fifo_bank_register.bank\[2\]\[70\] _05417_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07708_ sky130_fd_sc_hd__mux2_1
X_16583_ net484 _00031_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13795_ fifo_bank_register.bank\[7\]\[27\] _02128_ _02139_ fifo_bank_register.bank\[2\]\[27\]
+ _02203_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18322_ clknet_leaf_9_clk _01752_ net631 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_15534_ _03686_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__clkbuf_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12746_ _07671_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18253_ clknet_leaf_22_clk _01684_ net643 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ sub1.data_o\[67\] _05195_ _03633_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12677_ fifo_bank_register.bank\[2\]\[5\] _05280_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17204_ net471 _00647_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
X_14416_ fifo_bank_register.bank\[7\]\[95\] _02704_ _02713_ fifo_bank_register.bank\[2\]\[95\]
+ _02756_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a221o_1
X_18184_ clknet_leaf_1_clk _01615_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[78\]
+ sky130_fd_sc_hd__dfrtp_1
X_11628_ _07081_ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15396_ sub1.data_o\[74\] _03594_ _03595_ sub1.data_o\[10\] vssd1 vssd1 vccd1 vccd1
+ _03598_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17135_ net399 _00578_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_14347_ _02694_ fifo_bank_register.data_out\[87\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02696_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11559_ fifo_bank_register.bank\[7\]\[118\] _05518_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17066_ net447 _00509_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
X_14278_ _02142_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16017_ _03981_ _03983_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__xnor2_1
X_13229_ _07914_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__buf_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _04741_ _04754_ _04755_ _04757_ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__o221a_2
XFILLER_0_174_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ net465 _01411_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16919_ net565 _00362_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17899_ net417 _01342_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09322_ fifo_bank_register.bank\[9\]\[18\] _05307_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09253_ fifo_bank_register.read_ptr\[3\] _05256_ vssd1 vssd1 vccd1 vccd1 _05257_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08204_ sub1.state\[3\] vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09184_ _05172_ _05194_ _05060_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__mux2_8
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_6106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput205 key_i[52] vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_4
XFILLER_0_122_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput216 key_i[62] vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_4
Xinput227 key_i[72] vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_4
XTAP_5438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput238 key_i[82] vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_4
XTAP_4715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ addroundkey_data_o\[15\] mix1.data_o\[15\] _04663_ vssd1 vssd1 vccd1 vccd1
+ _04992_ sky130_fd_sc_hd__mux2_1
Xinput249 key_i[92] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__buf_2
XTAP_4726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08899_ _04648_ _04910_ _04922_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_224_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10930_ mix1.data_o\[116\] _04626_ _05617_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__o21a_1
XFILLER_0_223_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10861_ _06609_ _06610_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__xor2_1
XFILLER_0_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12600_ fifo_bank_register.bank\[3\]\[97\] _05474_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07594_ sky130_fd_sc_hd__mux2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ fifo_bank_register.bank\[6\]\[4\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ sub1.data_o\[102\] _06513_ _06547_ _06548_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06549_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ fifo_bank_register.bank\[3\]\[64\] _05405_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15250_ _03396_ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__xnor2_4
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12462_ fifo_bank_register.bank\[3\]\[31\] _05336_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14201_ fifo_bank_register.bank\[5\]\[71\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[71\]
+ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11413_ _06967_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__clkbuf_1
X_15181_ _03441_ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12393_ net597 _05249_ _05250_ _07483_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__and4_1
X_14132_ _02504_ fifo_bank_register.data_out\[63\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02505_ sky130_fd_sc_hd__mux2_1
X_11344_ fifo_bank_register.bank\[7\]\[16\] _05303_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14063_ fifo_bank_register.bank\[9\]\[56\] _02388_ _02440_ _02441_ _02442_ vssd1
+ vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a2111o_1
X_11275_ _05506_ fifo_bank_register.bank\[8\]\[112\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06894_ sky130_fd_sc_hd__mux2_1
X_13014_ fifo_bank_register.bank\[1\]\[36\] _05346_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10226_ net70 mix1.data_o\[47\] _05989_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10157_ _05899_ _05970_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__o21ai_4
X_17822_ net566 _01265_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[88\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 ks1.key_reg\[63\] vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ _04624_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__clkbuf_4
X_14965_ sub1.data_o\[79\] _03063_ _03092_ sub1.data_o\[47\] vssd1 vssd1 vccd1 vccd1
+ _03239_ sky130_fd_sc_hd__a22o_1
X_17753_ net516 _01196_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16704_ clknet_leaf_40_clk _00150_ net669 vssd1 vssd1 vccd1 vccd1 round\[1\] sky130_fd_sc_hd__dfrtp_4
X_13916_ fifo_bank_register.bank\[7\]\[40\] _02299_ _02308_ fifo_bank_register.bank\[2\]\[40\]
+ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a221o_1
XFILLER_0_159_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17684_ net517 _01127_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14896_ mix1.data_reg\[64\] _03170_ _03171_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16635_ net552 _00083_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13847_ fifo_bank_register.bank\[6\]\[32\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[32\]
+ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16566_ net477 _00014_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13778_ fifo_bank_register.bank\[5\]\[25\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[25\]
+ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15517_ _03668_ _04777_ _05219_ _03676_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a31o_1
X_18305_ clknet_leaf_34_clk _01736_ net662 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[71\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12729_ _07662_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__clkbuf_1
X_16497_ _03143_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_210_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18236_ clknet_leaf_32_clk _01667_ net653 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_143_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15448_ _03630_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ clknet_leaf_81_clk _01598_ net588 vssd1 vssd1 vccd1 vccd1 ks1.col\[21\] sky130_fd_sc_hd__dfrtp_1
X_15379_ _03586_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_170_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17118_ net485 _00561_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18098_ net458 _01541_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09940_ sub1.data_o\[18\] _05753_ _05779_ _05780_ _04611_ vssd1 vssd1 vccd1 vccd1
+ _05781_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17049_ net539 _00492_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09871_ _05717_ _05718_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__xor2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08822_ _04684_ _04844_ _04845_ _04689_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__a22o_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08753_ _04693_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__buf_4
XFILLER_0_224_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ addroundkey_data_o\[12\] mix1.data_o\[12\] _04666_ vssd1 vssd1 vccd1 vccd1
+ _04708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09305_ _05296_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09236_ _05233_ _05242_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09167_ _05119_ _05176_ _05157_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09098_ _05106_ _05107_ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__nand3_2
XFILLER_0_102_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11060_ _05290_ fifo_bank_register.bank\[8\]\[10\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10011_ _05844_ vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__clkbuf_1
XTAP_5224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ ks1.col\[27\] _05172_ _04911_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__mux2_1
XTAP_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11962_ _07257_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__clkbuf_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13701_ _02118_ fifo_bank_register.data_out\[17\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_196_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10913_ addroundkey_data_o\[114\] _06657_ _06612_ vssd1 vssd1 vccd1 vccd1 _06658_
+ sky130_fd_sc_hd__mux2_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ fifo_bank_register.bank\[1\]\[125\] _08111_ _08114_ fifo_bank_register.bank\[8\]\[125\]
+ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _07220_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16420_ net721 _04136_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__nand2_1
X_13632_ _08099_ vssd1 vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10844_ net138 ks1.key_reg\[107\] _06579_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16351_ net692 _04373_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13563_ fifo_bank_register.bank\[7\]\[2\] _08078_ _08093_ fifo_bank_register.bank\[2\]\[2\]
+ _08131_ vssd1 vssd1 vccd1 vccd1 _08132_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10775_ _06533_ vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__clkbuf_1
X_15302_ net735 _03324_ _03539_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12514_ fifo_bank_register.bank\[3\]\[56\] _05388_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07549_ sky130_fd_sc_hd__mux2_1
X_16282_ ks1.key_reg\[43\] _04008_ _04206_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__mux2_1
X_13494_ _08070_ _08071_ _08056_ vssd1 vssd1 vccd1 vccd1 _08072_ sky130_fd_sc_hd__and3b_1
XFILLER_0_168_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18021_ net483 _01464_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15233_ net755 _03491_ _03425_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ fifo_bank_register.bank\[3\]\[23\] _05319_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15164_ _03420_ _03429_ _05202_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12376_ _05522_ fifo_bank_register.bank\[4\]\[120\] _07341_ vssd1 vssd1 vccd1 vccd1
+ _07475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14115_ fifo_bank_register.bank\[0\]\[61\] _02489_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02490_ sky130_fd_sc_hd__mux2_1
X_11327_ fifo_bank_register.bank\[7\]\[8\] _05286_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06922_ sky130_fd_sc_hd__mux2_1
X_15095_ sub1.data_o\[4\] _04379_ _03059_ _03365_ vssd1 vssd1 vccd1 vccd1 _03366_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_205_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14046_ fifo_bank_register.bank\[1\]\[54\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[54\]
+ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11258_ _05489_ fifo_bank_register.bank\[8\]\[104\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10209_ _06023_ vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11189_ _05420_ fifo_bank_register.bank\[8\]\[71\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17805_ net525 _01248_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
X_15997_ _04865_ _03965_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__or2_1
XTAP_5780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14948_ addroundkey_data_o\[9\] _04377_ _03086_ _03222_ vssd1 vssd1 vccd1 vccd1 _03223_
+ sky130_fd_sc_hd__a211o_1
X_17736_ net420 _01179_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14879_ sub1.data_o\[7\] _04374_ _04658_ _03154_ vssd1 vssd1 vccd1 vccd1 _03155_
+ sky130_fd_sc_hd__a211o_1
X_17667_ net526 _01110_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16618_ net557 _00066_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_17598_ net441 _01041_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16549_ sub1.data_o\[82\] sub1.data_o\[18\] _03574_ vssd1 vssd1 vccd1 vccd1 _04360_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09021_ _04653_ _05017_ _05030_ _05042_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__a211o_2
XFILLER_0_143_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ clknet_leaf_19_clk _01650_ net640 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[49\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09923_ _05765_ vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09854_ _05617_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__clkbuf_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _04820_ _04822_ _04825_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__or4_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ net180 ks1.key_reg\[2\] _05625_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__mux2_2
XFILLER_0_213_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08736_ ks1.key_reg\[25\] _04730_ _04732_ net175 vssd1 vssd1 vccd1 vccd1 _04760_
+ sky130_fd_sc_hd__o31a_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 fifo_bank_register.data_out\[30\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 mix1.data_o\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_129 mix1.data_o\[33\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ _04669_ _04676_ _04683_ _04690_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__or4_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_163_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _04624_ sub1.ready_o vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__nand2_2
XFILLER_0_113_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_187_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10560_ _06338_ vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09219_ _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10491_ net228 ks1.key_reg\[73\] _06245_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__mux2_2
XFILLER_0_122_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ _05375_ fifo_bank_register.bank\[4\]\[50\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ _05307_ fifo_bank_register.bank\[4\]\[18\] _07353_ vssd1 vssd1 vccd1 vccd1
+ _07362_ sky130_fd_sc_hd__mux2_1
X_11112_ _06808_ vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__clkbuf_1
X_12092_ _07325_ vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15920_ sub1.data_o\[45\] _03576_ _03892_ sub1.data_o\[109\] vssd1 vssd1 vccd1 vccd1
+ _03898_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11043_ _05274_ fifo_bank_register.bank\[8\]\[2\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06772_ sky130_fd_sc_hd__mux2_1
XTAP_5021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15851_ mix1.data_o\[125\] net729 _03729_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__mux2_1
XTAP_5054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _03077_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__clkbuf_8
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15782_ _03822_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__clkbuf_1
X_18570_ clknet_leaf_80_clk _01999_ net580 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_203_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12994_ _07802_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__clkbuf_1
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17521_ net392 _00964_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ _03030_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__clkbuf_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ _07248_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ net465 _00895_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14664_ fifo_bank_register.bank\[6\]\[123\] _08104_ _08107_ fifo_bank_register.bank\[4\]\[123\]
+ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__a22o_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11876_ fifo_bank_register.bank\[5\]\[11\] _05293_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07212_ sky130_fd_sc_hd__mux2_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16403_ _04372_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__buf_4
XFILLER_0_223_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ fifo_bank_register.bank\[9\]\[8\] _08090_ _08175_ _08176_ _08177_ vssd1 vssd1
+ vccd1 vccd1 _08178_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17383_ net423 _00826_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10827_ _06578_ _06580_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__xor2_1
XFILLER_0_184_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14595_ _02916_ fifo_bank_register.data_out\[114\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16334_ _04242_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13546_ fifo_bank_register.bank\[9\]\[0\] _08090_ _08102_ _08109_ _08116_ vssd1 vssd1
+ vccd1 vccd1 _08117_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_54_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10758_ sub1.data_o\[99\] _06513_ _06516_ _06517_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06518_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16265_ ks1.key_reg\[35\] _03939_ _04106_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__mux2_1
X_13477_ fifo_bank_register.read_ptr\[3\] vssd1 vssd1 vccd1 vccd1 _08056_ sky130_fd_sc_hd__buf_2
X_10689_ sub1.data_o\[93\] _06454_ _06318_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15216_ net737 _03477_ _03425_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18004_ net425 _01447_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[6\] sky130_fd_sc_hd__dfxtp_1
X_12428_ _07503_ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16196_ net247 ks1.key_reg\[90\] _03918_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput306 net306 vssd1 vssd1 vccd1 vccd1 data_o[26] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput317 net317 vssd1 vssd1 vccd1 vccd1 data_o[36] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ _03207_ _03410_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__xnor2_2
Xoutput328 net328 vssd1 vssd1 vccd1 vccd1 data_o[46] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12359_ _07466_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__clkbuf_1
Xoutput339 net339 vssd1 vssd1 vccd1 vccd1 data_o[56] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15078_ addroundkey_data_o\[3\] _04378_ _05607_ _03349_ vssd1 vssd1 vccd1 vccd1 _03350_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14029_ fifo_bank_register.bank\[6\]\[52\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[52\]
+ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09570_ net255 vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__buf_2
XFILLER_0_222_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08521_ addroundkey_data_o\[99\] fifo_bank_register.data_out\[99\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17719_ net432 _01162_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08452_ _04542_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08383_ _04506_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09004_ _04677_ _05024_ _05025_ _04682_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout500 net507 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__buf_2
XFILLER_0_228_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout511 net530 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09906_ _05601_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__buf_4
Xfanout522 net529 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout533 net535 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
Xfanout544 net551 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_2
Xfanout555 net559 vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_2
Xfanout566 net569 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_2
X_09837_ _05686_ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__xor2_1
Xfanout577 fifo_bank_register.clk vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_4
Xfanout588 net595 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__buf_2
XFILLER_0_225_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout599 net601 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_2
X_09768_ _05624_ _05626_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__xor2_1
XFILLER_0_197_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1088 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08719_ ks1.key_reg\[20\] _04730_ _04732_ net170 vssd1 vssd1 vccd1 vccd1 _04743_
+ sky130_fd_sc_hd__o31a_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ sub1.data_o\[126\] _05236_ _04891_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__mux2_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ fifo_bank_register.bank\[6\]\[70\] _05417_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07135_ sky130_fd_sc_hd__mux2_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _07098_ vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__clkbuf_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_187_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13400_ _08016_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__clkbuf_1
X_10612_ _06126_ _06383_ _06385_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14380_ fifo_bank_register.bank\[0\]\[90\] _02724_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02726_ sky130_fd_sc_hd__mux2_1
X_11592_ fifo_bank_register.bank\[6\]\[5\] _05280_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13331_ _05392_ fifo_bank_register.bank\[0\]\[58\] _07971_ vssd1 vssd1 vccd1 vccd1
+ _07980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10543_ _06250_ _06319_ _06322_ _06254_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16050_ net231 ks1.key_reg\[76\] _03979_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13262_ _05323_ fifo_bank_register.bank\[0\]\[25\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07944_ sky130_fd_sc_hd__mux2_1
X_10474_ _06250_ _06260_ _06261_ _06254_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15001_ sub1.data_o\[1\] _03208_ _03081_ _03274_ vssd1 vssd1 vccd1 vccd1 _03275_
+ sky130_fd_sc_hd__a211o_1
X_12213_ _05359_ fifo_bank_register.bank\[4\]\[42\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13193_ _07906_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12144_ _07341_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__buf_4
XFILLER_0_209_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16952_ net456 _00395_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
X_12075_ _07316_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15903_ _05235_ sub1.data_o\[70\] _05199_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__mux2_1
X_11026_ net31 mix1.data_o\[127\] _05603_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16883_ net405 _00326_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18622_ clknet_leaf_20_clk _02051_ net640 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[115\]
+ sky130_fd_sc_hd__dfrtp_1
X_15834_ _03849_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__clkbuf_1
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_189_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18553_ clknet_leaf_78_clk _01982_ net589 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[80\]
+ sky130_fd_sc_hd__dfrtp_1
X_15765_ _03813_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__clkbuf_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ fifo_bank_register.bank\[1\]\[19\] _05309_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ net487 _00947_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14716_ sub1.data_o\[52\] sub1.data_o\[116\] _05598_ vssd1 vssd1 vccd1 vccd1 _03020_
+ sky130_fd_sc_hd__mux2_1
X_11928_ _07239_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15696_ _03777_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__clkbuf_1
X_18484_ clknet_leaf_56_clk _01913_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17435_ net565 _00878_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
X_14647_ fifo_bank_register.bank\[7\]\[121\] _08077_ _08092_ fifo_bank_register.bank\[2\]\[121\]
+ _02961_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a221o_1
X_11859_ fifo_bank_register.bank\[5\]\[3\] _05276_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 _04517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 _04596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17366_ net496 _00809_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_14578_ fifo_bank_register.bank\[0\]\[112\] _02901_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13529_ _08099_ vssd1 vssd1 vccd1 vccd1 _08100_ sky130_fd_sc_hd__clkbuf_4
X_16317_ net690 _04373_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__nor2_1
XFILLER_0_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17297_ net543 _00740_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16248_ _04138_ _04113_ _04125_ _04111_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or4b_4
XFILLER_0_207_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16179_ net154 ks1.key_reg\[121\] _03902_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__mux2_2
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09622_ _05511_ vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09553_ fifo_bank_register.bank\[9\]\[92\] _05464_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_214_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08504_ addroundkey_data_o\[91\] fifo_bank_register.data_out\[91\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__mux2_4
XFILLER_0_66_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09484_ _05312_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ _04533_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__buf_1
XFILLER_0_93_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08366_ _04497_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_184_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08297_ _04450_ _04451_ _04452_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__or4b_1
XFILLER_0_229_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10190_ net194 ks1.key_reg\[42\] _05997_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout396 net397 vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__clkbuf_2
X_12900_ _07752_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__clkbuf_1
X_13880_ fifo_bank_register.bank\[1\]\[36\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[36\]
+ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__a22o_1
XFILLER_0_199_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ fifo_bank_register.bank\[2\]\[78\] _05434_ _07707_ vssd1 vssd1 vccd1 vccd1
+ _07716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15550_ sub1.data_o\[98\] sub1.data_o\[34\] _03671_ vssd1 vssd1 vccd1 vccd1 _03696_
+ sky130_fd_sc_hd__mux2_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ fifo_bank_register.bank\[2\]\[45\] _05365_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07680_ sky130_fd_sc_hd__mux2_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ fifo_bank_register.bank\[1\]\[104\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[104\]
+ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a22o_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ fifo_bank_register.bank\[6\]\[62\] _05401_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15481_ _03581_ _04784_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__nor2_2
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _07643_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ net495 _00663_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
X_14432_ fifo_bank_register.bank\[7\]\[97\] _02704_ _02713_ fifo_bank_register.bank\[2\]\[97\]
+ _02770_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__a221o_1
X_11644_ _07089_ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17151_ net549 _00594_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14363_ fifo_bank_register.bank\[0\]\[89\] _02709_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02710_ sky130_fd_sc_hd__mux2_2
Xinput16 data_i[113] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11575_ fifo_bank_register.bank\[7\]\[126\] _05534_ _06912_ vssd1 vssd1 vccd1 vccd1
+ _07052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput27 data_i[123] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_4
X_16102_ net146 ks1.key_reg\[114\] _03905_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__mux2_2
Xinput38 data_i[18] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_2
XFILLER_0_220_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13314_ _07937_ vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__buf_4
Xinput49 data_i[28] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_2
X_17082_ net412 _00525_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10526_ addroundkey_data_o\[77\] _06307_ _06248_ vssd1 vssd1 vccd1 vccd1 _06308_
+ sky130_fd_sc_hd__mux2_1
X_14294_ fifo_bank_register.bank\[6\]\[81\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[81\]
+ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16033_ _05559_ _03997_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__xor2_2
X_13245_ _07934_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__clkbuf_1
X_10457_ _06244_ _06246_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13176_ fifo_bank_register.bank\[1\]\[113\] _05508_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07898_ sky130_fd_sc_hd__mux2_1
X_10388_ addroundkey_data_o\[61\] _06185_ _06169_ vssd1 vssd1 vccd1 vccd1 _06186_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12127_ _07344_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17984_ net491 _01427_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16935_ net454 _00378_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
X_12058_ _07307_ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__clkbuf_1
X_11009_ _06743_ vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__clkbuf_1
X_16866_ net486 _00309_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18605_ clknet_leaf_14_clk _02034_ net630 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[98\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15817_ _03840_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16797_ clknet_leaf_73_clk _00241_ net593 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[88\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18536_ clknet_leaf_61_clk _01965_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_1
X_15748_ _03804_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__clkbuf_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18467_ clknet_leaf_3_clk _01897_ net584 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[107\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_158_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_290 sub1.data_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15679_ _03768_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08220_ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__buf_4
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17418_ net521 _00861_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18398_ clknet_leaf_24_clk _01828_ net647 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[83\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17349_ net441 _00792_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08984_ _04863_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__clkbuf_8
XTAP_4908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09605_ fifo_bank_register.bank\[9\]\[109\] _05499_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09536_ net243 vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_210_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_167_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _05406_ vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08418_ addroundkey_data_o\[50\] fifo_bank_register.data_out\[50\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09398_ fifo_bank_register.bank\[9\]\[42\] _05359_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08349_ _04488_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ fifo_bank_register.bank\[7\]\[23\] _05319_ _06936_ vssd1 vssd1 vccd1 vccd1
+ _06940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10311_ _05949_ _06114_ _06115_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11291_ _05522_ fifo_bank_register.bank\[8\]\[120\] _06768_ vssd1 vssd1 vccd1 vccd1
+ _06902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13030_ _07821_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__clkbuf_1
X_10242_ _06051_ _06052_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10173_ _05609_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_218_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14981_ addroundkey_data_o\[10\] _04377_ _03086_ _03254_ vssd1 vssd1 vccd1 vccd1
+ _03255_ sky130_fd_sc_hd__a211o_1
XFILLER_0_195_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16720_ clknet_leaf_52_clk _00164_ net656 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_13932_ fifo_bank_register.bank\[9\]\[41\] _02307_ _02324_ _02325_ _02326_ vssd1
+ vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_96_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13863_ fifo_bank_register.bank\[6\]\[34\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[34\]
+ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__a22o_1
X_16651_ net403 _00099_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15602_ mix1.data_o\[7\] _03402_ mix1.next_ready_o vssd1 vssd1 vccd1 vccd1 _03727_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12814_ _07651_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_202_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13794_ fifo_bank_register.bank\[5\]\[27\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[27\]
+ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__a22o_1
X_16582_ net501 _00030_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18321_ clknet_leaf_8_clk _01751_ net634 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15533_ sub1.data_o\[59\] _05195_ _04884_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__mux2_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ fifo_bank_register.bank\[2\]\[37\] _05348_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18252_ clknet_leaf_21_clk _01683_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_15464_ _03641_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__clkbuf_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _07634_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ fifo_bank_register.bank\[5\]\[95\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[95\]
+ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__a22o_1
X_17203_ net459 _00646_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_167_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11627_ fifo_bank_register.bank\[6\]\[21\] _05315_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15395_ _03019_ _03593_ _05554_ _03597_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__a31o_1
X_18183_ clknet_leaf_1_clk _01614_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[77\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17134_ net395 _00577_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_14346_ _08063_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__buf_6
XFILLER_0_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11558_ _07043_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17065_ net446 _00508_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
X_10509_ addroundkey_data_o\[75\] _06292_ _06248_ vssd1 vssd1 vccd1 vccd1 _06293_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14277_ _02140_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11489_ _07007_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16016_ net192 ks1.key_reg\[40\] _03982_ vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__mux2_1
X_13228_ _07925_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ fifo_bank_register.bank\[1\]\[105\] _05491_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07889_ sky130_fd_sc_hd__mux2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ net467 _01410_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_178_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16918_ net566 _00361_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17898_ net425 _01341_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16849_ net533 _00292_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09321_ net167 vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__buf_2
X_18519_ clknet_leaf_64_clk _01948_ net607 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09252_ fifo_bank_register.write_ptr\[3\] _05251_ _05255_ vssd1 vssd1 vccd1 vccd1
+ _05256_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08203_ sub1.state\[0\] vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09183_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput206 key_i[53] vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_4
XTAP_5428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput217 key_i[63] vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_4
XFILLER_0_228_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ addroundkey_data_o\[111\] mix1.data_o\[111\] _04778_ vssd1 vssd1 vccd1 vccd1
+ _04991_ sky130_fd_sc_hd__mux2_1
Xinput228 key_i[73] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__buf_4
XTAP_4705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput239 key_i[83] vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__buf_4
XFILLER_0_216_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08898_ _04911_ _04913_ _04915_ _04916_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__a221o_2
XFILLER_0_224_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10860_ net140 ks1.key_reg\[109\] _06579_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09519_ fifo_bank_register.bank\[9\]\[81\] _05441_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10791_ mix1.data_o\[102\] _06494_ _06398_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _07557_ vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_192_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12461_ _07521_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14200_ _02565_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__clkbuf_1
X_11412_ fifo_bank_register.bank\[7\]\[48\] _05371_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06967_ sky130_fd_sc_hd__mux2_1
X_15180_ _03353_ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12392_ fifo_bank_register.write_ptr\[2\] _05254_ _05266_ vssd1 vssd1 vccd1 vccd1
+ _07483_ sky130_fd_sc_hd__and3b_1
XFILLER_0_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14131_ fifo_bank_register.bank\[0\]\[63\] _02503_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02504_ sky130_fd_sc_hd__mux2_2
X_11343_ _06930_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14062_ fifo_bank_register.bank\[1\]\[56\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[56\]
+ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__a22o_1
X_11274_ _06893_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13013_ _07812_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__clkbuf_1
X_10225_ _06037_ vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17821_ net561 _01264_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
X_10156_ sub1.data_o\[39\] _05971_ _05974_ _05975_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _05976_ sky130_fd_sc_hd__a221o_1
XTAP_5940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 sub1.state\[4\] vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17752_ net533 _01195_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14964_ _03168_ _03216_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__xnor2_1
X_10087_ sub1.data_o\[34\] _05911_ _05751_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__mux2_1
XTAP_5984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ clknet_leaf_40_clk _00149_ net669 vssd1 vssd1 vccd1 vccd1 round\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13915_ fifo_bank_register.bank\[5\]\[40\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[40\]
+ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_221_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17683_ net546 _01126_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
X_14895_ _03144_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16634_ net549 _00082_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
X_13846_ fifo_bank_register.bank\[7\]\[32\] _02218_ _02227_ fifo_bank_register.bank\[2\]\[32\]
+ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16565_ net473 _00013_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_13777_ _02188_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10989_ _06583_ _06724_ _06725_ _06587_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__a22o_1
X_18304_ clknet_leaf_34_clk _01735_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[70\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15516_ sub1.data_o\[52\] _03663_ _03675_ _03673_ vssd1 vssd1 vccd1 vccd1 _03676_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12728_ fifo_bank_register.bank\[2\]\[29\] _05331_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16496_ _04331_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18235_ clknet_leaf_29_clk _01666_ net635 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15447_ sub1.data_o\[29\] _05227_ _04879_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ _07624_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_210_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18166_ clknet_leaf_81_clk _01597_ net586 vssd1 vssd1 vccd1 vccd1 ks1.col\[20\] sky130_fd_sc_hd__dfrtp_4
X_15378_ sub1.data_o\[4\] _03585_ _03581_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17117_ net483 _00560_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_14329_ fifo_bank_register.bank\[0\]\[85\] _02679_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18097_ net463 _01540_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_180_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17048_ net538 _00491_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ net152 ks1.key_reg\[11\] _05708_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08821_ addroundkey_data_o\[6\] mix1.data_o\[6\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _04845_ sky130_fd_sc_hd__mux2_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _04766_ _04769_ _04772_ _04775_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__or4_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08683_ addroundkey_data_o\[108\] mix1.data_o\[108\] _04663_ vssd1 vssd1 vccd1 vccd1
+ _04707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09304_ fifo_bank_register.bank\[9\]\[12\] _05295_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ _05170_ _05226_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09166_ _05124_ _05125_ _05126_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09097_ sbox1.inversion_to_invert_var\[1\] sbox1.inversion_to_invert_var\[0\] vssd1
+ vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__or2b_1
XFILLER_0_160_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ addroundkey_data_o\[25\] _05843_ _05793_ vssd1 vssd1 vccd1 vccd1 _05844_
+ sky130_fd_sc_hd__mux2_1
XTAP_5214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09999_ _05829_ _05831_ _05832_ _05833_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_215_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11961_ fifo_bank_register.bank\[5\]\[51\] _05378_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ _06655_ _06656_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__xnor2_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _08068_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__clkbuf_8
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ fifo_bank_register.bank\[6\]\[125\] _08104_ _08107_ fifo_bank_register.bank\[4\]\[125\]
+ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11892_ fifo_bank_register.bank\[5\]\[19\] _05309_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13631_ _08096_ vssd1 vssd1 vccd1 vccd1 _08192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10843_ _06583_ _06593_ _06594_ _06587_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13562_ fifo_bank_register.bank\[5\]\[2\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[2\]
+ vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16350_ _04250_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__clkbuf_1
X_10774_ addroundkey_data_o\[100\] _06532_ _06522_ vssd1 vssd1 vccd1 vccd1 _06533_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15301_ _03542_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__clkbuf_1
X_12513_ _07548_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16281_ _04213_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_164_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13493_ _08063_ vssd1 vssd1 vccd1 vccd1 _08071_ sky130_fd_sc_hd__inv_2
XFILLER_0_212_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18020_ net513 _01463_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[22\]
+ sky130_fd_sc_hd__dfxtp_2
X_15232_ _03225_ _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ _07512_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15163_ _03394_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__xnor2_1
X_12375_ _07474_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14114_ fifo_bank_register.bank\[9\]\[61\] _02469_ _02486_ _02487_ _02488_ vssd1
+ vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_205_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11326_ _06921_ vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__clkbuf_1
X_15094_ sub1.data_o\[68\] _03072_ _03068_ sub1.data_o\[36\] vssd1 vssd1 vccd1 vccd1
+ _03365_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14045_ fifo_bank_register.bank\[6\]\[54\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[54\]
+ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11257_ _06884_ vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ addroundkey_data_o\[44\] _06022_ _05980_ vssd1 vssd1 vccd1 vccd1 _06023_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11188_ _06848_ vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17804_ net519 _01247_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
X_10139_ sub1.data_o\[38\] _05959_ _05936_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15996_ _03963_ _03964_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__xor2_4
XTAP_5781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17735_ net439 _01178_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14947_ addroundkey_data_o\[73\] _03063_ _03092_ addroundkey_data_o\[41\] vssd1 vssd1
+ vccd1 vccd1 _03222_ sky130_fd_sc_hd__a22o_1
XFILLER_0_221_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17666_ net513 _01109_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
X_14878_ sub1.data_o\[71\] _03061_ _03065_ sub1.data_o\[39\] vssd1 vssd1 vccd1 vccd1
+ _03154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_216_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16617_ net550 _00065_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_13829_ _02151_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_175_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17597_ net429 _01040_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16548_ _05103_ _04946_ _05554_ _04359_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__a31o_1
XFILLER_0_190_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16479_ net759 _03236_ _04321_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09020_ _05033_ _05035_ _05038_ _05041_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__or4_1
X_18218_ clknet_leaf_15_clk _01649_ net629 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[48\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18149_ clknet_leaf_82_clk _01580_ net585 vssd1 vssd1 vccd1 vccd1 ks1.col\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_142_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09922_ addroundkey_data_o\[16\] _05764_ _05697_ vssd1 vssd1 vccd1 vccd1 _05765_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09853_ sub1.data_o\[10\] _05700_ _05701_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__mux2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _04695_ _04826_ _04827_ _04689_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__a22o_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _05629_ _05639_ _05640_ _05633_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__a22o_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ ks1.key_reg\[1\] _04726_ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__a21oi_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 fifo_bank_register.data_out\[49\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_119 mix1.data_o\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _04684_ _04685_ _04686_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a22o_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08597_ net129 vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_166_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09218_ _05225_ _05226_ _05060_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__mux2_8
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10490_ _06250_ _06274_ _06275_ _06254_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09149_ sbox1.ah_reg\[1\] _05127_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ _07361_ vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11111_ _05342_ fifo_bank_register.bank\[8\]\[34\] _06803_ vssd1 vssd1 vccd1 vccd1
+ _06808_ sky130_fd_sc_hd__mux2_1
X_12091_ fifo_bank_register.bank\[5\]\[113\] _05508_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _06771_ vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_198_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_217_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _03857_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__clkbuf_1
XTAP_5055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _03054_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__buf_6
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ mix1.data_o\[91\] net736 _03819_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__mux2_1
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ fifo_bank_register.bank\[1\]\[26\] _05325_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07802_ sky130_fd_sc_hd__mux2_1
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17520_ net389 _00963_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14732_ ks1.col\[2\] _05559_ _04916_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_169_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ fifo_bank_register.bank\[5\]\[43\] _05361_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17451_ net451 _00894_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14663_ fifo_bank_register.bank\[7\]\[123\] _08077_ _08092_ fifo_bank_register.bank\[2\]\[123\]
+ _02975_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__a221o_1
X_11875_ _07211_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16402_ _04280_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__clkbuf_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13614_ fifo_bank_register.bank\[1\]\[8\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _08177_ sky130_fd_sc_hd__a22o_1
X_10826_ net136 ks1.key_reg\[105\] _06579_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17382_ net417 _00825_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14594_ fifo_bank_register.bank\[0\]\[114\] _02915_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16333_ ks1.key_reg\[66\] _03928_ _04240_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10757_ mix1.data_o\[99\] _06494_ _06398_ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__o21a_1
X_13545_ fifo_bank_register.bank\[1\]\[0\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13476_ _08055_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16264_ _04204_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10688_ net121 mix1.data_o\[93\] _06316_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18003_ net420 _01446_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[5\] sky130_fd_sc_hd__dfxtp_4
X_15215_ _03469_ _03476_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__xnor2_4
X_12427_ fifo_bank_register.bank\[3\]\[15\] _05301_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16195_ _04142_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__xnor2_4
Xoutput307 net307 vssd1 vssd1 vccd1 vccd1 data_o[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput318 net318 vssd1 vssd1 vccd1 vccd1 data_o[37] sky130_fd_sc_hd__clkbuf_4
X_15146_ _03152_ _03216_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ _05504_ fifo_bank_register.bank\[4\]\[111\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07466_ sky130_fd_sc_hd__mux2_1
Xoutput329 net329 vssd1 vssd1 vccd1 vccd1 data_o[47] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11309_ _06911_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__buf_4
X_15077_ addroundkey_data_o\[67\] _03064_ _03084_ addroundkey_data_o\[35\] vssd1 vssd1
+ vccd1 vccd1 _03349_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12289_ _07429_ vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14028_ fifo_bank_register.bank\[7\]\[52\] _02380_ _02389_ fifo_bank_register.bank\[2\]\[52\]
+ _02411_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a221o_1
XFILLER_0_219_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15979_ _03949_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__clkbuf_1
X_08520_ _04478_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__buf_6
XFILLER_0_222_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17718_ net432 _01161_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_188_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_194_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08451_ addroundkey_data_o\[66\] fifo_bank_register.data_out\[66\] _04534_ vssd1
+ vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__mux2_1
X_17649_ net392 _01092_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08382_ addroundkey_data_o\[33\] fifo_bank_register.data_out\[33\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__mux2_4
XFILLER_0_163_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09003_ addroundkey_data_o\[114\] mix1.data_o\[114\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _05025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout501 net507 vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__buf_2
X_09905_ _05748_ vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 net520 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__buf_2
Xfanout523 net529 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__buf_2
XFILLER_0_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout534 net535 vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_2
Xfanout545 net551 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__buf_2
Xfanout556 net559 vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_2
Xfanout567 net569 vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_2
X_09836_ net246 ks1.key_reg\[8\] _05625_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__mux2_1
Xfanout578 net580 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__clkbuf_4
Xfanout589 net595 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09767_ net130 ks1.key_reg\[0\] _05625_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _04735_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__buf_4
X_09698_ _05564_ vssd1 vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__clkbuf_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ sub1.state\[0\] vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__inv_2
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11660_ fifo_bank_register.bank\[6\]\[37\] _05348_ _07090_ vssd1 vssd1 vccd1 vccd1
+ _07098_ sky130_fd_sc_hd__mux2_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _06090_ _06342_ sub1.data_o\[85\] _06384_ vssd1 vssd1 vccd1 vccd1 _06385_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11591_ _07061_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13330_ _07979_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__clkbuf_1
X_10542_ mix1.data_o\[79\] _06296_ _06320_ _06321_ sub1.data_o\[79\] vssd1 vssd1 vccd1
+ vccd1 _06322_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13261_ _07943_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10473_ mix1.data_o\[71\] _06217_ _06241_ _06242_ sub1.data_o\[71\] vssd1 vssd1 vccd1
+ vccd1 _06261_ sky130_fd_sc_hd__a32o_1
XFILLER_0_228_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15000_ sub1.data_o\[65\] _03209_ _03067_ sub1.data_o\[33\] vssd1 vssd1 vccd1 vccd1
+ _03274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12212_ _07389_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13192_ fifo_bank_register.bank\[1\]\[121\] _05524_ _07771_ vssd1 vssd1 vccd1 vccd1
+ _07906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_202_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12143_ _07352_ vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16951_ net470 _00394_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
X_12074_ fifo_bank_register.bank\[5\]\[105\] _05491_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15902_ _03887_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__clkbuf_1
X_11025_ _06757_ vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16882_ net389 _00325_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18621_ clknet_leaf_16_clk _02050_ net634 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15833_ mix1.data_o\[116\] net688 _03841_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__mux2_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18552_ clknet_leaf_64_clk _01981_ net599 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[79\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15764_ mix1.data_o\[83\] net786 _03808_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__mux2_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12976_ _07792_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__clkbuf_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ net487 _00946_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_14715_ _05103_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_169_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ fifo_bank_register.bank\[5\]\[35\] _05344_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07239_ sky130_fd_sc_hd__mux2_1
X_18483_ clknet_leaf_55_clk _01912_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_15695_ mix1.data_o\[50\] net753 _03775_ vssd1 vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__mux2_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ net548 _00877_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
X_14646_ fifo_bank_register.bank\[5\]\[121\] _08096_ _08099_ fifo_bank_register.bank\[3\]\[121\]
+ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a22o_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11858_ _07202_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10809_ net6 mix1.data_o\[104\] _06316_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_19 _04529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17365_ net534 _00808_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14577_ fifo_bank_register.bank\[9\]\[112\] _02874_ _02898_ _02899_ _02900_ vssd1
+ vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a2111o_1
X_11789_ _07165_ vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16316_ _04215_ _04148_ _04232_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ _08098_ vssd1 vssd1 vccd1 vccd1 _08099_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17296_ net544 _00739_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_941 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16247_ net689 ks1.next_ready_o _04190_ _04191_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13459_ _05520_ fifo_bank_register.bank\[0\]\[119\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16178_ ks1.col\[25\] _04127_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__xor2_4
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15129_ _03372_ _03397_ _06630_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09621_ fifo_bank_register.bank\[9\]\[114\] _05510_ _05502_ vssd1 vssd1 vccd1 vccd1
+ _05511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09552_ net249 vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__buf_2
XFILLER_0_223_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_222_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08503_ _04569_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ net225 vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_176_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ addroundkey_data_o\[58\] fifo_bank_register.data_out\[58\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__mux2_2
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ addroundkey_data_o\[25\] fifo_bank_register.data_out\[25\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08296_ net240 net241 net239 net238 vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__and4b_1
XFILLER_0_18_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09819_ addroundkey_data_o\[6\] _05671_ next_addroundkey_ready_o vssd1 vssd1 vccd1
+ vccd1 _05672_ sky130_fd_sc_hd__mux2_1
Xfanout397 net444 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__buf_2
XFILLER_0_214_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _07715_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12761_ _07679_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ fifo_bank_register.bank\[6\]\[104\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[104\]
+ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__a22o_1
XFILLER_0_210_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _07125_ vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__clkbuf_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _05103_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__buf_4
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ fifo_bank_register.bank\[2\]\[12\] _05295_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ fifo_bank_register.bank\[6\]\[29\] _05331_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14431_ fifo_bank_register.bank\[5\]\[97\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[97\]
+ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__a22o_1
XFILLER_0_193_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17150_ net574 _00593_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11574_ _07051_ vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__clkbuf_1
X_14362_ fifo_bank_register.bank\[9\]\[89\] _02631_ _02706_ _02707_ _02708_ vssd1
+ vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_25_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput17 data_i[114] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
Xinput28 data_i[124] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__buf_2
XFILLER_0_135_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16101_ _04058_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__clkbuf_1
Xinput39 data_i[19] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_4
X_13313_ _07970_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__clkbuf_1
X_10525_ _06305_ _06306_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__xor2_1
X_14293_ fifo_bank_register.bank\[7\]\[81\] _02623_ _02632_ fifo_bank_register.bank\[2\]\[81\]
+ _02647_ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__a221o_1
X_17081_ net434 _00524_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13244_ _05305_ fifo_bank_register.bank\[0\]\[17\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07934_ sky130_fd_sc_hd__mux2_1
X_16032_ net137 ks1.key_reg\[106\] _03979_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10456_ net223 ks1.key_reg\[69\] _06245_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13175_ _07897_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__clkbuf_1
X_10387_ _06183_ _06184_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__xor2_1
XFILLER_0_209_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12126_ _05272_ fifo_bank_register.bank\[4\]\[1\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07344_ sky130_fd_sc_hd__mux2_1
X_17983_ net491 _01426_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
X_16934_ net445 _00377_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
X_12057_ fifo_bank_register.bank\[5\]\[97\] _05474_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07307_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11008_ addroundkey_data_o\[124\] _06742_ _05696_ vssd1 vssd1 vccd1 vccd1 _06743_
+ sky130_fd_sc_hd__mux2_1
X_16865_ net479 _00308_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18604_ clknet_leaf_14_clk _02033_ net630 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[97\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15816_ mix1.data_o\[108\] net758 _03830_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16796_ clknet_leaf_26_clk _00240_ net649 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[87\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18535_ clknet_leaf_60_clk _01964_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_158_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15747_ mix1.data_o\[75\] net760 _03797_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12959_ fifo_bank_register.bank\[1\]\[10\] _05290_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07784_ sky130_fd_sc_hd__mux2_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18466_ clknet_leaf_3_clk _01896_ net583 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[106\]
+ sky130_fd_sc_hd__dfrtp_2
X_15678_ mix1.data_o\[42\] net732 _03764_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 fifo_bank_register.data_out\[105\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_291 sub1.data_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17417_ net514 _00860_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_14629_ _02946_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__clkbuf_1
X_18397_ clknet_leaf_18_clk _01827_ net638 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[82\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17348_ net494 _00791_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17279_ net549 _00722_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ ks1.key_reg\[7\] _04725_ _05006_ net235 vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_228_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_223_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09604_ net140 vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__buf_2
XFILLER_0_196_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_218_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_196_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09535_ _05452_ vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ fifo_bank_register.bank\[9\]\[64\] _05405_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08417_ _04524_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__buf_1
XFILLER_0_175_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09397_ net194 vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_171_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08348_ addroundkey_data_o\[17\] fifo_bank_register.data_out\[17\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__mux2_2
XFILLER_0_149_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08279_ _04414_ _04419_ _04424_ _04435_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__or4_4
XFILLER_0_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10310_ _06090_ _05972_ sub1.data_o\[54\] _06079_ vssd1 vssd1 vccd1 vccd1 _06115_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_225_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11290_ _06901_ vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10241_ net200 ks1.key_reg\[48\] _05920_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__mux2_1
X_10172_ net64 mix1.data_o\[41\] _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14980_ addroundkey_data_o\[74\] _03209_ _03067_ addroundkey_data_o\[42\] vssd1 vssd1
+ vccd1 vccd1 _03254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13931_ fifo_bank_register.bank\[1\]\[41\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[41\]
+ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__a22o_1
XFILLER_0_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ net409 _00098_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
X_13862_ fifo_bank_register.bank\[7\]\[34\] _02218_ _02227_ fifo_bank_register.bank\[2\]\[34\]
+ _02263_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15601_ _03726_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12813_ _07706_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__clkbuf_1
X_16581_ net484 _00029_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13793_ _02202_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18320_ clknet_leaf_9_clk _01750_ net633 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15532_ _03685_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__clkbuf_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _07670_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_201_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ clknet_leaf_23_clk _01682_ net643 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ sub1.data_o\[34\] _03640_ _03636_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ fifo_bank_register.bank\[2\]\[4\] _05278_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17202_ net453 _00645_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ _02755_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__clkbuf_1
X_18182_ clknet_leaf_0_clk _01613_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[76\]
+ sky130_fd_sc_hd__dfrtp_1
X_11626_ _07080_ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15394_ sub1.data_o\[73\] _03594_ _03595_ sub1.data_o\[9\] vssd1 vssd1 vccd1 vccd1
+ _03597_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17133_ net415 _00576_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14345_ fifo_bank_register.bank\[0\]\[87\] _02693_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11557_ fifo_bank_register.bank\[7\]\[117\] _05516_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17064_ net446 _00507_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
X_10508_ _06290_ _06291_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14276_ _02138_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__clkbuf_4
X_11488_ fifo_bank_register.bank\[7\]\[84\] _05447_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_204_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16015_ _03918_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__buf_4
X_10439_ net93 mix1.data_o\[68\] _06158_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__mux2_1
X_13227_ _05288_ fifo_bank_register.bank\[0\]\[9\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ _07888_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_209_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ fifo_bank_register.bank\[5\]\[122\] _05526_ _07198_ vssd1 vssd1 vccd1 vccd1
+ _07334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13089_ _07852_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__clkbuf_1
X_17966_ net463 _01409_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16917_ net549 _00360_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17897_ net429 _01340_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16848_ net503 _00291_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16779_ clknet_leaf_79_clk _00223_ net579 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[70\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09320_ _05306_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18518_ clknet_leaf_64_clk _01947_ net603 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09251_ _05252_ _05253_ _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__a21o_1
XFILLER_0_186_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18449_ clknet_leaf_73_clk _01879_ net593 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[89\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_185_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08202_ sub1.state\[1\] vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09182_ _05163_ _05192_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput207 key_i[54] vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_4
XTAP_5429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput218 key_i[64] vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_4
Xinput229 key_i[74] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__buf_4
XFILLER_0_215_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08966_ mix1.data_o\[103\] _04698_ _04701_ _04989_ vssd1 vssd1 vccd1 vccd1 _04990_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_228_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08897_ _04645_ _04918_ _04863_ _04920_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_224_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_196_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09518_ net237 vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__clkbuf_4
X_10790_ _06491_ _06545_ _06546_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ net212 vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__buf_2
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12460_ fifo_bank_register.bank\[3\]\[30\] _05333_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _06966_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__clkbuf_1
X_12391_ _07482_ vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14130_ fifo_bank_register.bank\[9\]\[63\] _02469_ _02500_ _02501_ _02502_ vssd1
+ vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__a2111o_1
X_11342_ fifo_bank_register.bank\[7\]\[15\] _05301_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14061_ fifo_bank_register.bank\[6\]\[56\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[56\]
+ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__a22o_1
X_11273_ _05504_ fifo_bank_register.bank\[8\]\[111\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13012_ fifo_bank_register.bank\[1\]\[35\] _05344_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07812_ sky130_fd_sc_hd__mux2_1
X_10224_ addroundkey_data_o\[46\] _06036_ _05980_ vssd1 vssd1 vccd1 vccd1 _06037_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17820_ net548 _01263_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
X_10155_ mix1.data_o\[39\] _05952_ _05916_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__o21a_1
XTAP_5930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17751_ net532 _01194_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ net56 mix1.data_o\[34\] _05749_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__mux2_1
X_14963_ _03237_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 ks1.key_reg\[60\] vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16702_ clknet_leaf_40_clk _00148_ net669 vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_226_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13914_ _02142_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17682_ net543 _01125_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
X_14894_ _03090_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16633_ net554 _00081_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13845_ fifo_bank_register.bank\[5\]\[32\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[32\]
+ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_202_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16564_ net474 _00012_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_13776_ _02187_ fifo_bank_register.data_out\[24\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10988_ mix1.data_o\[122\] _05676_ _06575_ _06576_ sub1.data_o\[122\] vssd1 vssd1
+ vccd1 vccd1 _06725_ sky130_fd_sc_hd__a32o_1
X_18303_ clknet_leaf_34_clk _01734_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[69\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_146_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15515_ sub1.data_o\[20\] sub1.data_o\[84\] _03671_ vssd1 vssd1 vccd1 vccd1 _03675_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _07661_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__clkbuf_1
X_16495_ net687 _03424_ _04321_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18234_ clknet_leaf_27_clk _01665_ net641 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15446_ _03629_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12658_ fifo_bank_register.bank\[3\]\[125\] _05532_ _07485_ vssd1 vssd1 vccd1 vccd1
+ _07624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11609_ fifo_bank_register.bank\[6\]\[13\] _05297_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07071_ sky130_fd_sc_hd__mux2_1
X_18165_ clknet_leaf_75_clk _01596_ net587 vssd1 vssd1 vccd1 vccd1 ks1.col\[19\] sky130_fd_sc_hd__dfrtp_2
X_15377_ sub1.data_o\[36\] sub1.data_o\[100\] _05202_ vssd1 vssd1 vccd1 vccd1 _03585_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12589_ _07588_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_10_clk clknet_3_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17116_ net502 _00559_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14328_ fifo_bank_register.bank\[9\]\[85\] _02631_ _02676_ _02677_ _02678_ vssd1
+ vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18096_ net458 _01539_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_180_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17047_ net540 _00490_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14259_ fifo_bank_register.bank\[7\]\[78\] _02542_ _02551_ fifo_bank_register.bank\[2\]\[78\]
+ _02616_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ addroundkey_data_o\[62\] mix1.data_o\[62\] _04662_ vssd1 vssd1 vccd1 vccd1
+ _04844_ sky130_fd_sc_hd__mux2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _04661_ _04773_ _04774_ _04656_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ net564 _01392_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_77_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08682_ _04705_ _04681_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__nor2_4
XFILLER_0_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_221_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09303_ net161 vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__buf_2
XFILLER_0_118_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _05239_ _05240_ _05234_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__o21a_2
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09165_ sbox1.ah_reg\[2\] sbox1.ah_reg\[1\] vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__xor2_1
XFILLER_0_185_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09096_ _05105_ sbox1.inversion_to_invert_var\[3\] vssd1 vssd1 vccd1 vccd1 _05107_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_226_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09998_ _04609_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__clkbuf_4
XTAP_5237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08949_ addroundkey_data_o\[23\] mix1.data_o\[23\] _04656_ vssd1 vssd1 vccd1 vccd1
+ _04973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _07256_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__clkbuf_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ net146 ks1.key_reg\[114\] _04639_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__mux2_4
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _07219_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _08092_ vssd1 vssd1 vccd1 vccd1 _08191_ sky130_fd_sc_hd__clkbuf_4
X_10842_ mix1.data_o\[107\] _06463_ _06575_ _06576_ sub1.data_o\[107\] vssd1 vssd1
+ vccd1 vccd1 _06594_ sky130_fd_sc_hd__a32o_1
XFILLER_0_211_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13561_ _08130_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10773_ _06530_ _06531_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__xnor2_1
X_15300_ net693 _03283_ _03539_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12512_ fifo_bank_register.bank\[3\]\[55\] _05386_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07548_ sky130_fd_sc_hd__mux2_1
X_16280_ ks1.key_reg\[42\] _04000_ _04206_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__mux2_1
X_13492_ _05262_ _08069_ vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15231_ _03200_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_168_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12443_ fifo_bank_register.bank\[3\]\[22\] _05317_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_191_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15162_ _03152_ _03427_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_164_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12374_ _05520_ fifo_bank_register.bank\[4\]\[119\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14113_ fifo_bank_register.bank\[1\]\[61\] _02478_ _02479_ fifo_bank_register.bank\[8\]\[61\]
+ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a22o_1
X_11325_ fifo_bank_register.bank\[7\]\[7\] _05284_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06921_ sky130_fd_sc_hd__mux2_1
X_15093_ _03364_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14044_ fifo_bank_register.bank\[7\]\[54\] _02380_ _02389_ fifo_bank_register.bank\[2\]\[54\]
+ _02425_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__a221o_1
X_11256_ _05487_ fifo_bank_register.bank\[8\]\[103\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06884_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _06020_ _06021_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_1210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11187_ _05417_ fifo_bank_register.bank\[8\]\[70\] _06847_ vssd1 vssd1 vccd1 vccd1
+ _06848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10138_ net60 mix1.data_o\[38\] _05934_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__mux2_1
X_17803_ net518 _01246_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15995_ net189 ks1.key_reg\[38\] _03910_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__mux2_2
XFILLER_0_94_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_59_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17734_ net473 _01177_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14946_ sub1.data_o\[105\] _03078_ _03220_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__a21oi_2
X_10069_ net183 ks1.key_reg\[32\] _05762_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__mux2_2
XFILLER_0_221_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17665_ net572 _01108_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14877_ _03142_ _03152_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16616_ net574 _00064_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13828_ fifo_bank_register.bank\[6\]\[30\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a22o_1
XFILLER_0_203_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17596_ net408 _01039_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_175_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16547_ sub1.data_o\[113\] _05197_ _04358_ _03594_ vssd1 vssd1 vccd1 vccd1 _04359_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_169_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13759_ fifo_bank_register.bank\[0\]\[22\] _02172_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16478_ _04322_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18217_ clknet_leaf_0_clk _01648_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15429_ sub1.data_o\[21\] _03606_ _03619_ _03611_ vssd1 vssd1 vccd1 vccd1 _03620_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18148_ clknet_leaf_82_clk _01579_ net587 vssd1 vssd1 vccd1 vccd1 ks1.col\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18079_ net566 _01522_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[81\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09921_ _05761_ _05763_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09852_ _05609_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__buf_4
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ addroundkey_data_o\[3\] mix1.data_o\[3\] _04656_ vssd1 vssd1 vccd1 vccd1
+ _04827_ sky130_fd_sc_hd__mux2_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ mix1.data_o\[2\] _05586_ _05618_ _05621_ sub1.data_o\[2\] vssd1 vssd1 vccd1
+ vccd1 _05640_ sky130_fd_sc_hd__a32o_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08734_ ks1.key_reg\[1\] _04730_ _04732_ net169 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__o31a_1
XFILLER_0_197_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 fifo_bank_register.data_out\[87\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _04688_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_166_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _05137_ _05184_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09148_ _05156_ _05158_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__nor2_2
XFILLER_0_47_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09079_ _05091_ _05071_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_163_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11110_ _06807_ vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12090_ _07324_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11041_ _05272_ fifo_bank_register.bank\[8\]\[1\] _06769_ vssd1 vssd1 vccd1 vccd1
+ _06771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _03071_ _03075_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__nor2_4
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15780_ _03821_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__clkbuf_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12992_ _07801_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__clkbuf_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _03029_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_203_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _07247_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ net453 _00893_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ fifo_bank_register.bank\[5\]\[123\] _08096_ _08099_ fifo_bank_register.bank\[3\]\[123\]
+ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11874_ fifo_bank_register.bank\[5\]\[10\] _05290_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07211_ sky130_fd_sc_hd__mux2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16401_ ks1.key_reg\[96\] _03904_ _04264_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__mux2_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13613_ fifo_bank_register.bank\[6\]\[8\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _08176_ sky130_fd_sc_hd__a22o_1
XFILLER_0_211_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17381_ net437 _00824_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _05707_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__buf_4
X_14593_ fifo_bank_register.bank\[9\]\[114\] _02874_ _02912_ _02913_ _02914_ vssd1
+ vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_131_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16332_ _04241_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13544_ _08114_ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__clkbuf_4
X_10756_ _06491_ _06512_ _06515_ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16263_ net820 _03930_ _04106_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__mux2_1
X_13475_ _05536_ fifo_bank_register.bank\[0\]\[127\] _07914_ vssd1 vssd1 vccd1 vccd1
+ _08055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10687_ _06453_ vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18002_ net422 _01445_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[4\] sky130_fd_sc_hd__dfxtp_1
X_15214_ _03418_ _03475_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__xor2_2
XFILLER_0_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12426_ _07502_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__clkbuf_1
X_16194_ net155 ks1.key_reg\[122\] _03902_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__mux2_2
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15145_ _03412_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__clkbuf_1
Xoutput308 net308 vssd1 vssd1 vccd1 vccd1 data_o[28] sky130_fd_sc_hd__clkbuf_4
Xoutput319 net319 vssd1 vssd1 vccd1 vccd1 data_o[38] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12357_ _07465_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11308_ net597 _05249_ _05250_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__and4_1
X_15076_ sub1.data_o\[99\] _03079_ _03347_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_227_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12288_ _05434_ fifo_bank_register.bank\[4\]\[78\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07429_ sky130_fd_sc_hd__mux2_1
X_14027_ fifo_bank_register.bank\[5\]\[52\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[52\]
+ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a22o_1
X_11239_ _05470_ fifo_bank_register.bank\[8\]\[95\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15978_ ks1.key_reg\[4\] _03948_ _04373_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14929_ addroundkey_data_o\[89\] _03063_ _03092_ addroundkey_data_o\[57\] vssd1 vssd1
+ vccd1 vccd1 _03204_ sky130_fd_sc_hd__a22o_1
X_17717_ net412 _01160_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[111\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08450_ _04541_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_148_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17648_ net389 _01091_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ _04505_ vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17579_ net450 _01022_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09002_ addroundkey_data_o\[82\] mix1.data_o\[82\] _04662_ vssd1 vssd1 vccd1 vccd1
+ _05024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ addroundkey_data_o\[15\] _05747_ _05697_ vssd1 vssd1 vccd1 vccd1 _05748_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout502 net507 vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_2
Xfanout513 net520 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_2
Xfanout524 net529 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout535 net537 vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__clkbuf_2
Xfanout546 net551 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_2
X_09835_ _05629_ _05684_ _05685_ _05633_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a22o_1
Xfanout557 net559 vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_2
Xfanout568 net569 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout579 net580 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__buf_4
XFILLER_0_119_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09766_ _04639_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__buf_4
XFILLER_0_154_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08717_ _04740_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09697_ sub1.data_o\[125\] _05228_ _04891_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__mux2_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08648_ addroundkey_data_o\[28\] mix1.data_o\[28\] _04666_ vssd1 vssd1 vccd1 vccd1
+ _04672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _04608_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_187_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _05584_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__clkbuf_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11590_ fifo_bank_register.bank\[6\]\[4\] _05278_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10541_ _05619_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260_ _05321_ fifo_bank_register.bank\[0\]\[24\] _07938_ vssd1 vssd1 vccd1 vccd1
+ _07943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10472_ sub1.data_o\[71\] _06259_ _06239_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12211_ _05357_ fifo_bank_register.bank\[4\]\[41\] _07387_ vssd1 vssd1 vccd1 vccd1
+ _07389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ _07905_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_206_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12142_ _05288_ fifo_bank_register.bank\[4\]\[9\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16950_ net411 _00393_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
X_12073_ _07315_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_194_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15901_ sub1.data_o\[101\] _03886_ _03876_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__mux2_1
X_11024_ addroundkey_data_o\[126\] _06756_ _05696_ vssd1 vssd1 vccd1 vccd1 _06757_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16881_ net393 _00324_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15832_ _03848_ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__clkbuf_1
X_18620_ clknet_leaf_15_clk _02049_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[113\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_217_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _03812_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__clkbuf_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ clknet_leaf_78_clk _01980_ net580 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[78\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_204_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12975_ fifo_bank_register.bank\[1\]\[18\] _05307_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07792_ sky130_fd_sc_hd__mux2_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _05104_ _04927_ _05196_ _03018_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a31o_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17502_ net485 _00945_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _07238_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__clkbuf_1
X_18482_ clknet_leaf_57_clk _01911_ net602 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_15694_ _03776_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ net560 _00876_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14645_ _02960_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__clkbuf_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11857_ fifo_bank_register.bank\[5\]\[2\] _05274_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07202_ sky130_fd_sc_hd__mux2_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17364_ net534 _00807_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_10808_ _06563_ vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__clkbuf_1
X_14576_ fifo_bank_register.bank\[1\]\[112\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[112\]
+ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__a22o_1
X_11788_ fifo_bank_register.bank\[6\]\[98\] _05476_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16315_ net680 _04136_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13527_ _05262_ fifo_bank_register.read_ptr\[3\] fifo_bank_register.read_ptr\[0\]
+ fifo_bank_register.read_ptr\[1\] vssd1 vssd1 vccd1 vccd1 _08098_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_166_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17295_ net543 _00738_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
X_10739_ _06500_ vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16246_ _04869_ _04189_ _04371_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__a21o_1
XFILLER_0_179_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13458_ _08046_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12409_ _07493_ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16177_ _04112_ _04124_ _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__and3_1
X_13389_ _08010_ vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15128_ _03395_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_220_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15059_ sub1.data_o\[28\] _04379_ _03059_ _03330_ vssd1 vssd1 vccd1 vccd1 _03331_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_177_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09620_ net146 vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__buf_2
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09551_ _05463_ vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_179_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08502_ addroundkey_data_o\[90\] fifo_bank_register.data_out\[90\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09482_ _05416_ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08433_ _04532_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08364_ _04496_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08295_ net234 net236 net237 net233 vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09818_ _05669_ _05670_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__xor2_1
Xfanout398 net404 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__buf_2
X_09749_ _05607_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12760_ fifo_bank_register.bank\[2\]\[44\] _05363_ _07674_ vssd1 vssd1 vccd1 vccd1
+ _07679_ sky130_fd_sc_hd__mux2_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11711_ fifo_bank_register.bank\[6\]\[61\] _05399_ _07123_ vssd1 vssd1 vccd1 vccd1
+ _07125_ sky130_fd_sc_hd__mux2_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _07642_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_182_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _02769_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11642_ _07088_ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__clkbuf_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14361_ fifo_bank_register.bank\[1\]\[89\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[89\]
+ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ fifo_bank_register.bank\[7\]\[125\] _05532_ _06912_ vssd1 vssd1 vccd1 vccd1
+ _07051_ sky130_fd_sc_hd__mux2_1
Xinput18 data_i[115] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_4
X_16100_ ks1.key_reg\[17\] _04057_ _03958_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13312_ _05373_ fifo_bank_register.bank\[0\]\[49\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 data_i[125] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__buf_4
X_17080_ net407 _00523_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
X_10524_ net232 ks1.key_reg\[77\] _06245_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14292_ fifo_bank_register.bank\[5\]\[81\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[81\]
+ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16031_ net229 ks1.key_reg\[74\] _03907_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13243_ _07933_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10455_ _05707_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13174_ fifo_bank_register.bank\[1\]\[112\] _05506_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07897_ sky130_fd_sc_hd__mux2_1
X_10386_ net215 ks1.key_reg\[61\] _06166_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12125_ _07343_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17982_ net472 _01425_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16933_ net402 _00376_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
X_12056_ _07306_ vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _06740_ _06741_ vssd1 vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__xor2_1
X_16864_ net483 _00307_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_204_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18603_ clknet_leaf_13_clk _02032_ net628 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15815_ _03839_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__clkbuf_1
X_16795_ clknet_leaf_73_clk _00239_ net590 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[86\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_204_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15746_ _03803_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__clkbuf_1
X_18534_ clknet_leaf_61_clk _01963_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ _07771_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__buf_4
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11909_ _07229_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__clkbuf_1
X_15677_ _03767_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__clkbuf_1
X_18465_ clknet_leaf_83_clk _01895_ net584 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[105\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _07746_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_270 _05977_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_281 fifo_bank_register.data_out\[116\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_292 sub1.data_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17416_ net524 _00859_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
X_14628_ _02945_ fifo_bank_register.data_out\[118\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _02946_ sky130_fd_sc_hd__mux2_1
X_18396_ clknet_leaf_19_clk _01826_ net640 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[81\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17347_ net494 _00790_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14559_ fifo_bank_register.bank\[1\]\[110\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[110\]
+ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17278_ net570 _00721_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16229_ _04173_ _04174_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_140_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08982_ ks1.key_reg\[7\] _04729_ _04731_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__or3_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09603_ _05498_ vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_196_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09534_ fifo_bank_register.bank\[9\]\[86\] _05451_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_223_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ net218 vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08416_ addroundkey_data_o\[49\] fifo_bank_register.data_out\[49\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09396_ _05358_ vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08347_ _04487_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _04427_ _04428_ _04429_ _04434_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__or4_4
XFILLER_0_225_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10240_ _05899_ _06046_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_225_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ _05603_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__buf_4
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13930_ fifo_bank_register.bank\[6\]\[41\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[41\]
+ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13861_ fifo_bank_register.bank\[5\]\[34\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[34\]
+ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15600_ mix1.data_o\[6\] _03392_ mix1.next_ready_o vssd1 vssd1 vccd1 vccd1 _03726_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12812_ fifo_bank_register.bank\[2\]\[69\] _05415_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_198_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16580_ net512 _00028_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13792_ _02201_ fifo_bank_register.data_out\[26\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15531_ sub1.data_o\[58\] _05559_ _04884_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__mux2_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ fifo_bank_register.bank\[2\]\[36\] _05346_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18250_ clknet_leaf_21_clk _01681_ net643 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ sub1.data_o\[66\] _05559_ _03633_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__mux2_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _07633_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ net451 _00644_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
X_14413_ _02754_ fifo_bank_register.data_out\[94\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18181_ clknet_leaf_1_clk _01612_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[75\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ fifo_bank_register.bank\[6\]\[20\] _05311_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07080_ sky130_fd_sc_hd__mux2_1
X_15393_ _03019_ _03593_ _05548_ _03596_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17132_ net417 _00575_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14344_ fifo_bank_register.bank\[9\]\[87\] _02631_ _02690_ _02691_ _02692_ vssd1
+ vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__a2111o_1
X_11556_ _07042_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17063_ net402 _00506_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
X_10507_ net230 ks1.key_reg\[75\] _06245_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__mux2_1
X_14275_ _02136_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__clkbuf_4
X_11487_ _07006_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__clkbuf_1
X_16014_ _03978_ _03980_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__xor2_2
XFILLER_0_111_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13226_ _07924_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_204_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10438_ _06229_ vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ fifo_bank_register.bank\[1\]\[104\] _05489_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07888_ sky130_fd_sc_hd__mux2_1
X_10369_ _05792_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__buf_4
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _07333_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__clkbuf_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ fifo_bank_register.bank\[1\]\[71\] _05420_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07852_ sky130_fd_sc_hd__mux2_1
X_17965_ net467 _01408_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12039_ _07297_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16916_ net525 _00359_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17896_ net431 _01339_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16847_ net426 _00290_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16778_ clknet_leaf_79_clk _00222_ net579 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[69\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_220_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18517_ clknet_leaf_63_clk _01946_ net599 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_15729_ _03794_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_158_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09250_ fifo_bank_register.write_ptr\[3\] vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__inv_2
X_18448_ clknet_leaf_74_clk _01878_ net593 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[88\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09181_ _05184_ _05191_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__xor2_2
XFILLER_0_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18379_ clknet_3_3__leaf_clk _01809_ net635 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[64\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_6109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08965_ addroundkey_data_o\[103\] _04666_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__or2_1
Xinput208 key_i[55] vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
XFILLER_0_228_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput219 key_i[65] vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_2
XFILLER_0_215_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08896_ ks1.key_reg\[0\] _04725_ _04919_ net130 vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09517_ _05440_ vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _05393_ vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_164_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ fifo_bank_register.bank\[9\]\[36\] _05346_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11410_ fifo_bank_register.bank\[7\]\[47\] _05369_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12390_ _05536_ fifo_bank_register.bank\[4\]\[127\] _07341_ vssd1 vssd1 vccd1 vccd1
+ _07482_ sky130_fd_sc_hd__mux2_1
X_11341_ _06929_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14060_ fifo_bank_register.bank\[7\]\[56\] _02380_ _02389_ fifo_bank_register.bank\[2\]\[56\]
+ _02439_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11272_ _06892_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13011_ _07811_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10223_ _06034_ _06035_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__xor2_1
XFILLER_0_218_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10154_ _05949_ _05970_ _05973_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__a21o_1
XTAP_5920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14962_ mix1.data_reg\[65\] _03236_ _03171_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__mux2_1
X_17750_ net497 _01193_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
X_10085_ _05910_ vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__clkbuf_1
Xhold7 ks1.key_reg\[40\] vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16701_ clknet_leaf_44_clk next_state net653 vssd1 vssd1 vccd1 vccd1 state sky130_fd_sc_hd__dfrtp_2
XTAP_5997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13913_ _02140_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__clkbuf_4
X_14893_ _03153_ _03168_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__xnor2_1
X_17681_ net544 _01124_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13844_ _02248_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__clkbuf_1
X_16632_ net553 _00080_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_226_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16563_ net473 _00011_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_13775_ fifo_bank_register.bank\[0\]\[24\] _02186_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02187_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10987_ sub1.data_o\[122\] _06723_ _06573_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__mux2_1
X_18302_ clknet_leaf_32_clk _01733_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[68\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15514_ _03668_ _04777_ _05196_ _03674_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__a31o_1
XFILLER_0_167_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12726_ fifo_bank_register.bank\[2\]\[28\] _05329_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16494_ _04330_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15445_ sub1.data_o\[28\] _05218_ _04879_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__mux2_1
X_18233_ clknet_leaf_11_clk _01664_ net622 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[63\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12657_ _07623_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ _07070_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__clkbuf_1
X_15376_ _03584_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18164_ clknet_leaf_82_clk _01595_ net587 vssd1 vssd1 vccd1 vccd1 ks1.col\[18\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_182_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12588_ fifo_bank_register.bank\[3\]\[91\] _05462_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14327_ fifo_bank_register.bank\[1\]\[85\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[85\]
+ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
X_17115_ net484 _00558_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18095_ net457 _01538_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[97\]
+ sky130_fd_sc_hd__dfxtp_1
X_11539_ _07033_ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17046_ net541 _00489_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14258_ fifo_bank_register.bank\[5\]\[78\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[78\]
+ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ _05248_ fifo_bank_register.bank\[0\]\[0\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14189_ fifo_bank_register.bank\[7\]\[70\] _02542_ _02551_ fifo_bank_register.bank\[2\]\[70\]
+ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a221o_1
XFILLER_0_209_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08750_ mix1.data_o\[25\] _04675_ _04670_ mix1.data_o\[49\] vssd1 vssd1 vccd1 vccd1
+ _04774_ sky130_fd_sc_hd__a22o_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ net538 _01391_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08681_ _04362_ _04673_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17879_ net532 _01322_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_221_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_215_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09302_ _05294_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _05193_ _05224_ _05060_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09164_ _05111_ _05173_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__and3_2
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09095_ _05105_ sbox1.inversion_to_invert_var\[3\] sbox1.inversion_to_invert_var\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_222_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ mix1.data_o\[24\] _05797_ _05821_ _05822_ sub1.data_o\[24\] vssd1 vssd1 vccd1
+ vccd1 _05832_ sky130_fd_sc_hd__a32o_1
XTAP_5227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_177_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ addroundkey_data_o\[127\] mix1.data_o\[127\] _04658_ vssd1 vssd1 vccd1 vccd1
+ _04972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ addroundkey_data_o\[104\] mix1.data_o\[104\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04903_ sky130_fd_sc_hd__mux2_1
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10910_ _05623_ _06650_ _06654_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_157_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11890_ fifo_bank_register.bank\[5\]\[18\] _05307_ _07210_ vssd1 vssd1 vccd1 vccd1
+ _07219_ sky130_fd_sc_hd__mux2_1
X_10841_ sub1.data_o\[107\] _06592_ _06573_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ _08129_ fifo_bank_register.data_out\[1\] _08064_ vssd1 vssd1 vccd1 vccd1
+ _08130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ net131 ks1.key_reg\[100\] _06402_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12511_ _07547_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ fifo_bank_register.read_ptr\[0\] fifo_bank_register.read_ptr\[1\] vssd1 vssd1
+ vccd1 vccd1 _08069_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15230_ _03281_ _03288_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12442_ _07511_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15161_ _03089_ _03410_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12373_ _07473_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14112_ fifo_bank_register.bank\[6\]\[61\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[61\]
+ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_205_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ _06920_ vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15092_ mix1.data_reg\[68\] _03363_ _03171_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_160_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14043_ fifo_bank_register.bank\[5\]\[54\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[54\]
+ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__a22o_1
X_11255_ _06883_ vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__clkbuf_1
X_10206_ net196 ks1.key_reg\[44\] _05997_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__mux2_1
X_11186_ _06791_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__buf_4
XFILLER_0_207_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17802_ net511 _01245_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_175_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10137_ _05958_ vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__clkbuf_1
XTAP_5750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15994_ _03961_ _03962_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__xor2_4
XTAP_5761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17733_ net441 _01176_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
X_10068_ _05568_ _05890_ _05894_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__o21ai_4
X_14945_ sub1.data_o\[9\] _04377_ _03081_ _03219_ vssd1 vssd1 vccd1 vccd1 _03220_
+ sky130_fd_sc_hd__a211o_1
XTAP_5794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17664_ net557 _01107_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_14876_ _03148_ _03151_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__nor2_8
XFILLER_0_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16615_ net572 _00063_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13827_ _02148_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__clkbuf_4
X_17595_ net432 _01038_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[117\]
+ sky130_fd_sc_hd__dfxtp_1
X_16546_ sub1.data_o\[81\] sub1.data_o\[17\] _03574_ vssd1 vssd1 vccd1 vccd1 _04358_
+ sky130_fd_sc_hd__mux2_1
X_13758_ fifo_bank_register.bank\[9\]\[22\] _02137_ _02169_ _02170_ _02171_ vssd1
+ vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_169_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12709_ _07651_ vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16477_ net739 _03170_ _04321_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__mux2_1
X_13689_ fifo_bank_register.bank\[1\]\[16\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18216_ clknet_leaf_84_clk _01647_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15428_ sub1.data_o\[117\] sub1.data_o\[53\] _03609_ vssd1 vssd1 vccd1 vccd1 _03619_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15359_ _03572_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__clkbuf_1
X_18147_ clknet_leaf_78_clk _01578_ net579 vssd1 vssd1 vccd1 vccd1 ks1.col\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_171_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18078_ net566 _01521_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[80\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09920_ net165 ks1.key_reg\[16\] _05762_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__mux2_4
XFILLER_0_180_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17029_ net524 _00472_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09851_ net12 mix1.data_o\[10\] _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ addroundkey_data_o\[35\] mix1.data_o\[35\] _04805_ vssd1 vssd1 vccd1 vccd1
+ _04826_ sky130_fd_sc_hd__mux2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ sub1.data_o\[2\] _05638_ _05610_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__mux2_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ ks1.key_reg\[9\] _04742_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08664_ _04364_ _04365_ _04687_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__and3_1
XFILLER_0_178_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08595_ _04615_ _04621_ _04617_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ _05215_ _05224_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_118_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_161_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09147_ sbox1.ah_reg\[3\] _05119_ _05157_ _05155_ vssd1 vssd1 vccd1 vccd1 _05158_
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09078_ sbox1.ah\[0\] vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11040_ _06770_ vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ fifo_bank_register.bank\[1\]\[25\] _05323_ _07795_ vssd1 vssd1 vccd1 vccd1
+ _07801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11942_ fifo_bank_register.bank\[5\]\[42\] _05359_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07247_ sky130_fd_sc_hd__mux2_1
X_14730_ ks1.col\[1\] _05553_ _04916_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _02974_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11873_ _07198_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__buf_4
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13612_ fifo_bank_register.bank\[7\]\[8\] _08078_ _08093_ fifo_bank_register.bank\[2\]\[8\]
+ _08174_ vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__a221o_1
X_16400_ _04279_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__clkbuf_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _06416_ _06574_ _06577_ _06420_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ net430 _00823_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_14592_ fifo_bank_register.bank\[1\]\[114\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[114\]
+ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a22o_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13543_ _08113_ vssd1 vssd1 vccd1 vccd1 _08114_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16331_ net838 _03920_ _04240_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ _06395_ _06514_ sub1.data_o\[99\] _06384_ vssd1 vssd1 vccd1 vccd1 _06515_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_153_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16262_ _04203_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__clkbuf_1
X_13474_ _08054_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_180_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10686_ addroundkey_data_o\[92\] _06452_ _06431_ vssd1 vssd1 vccd1 vccd1 _06453_
+ sky130_fd_sc_hd__mux2_1
X_15213_ _03473_ _03474_ _05198_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__a21o_2
XFILLER_0_152_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18001_ net420 _01444_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12425_ fifo_bank_register.bank\[3\]\[14\] _05299_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07502_ sky130_fd_sc_hd__mux2_1
X_16193_ ks1.col\[26\] _04141_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15144_ net769 _03411_ _03171_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12356_ _05501_ fifo_bank_register.bank\[4\]\[110\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput309 net309 vssd1 vssd1 vccd1 vccd1 data_o[29] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_168_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11307_ fifo_bank_register.write_ptr\[2\] _05254_ _05266_ vssd1 vssd1 vccd1 vccd1
+ _06910_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15075_ sub1.data_o\[3\] _04378_ _03059_ _03346_ vssd1 vssd1 vccd1 vccd1 _03347_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12287_ _07428_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__clkbuf_1
X_14026_ _02410_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11238_ _06874_ vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11169_ _06838_ vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15977_ _04734_ _03947_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__xnor2_1
XTAP_5591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17716_ net434 _01159_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[110\]
+ sky130_fd_sc_hd__dfxtp_1
X_14928_ sub1.data_o\[121\] _03056_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17647_ net398 _01090_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
X_14859_ addroundkey_data_o\[93\] _03108_ _03066_ addroundkey_data_o\[61\] vssd1 vssd1
+ vccd1 vccd1 _03135_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ addroundkey_data_o\[32\] fifo_bank_register.data_out\[32\] _04501_ vssd1
+ vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__mux2_1
X_17578_ net447 _01021_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16529_ net757 _03516_ _04343_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09001_ _04670_ _05021_ _05022_ _04675_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09903_ _05745_ _05746_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout503 net504 vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
Xfanout514 net520 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__buf_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout525 net526 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__buf_2
Xfanout536 net537 vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_2
X_09834_ mix1.data_o\[8\] _05677_ _05618_ _05621_ sub1.data_o\[8\] vssd1 vssd1 vccd1
+ vccd1 _05685_ sky130_fd_sc_hd__a32o_1
Xfanout547 net551 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__buf_2
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout558 net559 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout569 net577 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_214_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09765_ _05611_ _05615_ _05622_ _05623_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__a22o_2
XFILLER_0_119_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_197_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08716_ ks1.state\[1\] ks1.state\[2\] ks1.state\[0\] vssd1 vssd1 vccd1 vccd1 _04740_
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_55_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09696_ _05563_ vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08647_ addroundkey_data_o\[52\] mix1.data_o\[52\] _04663_ vssd1 vssd1 vccd1 vccd1
+ _04671_ sky130_fd_sc_hd__mux2_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08578_ addroundkey_data_o\[127\] fifo_bank_register.data_out\[127\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__mux2_2
XFILLER_0_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10540_ _05757_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10471_ net97 mix1.data_o\[71\] _06237_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_162_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12210_ _07388_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13190_ fifo_bank_register.bank\[1\]\[120\] _05522_ _07771_ vssd1 vssd1 vccd1 vccd1
+ _07905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_161_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ _07351_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12072_ fifo_bank_register.bank\[5\]\[104\] _05489_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15900_ _05227_ sub1.data_o\[69\] _05199_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__mux2_1
X_11023_ _06754_ _06755_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__xor2_1
XFILLER_0_194_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16880_ net405 _00323_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_198_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_217_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15831_ mix1.data_o\[115\] net696 _03841_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__mux2_1
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18550_ clknet_leaf_64_clk _01979_ net603 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[77\]
+ sky130_fd_sc_hd__dfrtp_1
X_15762_ mix1.data_o\[82\] net748 _03808_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__mux2_1
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ _07791_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__clkbuf_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ net487 _00944_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14713_ sub1.data_o\[83\] _03010_ _03017_ sub1.next_ready_o vssd1 vssd1 vccd1 vccd1
+ _03018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ fifo_bank_register.bank\[5\]\[34\] _05342_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07238_ sky130_fd_sc_hd__mux2_1
X_18481_ clknet_leaf_59_clk _01910_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_15693_ mix1.data_o\[49\] net788 _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__mux2_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ net560 _00875_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11856_ _07201_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14644_ _02959_ fifo_bank_register.data_out\[120\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _02960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10807_ addroundkey_data_o\[103\] _06562_ _06522_ vssd1 vssd1 vccd1 vccd1 _06563_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17363_ net505 _00806_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14575_ fifo_bank_register.bank\[6\]\[112\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[112\]
+ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11787_ _07164_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__clkbuf_1
X_16314_ _04215_ _04134_ _04231_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__o21ai_1
X_13526_ _08096_ vssd1 vssd1 vccd1 vccd1 _08097_ sky130_fd_sc_hd__clkbuf_4
X_10738_ addroundkey_data_o\[97\] _06499_ _06431_ vssd1 vssd1 vccd1 vccd1 _06500_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17294_ net544 _00737_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13457_ _05518_ fifo_bank_register.bank\[0\]\[118\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08046_ sky130_fd_sc_hd__mux2_1
X_16245_ _04869_ _04189_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__nor2_1
X_10669_ _06436_ _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__xor2_1
XFILLER_0_179_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12408_ fifo_bank_register.bank\[3\]\[6\] _05282_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13388_ _05449_ fifo_bank_register.bank\[0\]\[85\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08010_ sky130_fd_sc_hd__mux2_1
X_16176_ _04113_ _04125_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15127_ _03343_ _03361_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_121_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12339_ _05485_ fifo_bank_register.bank\[4\]\[102\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15058_ sub1.data_o\[92\] _03144_ _03145_ sub1.data_o\[60\] vssd1 vssd1 vccd1 vccd1
+ _03330_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14009_ _02148_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09550_ fifo_bank_register.bank\[9\]\[91\] _05462_ _05460_ vssd1 vssd1 vccd1 vccd1
+ _05463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08501_ _04568_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_2
X_09481_ fifo_bank_register.bank\[9\]\[69\] _05415_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ addroundkey_data_o\[57\] fifo_bank_register.data_out\[57\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__mux2_2
XFILLER_0_153_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08363_ addroundkey_data_o\[24\] fifo_bank_register.data_out\[24\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08294_ net226 net228 net227 net225 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_50_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09817_ net224 ks1.key_reg\[6\] _05625_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout399 net404 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_213_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09748_ _05606_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _05154_ _05243_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__nor2_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _07124_ vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__clkbuf_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12690_ fifo_bank_register.bank\[2\]\[11\] _05293_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07642_ sky130_fd_sc_hd__mux2_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11641_ fifo_bank_register.bank\[6\]\[28\] _05329_ _07079_ vssd1 vssd1 vccd1 vccd1
+ _07088_ sky130_fd_sc_hd__mux2_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_181_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14360_ fifo_bank_register.bank\[6\]\[89\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[89\]
+ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a22o_1
X_11572_ _07050_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _07969_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10523_ _06250_ _06303_ _06304_ _06254_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__a22o_1
Xinput19 data_i[116] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14291_ _02646_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13242_ _05303_ fifo_bank_register.bank\[0\]\[16\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07933_ sky130_fd_sc_hd__mux2_1
X_16030_ net194 ks1.key_reg\[42\] _03910_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10454_ _06171_ _06240_ _06243_ _06175_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__a22o_2
XFILLER_0_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13173_ _07896_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__clkbuf_1
X_10385_ _06171_ _06181_ _06182_ _06175_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12124_ _05248_ fifo_bank_register.bank\[4\]\[0\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17981_ net435 _01424_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12055_ fifo_bank_register.bank\[5\]\[96\] _05472_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07306_ sky130_fd_sc_hd__mux2_1
X_16932_ net454 _00375_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
X_11006_ net157 ks1.key_reg\[124\] _05762_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16863_ net488 _00306_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_18602_ clknet_leaf_14_clk _02031_ net629 vssd1 vssd1 vccd1 vccd1 mix1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_15814_ mix1.data_o\[107\] net746 _03830_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_204_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16794_ clknet_leaf_39_clk _00238_ net663 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[85\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18533_ clknet_leaf_61_clk _01962_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
X_15745_ mix1.data_o\[74\] net727 _03797_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__mux2_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _07782_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18464_ clknet_leaf_3_clk _01894_ net583 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[104\]
+ sky130_fd_sc_hd__dfrtp_4
X_11908_ fifo_bank_register.bank\[5\]\[26\] _05325_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07229_ sky130_fd_sc_hd__mux2_1
X_15676_ mix1.data_o\[41\] net754 _03764_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_260 net266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ fifo_bank_register.bank\[2\]\[105\] _05491_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07746_ sky130_fd_sc_hd__mux2_1
XANTENNA_271 addroundkey_data_o\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17415_ net518 _00858_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_282 fifo_bank_register.data_out\[116\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_293 sub1.data_o\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14627_ fifo_bank_register.bank\[0\]\[118\] _02944_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02945_ sky130_fd_sc_hd__mux2_1
X_18395_ clknet_leaf_18_clk _01825_ net638 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[80\]
+ sky130_fd_sc_hd__dfrtp_4
X_11839_ _07191_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17346_ net494 _00789_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14558_ _02153_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13509_ _05250_ _08082_ _05266_ vssd1 vssd1 vccd1 vccd1 _08083_ sky130_fd_sc_hd__mux2_1
X_17277_ net570 _00720_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14489_ _02822_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16228_ net158 ks1.key_reg\[125\] _03976_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__mux2_2
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16159_ _04644_ _05539_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08981_ ks1.key_reg\[15\] _04726_ _05004_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_228_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09602_ fifo_bank_register.bank\[9\]\[108\] _05497_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09533_ net242 vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_211_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09464_ _05404_ vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08415_ _04478_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__buf_12
X_09395_ fifo_bank_register.bank\[9\]\[41\] _05357_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08346_ addroundkey_data_o\[16\] fifo_bank_register.data_out\[16\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__mux2_4
XFILLER_0_184_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08277_ _04430_ _04431_ _04432_ _04433_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__or4_1
XFILLER_0_190_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10170_ _05988_ vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13860_ _02262_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12811_ _07705_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13791_ fifo_bank_register.bank\[0\]\[26\] _02200_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15530_ _03684_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__clkbuf_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _07669_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_210_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_166_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _03639_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__clkbuf_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ fifo_bank_register.bank\[2\]\[3\] _05276_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ net465 _00643_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_182_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__buf_4
X_14412_ fifo_bank_register.bank\[0\]\[94\] _02753_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18180_ clknet_leaf_0_clk _01611_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[74\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15392_ sub1.data_o\[72\] _03594_ _03595_ sub1.data_o\[8\] vssd1 vssd1 vccd1 vccd1
+ _03596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17131_ net414 _00574_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
X_11555_ fifo_bank_register.bank\[7\]\[116\] _05514_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07042_ sky130_fd_sc_hd__mux2_1
X_14343_ fifo_bank_register.bank\[1\]\[87\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[87\]
+ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10506_ _06250_ _06288_ _06289_ _06254_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__a22o_1
X_14274_ _02630_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__clkbuf_1
X_17062_ net401 _00505_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11486_ fifo_bank_register.bank\[7\]\[83\] _05445_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13225_ _05286_ fifo_bank_register.bank\[0\]\[8\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07924_ sky130_fd_sc_hd__mux2_1
X_16013_ net227 ks1.key_reg\[72\] _03979_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__mux2_1
X_10437_ addroundkey_data_o\[67\] _06228_ _06169_ vssd1 vssd1 vccd1 vccd1 _06229_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13156_ _07887_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__clkbuf_1
X_10368_ _06165_ _06167_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__xor2_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ fifo_bank_register.bank\[5\]\[121\] _05524_ _07198_ vssd1 vssd1 vccd1 vccd1
+ _07333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _07851_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__clkbuf_1
X_17964_ net466 _01407_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
X_10299_ mix1.data_o\[53\] _05952_ _06093_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__o21a_1
XFILLER_0_224_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_178_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12038_ fifo_bank_register.bank\[5\]\[88\] _05455_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07297_ sky130_fd_sc_hd__mux2_1
X_16915_ net553 _00358_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_218_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17895_ net425 _01338_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16846_ net425 _00289_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16777_ clknet_leaf_48_clk _00221_ net611 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[68\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13989_ fifo_bank_register.bank\[9\]\[48\] _02307_ _02374_ _02375_ _02376_ vssd1
+ vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a2111o_1
X_18516_ clknet_leaf_62_clk _01945_ net599 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15728_ mix1.data_o\[66\] mix1.data_reg\[66\] _03786_ vssd1 vssd1 vccd1 vccd1 _03794_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_186_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18447_ clknet_leaf_9_clk _01877_ net631 vssd1 vssd1 vccd1 vccd1 sub1.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15659_ mix1.data_o\[33\] net772 _03753_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09180_ _05187_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18378_ clknet_leaf_46_clk _01808_ net652 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[63\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17329_ net462 _00772_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput209 key_i[56] vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_4
X_08964_ _04986_ _04987_ _04698_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__mux2_1
XFILLER_0_227_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08895_ ks1.key_reg\[0\] _04729_ _04731_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__or3_1
XFILLER_0_192_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_918 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09516_ fifo_bank_register.bank\[9\]\[80\] _05438_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_182_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09447_ fifo_bank_register.bank\[9\]\[58\] _05392_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05393_ sky130_fd_sc_hd__mux2_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_176_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09378_ net187 vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08329_ _04477_ vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_2
XFILLER_0_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ fifo_bank_register.bank\[7\]\[14\] _05299_ _06924_ vssd1 vssd1 vccd1 vccd1
+ _06929_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11271_ _05501_ fifo_bank_register.bank\[8\]\[110\] _06891_ vssd1 vssd1 vccd1 vccd1
+ _06892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ fifo_bank_register.bank\[1\]\[34\] _05342_ _07806_ vssd1 vssd1 vccd1 vccd1
+ _07811_ sky130_fd_sc_hd__mux2_1
X_10222_ net198 ks1.key_reg\[46\] _05997_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10153_ _05913_ _05972_ sub1.data_o\[39\] _05902_ vssd1 vssd1 vccd1 vccd1 _05973_
+ sky130_fd_sc_hd__a31o_1
XTAP_5910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14961_ _03200_ _03235_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__xnor2_2
X_10084_ addroundkey_data_o\[33\] _05909_ _05872_ vssd1 vssd1 vccd1 vccd1 _05910_
+ sky130_fd_sc_hd__mux2_1
XTAP_5954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 ks1.key_reg\[108\] vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16700_ clknet_leaf_71_clk _00147_ net652 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[127\]
+ sky130_fd_sc_hd__dfrtp_2
X_13912_ _02138_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__clkbuf_4
XTAP_5987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ net549 _01123_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14892_ _03160_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16631_ net528 _00079_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13843_ _02247_ fifo_bank_register.data_out\[31\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_199_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16562_ net474 _00010_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_10986_ net26 mix1.data_o\[122\] _06571_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__mux2_1
X_13774_ fifo_bank_register.bank\[9\]\[24\] _02137_ _02183_ _02184_ _02185_ vssd1
+ vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_69_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18301_ clknet_leaf_27_clk _01732_ net642 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[67\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15513_ sub1.data_o\[51\] _03663_ _03672_ _03673_ vssd1 vssd1 vccd1 vccd1 _03674_
+ sky130_fd_sc_hd__a22o_1
X_12725_ _07660_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__clkbuf_1
X_16493_ net781 _03411_ _04321_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18232_ clknet_leaf_9_clk _01663_ net631 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[62\]
+ sky130_fd_sc_hd__dfrtp_2
X_15444_ _03628_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12656_ fifo_bank_register.bank\[3\]\[124\] _05530_ _07485_ vssd1 vssd1 vccd1 vccd1
+ _07623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11607_ fifo_bank_register.bank\[6\]\[12\] _05295_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07070_ sky130_fd_sc_hd__mux2_1
X_18163_ clknet_leaf_76_clk _01594_ net589 vssd1 vssd1 vccd1 vccd1 ks1.col\[17\] sky130_fd_sc_hd__dfrtp_4
X_15375_ sub1.data_o\[3\] _03583_ _03581_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12587_ _07587_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17114_ net512 _00557_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
X_14326_ fifo_bank_register.bank\[6\]\[85\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[85\]
+ vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18094_ net398 _01537_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[96\]
+ sky130_fd_sc_hd__dfxtp_1
X_11538_ fifo_bank_register.bank\[7\]\[108\] _05497_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17045_ net547 _00488_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11469_ fifo_bank_register.bank\[7\]\[75\] _05428_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _06997_ sky130_fd_sc_hd__mux2_1
X_14257_ _02615_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13208_ _07914_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14188_ fifo_bank_register.bank\[5\]\[70\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[70\]
+ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__a22o_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13139_ _07878_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__clkbuf_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ net568 _01390_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08680_ mix1.data_o\[100\] _04698_ _04701_ _04703_ vssd1 vssd1 vccd1 vccd1 _04704_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17878_ net497 _01321_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16829_ clknet_leaf_74_clk _00273_ net591 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[120\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_221_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09301_ fifo_bank_register.bank\[9\]\[11\] _05293_ _05291_ vssd1 vssd1 vccd1 vccd1
+ _05294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_215_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09232_ _05193_ _05224_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09163_ sbox1.ah_reg\[3\] sbox1.ah_reg\[2\] vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09094_ sbox1.inversion_to_invert_var\[2\] vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__buf_2
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ sub1.data_o\[24\] _05830_ _05819_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__mux2_1
XTAP_5217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _04877_ _04970_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__xor2_4
XTAP_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08878_ mix1.data_o\[96\] _04900_ _04701_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_
+ sky130_fd_sc_hd__o211a_1
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_224_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10840_ net9 mix1.data_o\[107\] _06571_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10771_ _06381_ _06525_ _06529_ vssd1 vssd1 vccd1 vccd1 _06530_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12510_ fifo_bank_register.bank\[3\]\[54\] _05384_ _07542_ vssd1 vssd1 vccd1 vccd1
+ _07547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13490_ _08063_ vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_165_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ fifo_bank_register.bank\[3\]\[21\] _05315_ _07509_ vssd1 vssd1 vccd1 vccd1
+ _07511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15160_ _03426_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12372_ _05518_ fifo_bank_register.bank\[4\]\[118\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11323_ fifo_bank_register.bank\[7\]\[6\] _05282_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06920_ sky130_fd_sc_hd__mux2_1
X_14111_ fifo_bank_register.bank\[7\]\[61\] _02461_ _02470_ fifo_bank_register.bank\[2\]\[61\]
+ _02485_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a221o_1
X_15091_ _03345_ _03362_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_26_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14042_ _02424_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__clkbuf_1
X_11254_ _05485_ fifo_bank_register.bank\[8\]\[102\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_205_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10205_ _06001_ _06018_ _06019_ _06005_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11185_ _06846_ vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17801_ net511 _01244_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
X_10136_ addroundkey_data_o\[37\] _05957_ _05872_ vssd1 vssd1 vccd1 vccd1 _05958_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15993_ net225 ks1.key_reg\[70\] _03907_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__mux2_2
XTAP_5751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17732_ net494 _01175_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10067_ sub1.data_o\[32\] _05753_ _05892_ _05893_ _04611_ vssd1 vssd1 vccd1 vccd1
+ _05894_ sky130_fd_sc_hd__a221o_1
X_14944_ sub1.data_o\[73\] _03063_ _03092_ sub1.data_o\[41\] vssd1 vssd1 vccd1 vccd1
+ _03219_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17663_ net550 _01106_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14875_ addroundkey_data_o\[104\] _03143_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_202_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16614_ net556 _00062_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13826_ _02146_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17594_ net409 _01037_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16545_ _05103_ _04946_ _05548_ _04357_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ fifo_bank_register.bank\[1\]\[22\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__a22o_1
X_10969_ _06708_ vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12708_ _07627_ vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__buf_6
X_16476_ _03143_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__buf_4
XFILLER_0_31_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13688_ fifo_bank_register.bank\[6\]\[16\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18215_ clknet_leaf_84_clk _01646_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[45\]
+ sky130_fd_sc_hd__dfrtp_1
X_15427_ _03603_ _04949_ _05219_ _03618_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ _07614_ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_208_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18146_ clknet_leaf_64_clk _01577_ net603 vssd1 vssd1 vccd1 vccd1 ks1.col\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ mix1.data_reg\[62\] _03533_ _03145_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14309_ fifo_bank_register.bank\[7\]\[83\] _02623_ _02632_ fifo_bank_register.bank\[2\]\[83\]
+ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__a221o_1
X_18077_ net568 _01520_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_223_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15289_ _03534_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17028_ net523 _00471_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09850_ _05603_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__buf_4
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08801_ _04701_ _04823_ _04824_ _04682_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__a22o_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ net51 mix1.data_o\[2\] _05604_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__mux2_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ ks1.key_reg\[9\] _04730_ _04732_ net257 vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__o31a_1
X_08663_ sub1.state\[1\] sub1.state\[0\] vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__and2_1
XFILLER_0_205_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08594_ round\[1\] round\[2\] round\[3\] _04613_ vssd1 vssd1 vccd1 vccd1 _04621_
+ sky130_fd_sc_hd__and4bb_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09215_ _05212_ _05223_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09146_ sbox1.ah_reg\[0\] sbox1.ah_reg\[3\] vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09077_ _04877_ _05090_ vssd1 vssd1 vccd1 vccd1 sbox1.intermediate_to_invert_var\[2\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_228_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09979_ addroundkey_data_o\[22\] _05815_ _05793_ vssd1 vssd1 vccd1 vccd1 _05816_
+ sky130_fd_sc_hd__mux2_1
XTAP_5047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _07800_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__clkbuf_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _07246_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__clkbuf_1
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14660_ _02973_ fifo_bank_register.data_out\[122\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _02974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _07209_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ fifo_bank_register.bank\[5\]\[8\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[8\]
+ vssd1 vssd1 vccd1 vccd1 _08174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ mix1.data_o\[105\] _06463_ _06575_ _06576_ sub1.data_o\[105\] vssd1 vssd1
+ vccd1 vccd1 _06577_ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14591_ fifo_bank_register.bank\[6\]\[114\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[114\]
+ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a22o_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16330_ _04372_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ _08056_ _08070_ vssd1 vssd1 vccd1 vccd1 _08113_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10754_ sub1.ready_o vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16261_ net813 _03922_ _04106_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13473_ _05534_ fifo_bank_register.bank\[0\]\[126\] _07914_ vssd1 vssd1 vccd1 vccd1
+ _08054_ sky130_fd_sc_hd__mux2_1
X_10685_ _06450_ _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18000_ net420 _01443_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[2\] sky130_fd_sc_hd__dfxtp_1
X_15212_ _03455_ _03472_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__or2_1
X_12424_ _07501_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16192_ _04111_ _04138_ _04140_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__or3_2
XFILLER_0_106_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15143_ _03409_ _03410_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12355_ _07364_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__buf_4
XFILLER_0_11_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11306_ _06909_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15074_ sub1.data_o\[67\] _03064_ _03084_ sub1.data_o\[35\] vssd1 vssd1 vccd1 vccd1
+ _03346_ sky130_fd_sc_hd__a22o_1
X_12286_ _05432_ fifo_bank_register.bank\[4\]\[77\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14025_ _02409_ fifo_bank_register.data_out\[51\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02410_ sky130_fd_sc_hd__mux2_1
X_11237_ _05468_ fifo_bank_register.bank\[8\]\[94\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11168_ _05399_ fifo_bank_register.bank\[8\]\[61\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10119_ sub1.data_o\[36\] _05753_ _05939_ _05940_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _05942_ sky130_fd_sc_hd__a221o_1
XTAP_5570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ _06801_ vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__clkbuf_1
X_15976_ _03945_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__xor2_2
XTAP_5581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17715_ net458 _01158_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_188_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14927_ sub1.data_o\[25\] _04377_ _03081_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17646_ net397 _01089_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_14858_ sub1.data_o\[125\] _03055_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_37_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13809_ _02216_ fifo_bank_register.data_out\[28\] _02209_ vssd1 vssd1 vccd1 vccd1
+ _02217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_212_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17577_ net445 _01020_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ mix1.state\[0\] _03060_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__nor2_2
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16528_ _04348_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16459_ net682 _04373_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nor2_1
XFILLER_0_186_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09000_ addroundkey_data_o\[26\] mix1.data_o\[26\] _04803_ vssd1 vssd1 vccd1 vccd1
+ _05022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18129_ clknet_leaf_24_clk _01572_ net643 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[83\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09902_ net164 ks1.key_reg\[15\] _05708_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout504 net507 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__buf_2
XFILLER_0_1_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout515 net520 vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout526 net528 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_2
X_09833_ sub1.data_o\[8\] _05683_ _05610_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__mux2_1
Xfanout537 net577 vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_2
Xfanout548 net551 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout559 net577 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09764_ _04609_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__buf_6
XFILLER_0_213_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08715_ _04721_ _04734_ _04736_ _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_213_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09695_ sub1.data_o\[124\] _05219_ _04891_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ sub1.state\[1\] sub1.state\[2\] sub1.state\[3\] _04363_ vssd1 vssd1 vccd1
+ vccd1 _04670_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _04607_ vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10470_ _06258_ vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09129_ _05138_ _05139_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__xor2_2
XFILLER_0_126_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12140_ _05286_ fifo_bank_register.bank\[4\]\[8\] _07342_ vssd1 vssd1 vccd1 vccd1
+ _07351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ _07314_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11022_ net159 ks1.key_reg\[126\] _05762_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15830_ _03847_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__clkbuf_1
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _03811_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__clkbuf_1
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ fifo_bank_register.bank\[1\]\[17\] _05305_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07791_ sky130_fd_sc_hd__mux2_1
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ net488 _00943_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_14712_ sub1.data_o\[51\] sub1.data_o\[115\] _05598_ vssd1 vssd1 vccd1 vccd1 _03017_
+ sky130_fd_sc_hd__mux2_1
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _07237_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__clkbuf_1
X_18480_ clknet_leaf_59_clk _01909_ net613 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_15692_ _03741_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__buf_4
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ net565 _00874_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
X_14643_ fifo_bank_register.bank\[0\]\[120\] _02958_ _08120_ vssd1 vssd1 vccd1 vccd1
+ _02959_ sky130_fd_sc_hd__mux2_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11855_ fifo_bank_register.bank\[5\]\[1\] _05272_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07201_ sky130_fd_sc_hd__mux2_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17362_ net504 _00805_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_10806_ _06560_ _06561_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14574_ fifo_bank_register.bank\[7\]\[112\] _02866_ _02875_ fifo_bank_register.bank\[2\]\[112\]
+ _02897_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a221o_1
X_11786_ fifo_bank_register.bank\[6\]\[97\] _05474_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_172_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16313_ net673 _04136_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13525_ _08095_ vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__clkbuf_4
X_17293_ net517 _00736_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[71\]
+ sky130_fd_sc_hd__dfxtp_1
X_10737_ _06497_ _06498_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_165_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16244_ _04187_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__xor2_2
X_13456_ _08045_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__clkbuf_1
X_10668_ net247 ks1.key_reg\[90\] _06324_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12407_ _07492_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16175_ addroundkey_round\[3\] _04642_ _04644_ _05544_ vssd1 vssd1 vccd1 vccd1 _04125_
+ sky130_fd_sc_hd__a31oi_4
X_10599_ _06126_ _06372_ _06373_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__a21o_1
X_13387_ _08009_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15126_ _03115_ _03131_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_51_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _07455_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15057_ _03199_ _03327_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__a21o_1
X_12269_ _05415_ fifo_bank_register.bank\[4\]\[69\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14008_ _02146_ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__buf_4
XFILLER_0_49_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15959_ _05050_ _03930_ _03914_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_211_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08500_ addroundkey_data_o\[89\] fifo_bank_register.data_out\[89\] _04567_ vssd1
+ vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__mux2_2
XFILLER_0_204_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09480_ net223 vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_210_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08431_ _04531_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_187_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17629_ net487 _01072_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ _04495_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08293_ net230 net229 net232 net231 vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__or4_1
XFILLER_0_160_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09816_ _05629_ _05667_ _05668_ _05633_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a22o_1
Xfanout389 net391 vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_2
XFILLER_0_214_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09747_ _04900_ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09678_ _05549_ vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ sub1.state\[4\] _04366_ _04652_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__and3b_4
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _07087_ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11571_ fifo_bank_register.bank\[7\]\[124\] _05530_ _06912_ vssd1 vssd1 vccd1 vccd1
+ _07050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13310_ _05371_ fifo_bank_register.bank\[0\]\[48\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10522_ mix1.data_o\[77\] _06296_ _06241_ _06242_ sub1.data_o\[77\] vssd1 vssd1 vccd1
+ vccd1 _06304_ sky130_fd_sc_hd__a32o_1
X_14290_ _02645_ fifo_bank_register.data_out\[80\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_162_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_190_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10453_ mix1.data_o\[69\] _06217_ _06241_ _06242_ sub1.data_o\[69\] vssd1 vssd1 vccd1
+ vccd1 _06243_ sky130_fd_sc_hd__a32o_1
X_13241_ _07932_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10384_ mix1.data_o\[61\] _06138_ _06162_ _06163_ sub1.data_o\[61\] vssd1 vssd1 vccd1
+ vccd1 _06182_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13172_ fifo_bank_register.bank\[1\]\[111\] _05504_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12123_ _07341_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17980_ net457 _01423_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
X_16931_ net400 _00374_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_12054_ _07305_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11005_ _05615_ _06738_ _06739_ _05567_ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__a22o_1
X_16862_ net482 _00305_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[24\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_217_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18601_ clknet_leaf_33_clk _02030_ net660 vssd1 vssd1 vccd1 vccd1 mix1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_15813_ _03838_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__clkbuf_1
X_16793_ clknet_leaf_73_clk _00237_ net593 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[84\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18532_ clknet_leaf_59_clk _01961_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[59\]
+ sky130_fd_sc_hd__dfrtp_1
X_15744_ _03802_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ fifo_bank_register.bank\[1\]\[9\] _05288_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18463_ clknet_leaf_34_clk _01893_ net662 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[103\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11907_ _07228_ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _03766_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_250 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ _07745_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__clkbuf_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_261 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17414_ net514 _00857_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_272 addroundkey_data_o\[112\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14626_ fifo_bank_register.bank\[9\]\[118\] _02874_ _02941_ _02942_ _02943_ vssd1
+ vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a2111o_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18394_ clknet_leaf_14_clk _01824_ net629 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[79\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_283 fifo_bank_register.data_out\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11838_ fifo_bank_register.bank\[6\]\[122\] _05526_ _07055_ vssd1 vssd1 vccd1 vccd1
+ _07191_ sky130_fd_sc_hd__mux2_1
XANTENNA_294 sub1.data_o\[22\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17345_ net439 _00788_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _02151_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__clkbuf_4
X_11769_ fifo_bank_register.bank\[6\]\[89\] _05457_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_clk clknet_3_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13508_ _05260_ vssd1 vssd1 vccd1 vccd1 _08082_ sky130_fd_sc_hd__inv_2
X_17276_ net555 _00719_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14488_ _02821_ fifo_bank_register.data_out\[102\] _02776_ vssd1 vssd1 vccd1 vccd1
+ _02822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16227_ ks1.col\[29\] _04172_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_148_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13439_ _08036_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16158_ _04727_ _04638_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15109_ _03115_ _03138_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16089_ _04046_ _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__xor2_2
X_08980_ ks1.key_reg\[15\] _04745_ _04746_ net164 vssd1 vssd1 vccd1 vccd1 _05004_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_227_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09601_ net139 vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__buf_2
XFILLER_0_194_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09532_ _05450_ vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ fifo_bank_register.bank\[9\]\[63\] _05403_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08414_ _04522_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__clkbuf_1
X_09394_ net193 vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08345_ _04486_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_188_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08276_ net255 net131 net132 net256 vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12810_ fifo_bank_register.bank\[2\]\[68\] _05413_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13790_ fifo_bank_register.bank\[9\]\[26\] _02137_ _02197_ _02198_ _02199_ vssd1
+ vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_186_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ fifo_bank_register.bank\[2\]\[35\] _05344_ _07663_ vssd1 vssd1 vccd1 vccd1
+ _07669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15460_ sub1.data_o\[33\] _03638_ _03636_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__mux2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12672_ _07632_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ fifo_bank_register.bank\[9\]\[94\] _02712_ _02750_ _02751_ _02752_ vssd1
+ vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__a2111o_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _07054_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__buf_8
XFILLER_0_93_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15391_ _03581_ _04689_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__nor2_2
XFILLER_0_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_16
X_17130_ net422 _00573_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14342_ fifo_bank_register.bank\[6\]\[87\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[87\]
+ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11554_ _07041_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ mix1.data_o\[75\] _06217_ _06241_ _06242_ sub1.data_o\[75\] vssd1 vssd1 vccd1
+ vccd1 _06289_ sky130_fd_sc_hd__a32o_1
X_17061_ net400 _00504_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
X_14273_ _02629_ fifo_bank_register.data_out\[79\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11485_ _07005_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _03905_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__buf_4
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13224_ _07923_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__clkbuf_1
X_10436_ _06226_ _06227_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13155_ fifo_bank_register.bank\[1\]\[103\] _05487_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10367_ net212 ks1.key_reg\[59\] _06166_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _07332_ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10298_ _05949_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__a21o_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ fifo_bank_register.bank\[1\]\[70\] _05417_ _07850_ vssd1 vssd1 vccd1 vccd1
+ _07851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17963_ net450 _01406_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16914_ net545 _00357_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
X_12037_ _07296_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17894_ net418 _01337_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16845_ net425 _00288_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16776_ clknet_leaf_48_clk _00220_ net610 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[67\]
+ sky130_fd_sc_hd__dfrtp_4
X_13988_ fifo_bank_register.bank\[1\]\[48\] _02316_ _02317_ fifo_bank_register.bank\[8\]\[48\]
+ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__a22o_1
XFILLER_0_220_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15727_ _03793_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18515_ clknet_leaf_65_clk _01944_ net604 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_12939_ _07773_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_220_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15658_ _03757_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__clkbuf_1
X_18446_ clknet_leaf_10_clk _01876_ net623 vssd1 vssd1 vccd1 vccd1 sub1.state\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14609_ fifo_bank_register.bank\[9\]\[116\] _02874_ _02926_ _02927_ _02928_ vssd1
+ vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_111_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18377_ clknet_3_6__leaf_clk _01807_ net653 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[62\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15589_ _03720_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_13_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17328_ net464 _00771_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17259_ net414 _00702_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08963_ addroundkey_data_o\[47\] _04693_ _04695_ addroundkey_data_o\[39\] vssd1 vssd1
+ vccd1 vccd1 _04987_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08894_ ks1.key_reg\[24\] _04735_ _04917_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_166_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09515_ _05312_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09446_ net211 vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_191_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09377_ _05345_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08328_ addroundkey_data_o\[8\] fifo_bank_register.data_out\[8\] _04468_ vssd1 vssd1
+ vccd1 vccd1 _04477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ net106 net95 net128 net117 vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__or4_1
XFILLER_0_201_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11270_ _06791_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10221_ _06001_ _06032_ _06033_ _06005_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10152_ sub1.ready_o vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_207_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput290 net290 vssd1 vssd1 vccd1 vccd1 data_o[127] sky130_fd_sc_hd__clkbuf_4
XTAP_5911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14960_ _03207_ _03234_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__xnor2_1
X_10083_ _05907_ _05908_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__xnor2_1
XTAP_5944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold9 ks1.key_reg\[44\] vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13911_ _02136_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__clkbuf_4
XTAP_5977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14891_ _03163_ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__nor2_8
XTAP_5999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16630_ net519 _00078_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_214_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13842_ fifo_bank_register.bank\[0\]\[31\] _02246_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16561_ net490 _00009_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_13773_ fifo_bank_register.bank\[1\]\[24\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10985_ _06722_ vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15512_ _03581_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__clkbuf_4
X_18300_ clknet_leaf_30_clk _01731_ net642 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[66\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12724_ fifo_bank_register.bank\[2\]\[27\] _05327_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07660_ sky130_fd_sc_hd__mux2_1
X_16492_ _04329_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_195_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18231_ clknet_leaf_36_clk _01662_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[61\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_183_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15443_ sub1.data_o\[27\] _05195_ _04879_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__mux2_1
X_12655_ _07622_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11606_ _07069_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18162_ clknet_leaf_81_clk _01593_ net578 vssd1 vssd1 vccd1 vccd1 ks1.col\[16\] sky130_fd_sc_hd__dfrtp_1
X_15374_ sub1.data_o\[35\] sub1.data_o\[99\] _03574_ vssd1 vssd1 vccd1 vccd1 _03583_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12586_ fifo_bank_register.bank\[3\]\[90\] _05459_ _07586_ vssd1 vssd1 vccd1 vccd1
+ _07587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17113_ net505 _00556_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14325_ fifo_bank_register.bank\[7\]\[85\] _02623_ _02632_ fifo_bank_register.bank\[2\]\[85\]
+ _02675_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a221o_1
X_18093_ net399 _01536_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[95\]
+ sky130_fd_sc_hd__dfxtp_1
X_11537_ _07032_ vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17044_ net516 _00487_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14256_ _02613_ fifo_bank_register.data_out\[77\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02615_ sky130_fd_sc_hd__mux2_1
X_11468_ _06996_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13207_ _07913_ vssd1 vssd1 vccd1 vccd1 _07914_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ _06211_ _06212_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14187_ _02142_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11399_ _06960_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ fifo_bank_register.bank\[1\]\[95\] _05470_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07878_ sky130_fd_sc_hd__mux2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ fifo_bank_register.bank\[1\]\[62\] _05401_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07842_ sky130_fd_sc_hd__mux2_1
X_17946_ net536 _01389_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_2_clk clknet_3_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17877_ net535 _01320_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16828_ clknet_leaf_73_clk _00272_ net590 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[119\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_215_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16759_ clknet_leaf_39_clk _00203_ net663 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[50\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_177_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09300_ net152 vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__buf_2
XFILLER_0_220_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_201_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09231_ _05104_ _04946_ _05236_ _05238_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a31o_1
X_18429_ clknet_leaf_16_clk _01859_ net630 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[114\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09162_ sbox1.ah_reg\[3\] sbox1.ah_reg\[2\] vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09093_ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_185_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_200_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09995_ net45 mix1.data_o\[24\] _05817_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__mux2_1
XTAP_5207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_229_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08946_ _04874_ _04872_ _04968_ _04969_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__o22a_2
XFILLER_0_215_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_192_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08877_ addroundkey_data_o\[96\] _04657_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__or2_1
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10770_ sub1.data_o\[100\] _06513_ _06527_ _06528_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06529_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09429_ fifo_bank_register.bank\[9\]\[52\] _05380_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12440_ _07510_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12371_ _07472_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14110_ fifo_bank_register.bank\[5\]\[61\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[61\]
+ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__a22o_1
X_11322_ _06919_ vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15090_ _03354_ _03361_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14041_ _02423_ fifo_bank_register.data_out\[53\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02424_ sky130_fd_sc_hd__mux2_1
X_11253_ _06882_ vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10204_ mix1.data_o\[44\] _05876_ _05993_ _05994_ sub1.data_o\[44\] vssd1 vssd1 vccd1
+ vccd1 _06019_ sky130_fd_sc_hd__a32o_1
XFILLER_0_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11184_ _05415_ fifo_bank_register.bank\[8\]\[69\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06846_ sky130_fd_sc_hd__mux2_1
X_17800_ net527 _01243_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
X_10135_ _05955_ _05956_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_207_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15992_ ks1.col\[6\] _03960_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__xor2_4
XTAP_5730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14943_ _03168_ _03217_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__xor2_2
X_10066_ mix1.data_o\[32\] _05576_ _05758_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__o21a_1
X_17731_ net494 _01174_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14874_ addroundkey_data_o\[8\] _04379_ _05607_ _03149_ vssd1 vssd1 vccd1 vccd1 _03150_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17662_ net571 _01105_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13825_ fifo_bank_register.bank\[7\]\[30\] _02218_ _02227_ fifo_bank_register.bank\[2\]\[30\]
+ _02230_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__a221o_1
X_16613_ net562 _00061_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_17593_ net432 _01036_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[115\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16544_ sub1.data_o\[112\] _05197_ _04356_ _03594_ vssd1 vssd1 vccd1 vccd1 _04357_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13756_ fifo_bank_register.bank\[6\]\[22\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10968_ addroundkey_data_o\[119\] _06707_ _05696_ vssd1 vssd1 vccd1 vccd1 _06708_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12707_ _07650_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16475_ _04320_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_1038 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13687_ fifo_bank_register.bank\[7\]\[16\] _08182_ _08191_ fifo_bank_register.bank\[2\]\[16\]
+ _02106_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10899_ _05623_ _06640_ _06644_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_155_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15426_ sub1.data_o\[20\] _03606_ _03617_ _03611_ vssd1 vssd1 vccd1 vccd1 _03618_
+ sky130_fd_sc_hd__a22o_1
X_18214_ clknet_leaf_84_clk _01645_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[44\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12638_ fifo_bank_register.bank\[3\]\[115\] _05512_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15357_ _03571_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__clkbuf_1
X_18145_ clknet_leaf_53_clk sbox1.ah\[3\] net656 vssd1 vssd1 vccd1 vccd1 sbox1.ah_reg\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12569_ fifo_bank_register.bank\[3\]\[82\] _05443_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14308_ fifo_bank_register.bank\[5\]\[83\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[83\]
+ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__a22o_1
X_18076_ net519 _01519_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[78\]
+ sky130_fd_sc_hd__dfxtp_1
X_15288_ net716 _03533_ _03144_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17027_ net525 _00470_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14239_ _02599_ fifo_bank_register.data_out\[75\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ addroundkey_data_o\[115\] mix1.data_o\[115\] _04656_ vssd1 vssd1 vccd1 vccd1
+ _04824_ sky130_fd_sc_hd__mux2_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09780_ _05637_ vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__clkbuf_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ ks1.state\[1\] _04737_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__nand2_2
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ net514 _01372_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_213_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08662_ addroundkey_data_o\[4\] mix1.data_o\[4\] _04666_ vssd1 vssd1 vccd1 vccd1
+ _04686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_205_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08593_ _04620_ vssd1 vssd1 vccd1 vccd1 next_state sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09214_ _05137_ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09145_ sbox1.ah_reg\[0\] _05155_ _05119_ sbox1.ah_reg\[3\] vssd1 vssd1 vccd1 vccd1
+ _05156_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09076_ _05087_ _05089_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09978_ _05813_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__xor2_1
XFILLER_0_60_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08929_ _04713_ _04951_ _04952_ _04716_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ fifo_bank_register.bank\[5\]\[41\] _05357_ _07244_ vssd1 vssd1 vccd1 vccd1
+ _07246_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ fifo_bank_register.bank\[5\]\[9\] _05288_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07209_ sky130_fd_sc_hd__mux2_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_197_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13610_ _08173_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10822_ _05619_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__clkbuf_4
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14590_ fifo_bank_register.bank\[7\]\[114\] _02866_ _02875_ fifo_bank_register.bank\[2\]\[114\]
+ _02911_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13541_ _08111_ vssd1 vssd1 vccd1 vccd1 _08112_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10753_ _05613_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16260_ _04202_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13472_ _08053_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10684_ net249 ks1.key_reg\[92\] _06324_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _03455_ _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12423_ fifo_bank_register.bank\[3\]\[13\] _05297_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16191_ _04126_ _04139_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15142_ _03160_ _03245_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_140_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12354_ _07463_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11305_ _05536_ fifo_bank_register.bank\[8\]\[127\] _06768_ vssd1 vssd1 vccd1 vccd1
+ _06909_ sky130_fd_sc_hd__mux2_1
X_15073_ _03329_ _03344_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_205_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12285_ _07427_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__clkbuf_1
X_14024_ fifo_bank_register.bank\[0\]\[51\] _02408_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02409_ sky130_fd_sc_hd__mux2_1
X_11236_ _06873_ vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_205_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11167_ _06837_ vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_207_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10118_ _04610_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11098_ _05329_ fifo_bank_register.bank\[8\]\[28\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06801_ sky130_fd_sc_hd__mux2_1
X_15975_ net187 ks1.key_reg\[36\] _03937_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__mux2_1
XTAP_5571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17714_ net450 _01157_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
X_10049_ _05829_ _05875_ _05877_ _05833_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14926_ sub1.data_o\[89\] _03063_ _03092_ sub1.data_o\[57\] vssd1 vssd1 vccd1 vccd1
+ _03201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_175_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17645_ net414 _01088_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14857_ sub1.data_o\[29\] _03100_ _03058_ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_202_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_216_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13808_ fifo_bank_register.bank\[0\]\[28\] _02215_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02216_ sky130_fd_sc_hd__mux2_1
X_14788_ _03063_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17576_ net445 _01019_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16527_ net744 _03514_ _04343_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__mux2_1
X_13739_ fifo_bank_register.bank\[1\]\[20\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16458_ _04310_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_170_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15409_ _03603_ _03593_ _05245_ _03605_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__a31o_1
XFILLER_0_171_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16389_ _04167_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18128_ clknet_leaf_21_clk _01571_ net639 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[82\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18059_ net528 _01502_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09901_ _05712_ _05743_ _05744_ _05716_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_223_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout505 net507 vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_2
XFILLER_0_226_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout516 net520 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09832_ net117 mix1.data_o\[8\] _05604_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__mux2_1
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__buf_2
Xfanout538 net542 vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__buf_2
XFILLER_0_158_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout549 net551 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__buf_2
X_09763_ mix1.data_o\[0\] _05586_ _05618_ _05621_ sub1.data_o\[0\] vssd1 vssd1 vccd1
+ vccd1 _05622_ sky130_fd_sc_hd__a32o_1
XFILLER_0_193_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08714_ ks1.state\[1\] _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09694_ _05562_ vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08645_ _04661_ _04664_ _04667_ _04668_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08576_ addroundkey_data_o\[126\] fifo_bank_register.data_out\[126\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__mux2_2
XFILLER_0_117_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_165_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09128_ sbox1.ah_reg\[3\] _05127_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__nand2_1
XFILLER_0_165_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09059_ _05074_ vssd1 vssd1 vccd1 vccd1 sbox1.next_alph\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_202_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12070_ fifo_bank_register.bank\[5\]\[103\] _05487_ _07310_ vssd1 vssd1 vccd1 vccd1
+ _07314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11021_ _05615_ _06752_ _06753_ _05567_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15760_ mix1.data_o\[81\] net755 _03808_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__mux2_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _07790_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14711_ _05104_ _04927_ _05560_ _03016_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__a31o_1
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11923_ fifo_bank_register.bank\[5\]\[33\] _05340_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07237_ sky130_fd_sc_hd__mux2_1
X_15691_ _03774_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__clkbuf_1
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ net565 _00873_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
X_14642_ fifo_bank_register.bank\[9\]\[120\] _08089_ _02955_ _02956_ _02957_ vssd1
+ vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__a2111o_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11854_ _07200_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__clkbuf_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10805_ net134 ks1.key_reg\[103\] _06402_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__mux2_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14573_ fifo_bank_register.bank\[5\]\[112\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[112\]
+ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a22o_1
X_17361_ net533 _00804_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11785_ _07163_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13524_ _08065_ _08094_ vssd1 vssd1 vccd1 vccd1 _08095_ sky130_fd_sc_hd__nor2_1
X_16312_ _04230_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17292_ net517 _00735_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[70\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10736_ net254 ks1.key_reg\[97\] _06402_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16243_ net216 ks1.key_reg\[62\] _03937_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13455_ _05516_ fifo_bank_register.bank\[0\]\[117\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ _06416_ _06434_ _06435_ _06420_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ fifo_bank_register.bank\[3\]\[5\] _05280_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07492_ sky130_fd_sc_hd__mux2_1
X_16174_ _04111_ _04113_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13386_ _05447_ fifo_bank_register.bank\[0\]\[84\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08009_ sky130_fd_sc_hd__mux2_1
X_10598_ _06090_ _06342_ sub1.data_o\[84\] _06079_ vssd1 vssd1 vccd1 vccd1 _06373_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_180_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15125_ _03167_ _03187_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_121_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12337_ _05483_ fifo_bank_register.bank\[4\]\[101\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15056_ _03199_ _03327_ _04624_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_220_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12268_ _07418_ vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_208_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14007_ fifo_bank_register.bank\[7\]\[50\] _02380_ _02389_ fifo_bank_register.bank\[2\]\[50\]
+ _02392_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a221o_1
X_11219_ _06864_ vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12199_ _07382_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__clkbuf_1
XTAP_6080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15958_ _05050_ _03930_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__or2_1
Xinput190 key_i[39] vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14909_ addroundkey_data_o\[87\] _03062_ _03091_ addroundkey_data_o\[55\] vssd1 vssd1
+ vccd1 vccd1 _03184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_204_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15889_ sub1.data_o\[97\] _03878_ _03876_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08430_ addroundkey_data_o\[56\] fifo_bank_register.data_out\[56\] _04523_ vssd1
+ vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__mux2_1
X_17628_ net501 _01071_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08361_ addroundkey_data_o\[23\] fifo_bank_register.data_out\[23\] _04490_ vssd1
+ vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17559_ net540 _01002_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08292_ _04445_ _04446_ _04447_ _04448_ vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09815_ mix1.data_o\[6\] _05586_ _05618_ _05621_ sub1.data_o\[6\] vssd1 vssd1 vccd1
+ vccd1 _05668_ sky130_fd_sc_hd__a32o_1
XFILLER_0_214_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09746_ net1 mix1.data_o\[0\] _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09677_ sub1.data_o\[120\] _05548_ _04891_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__mux2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_222_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08628_ state _04618_ _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _04598_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11570_ _07049_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10521_ sub1.data_o\[77\] _06302_ _06239_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13240_ _05301_ fifo_bank_register.bank\[0\]\[15\] _07926_ vssd1 vssd1 vccd1 vccd1
+ _07932_ sky130_fd_sc_hd__mux2_1
X_10452_ _05619_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13171_ _07895_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__clkbuf_1
X_10383_ sub1.data_o\[61\] _06180_ _06160_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12122_ _07340_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__buf_4
XFILLER_0_206_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12053_ fifo_bank_register.bank\[5\]\[95\] _05470_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07305_ sky130_fd_sc_hd__mux2_1
X_16930_ net410 _00373_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11004_ mix1.data_o\[124\] _05676_ _05758_ _05620_ sub1.data_o\[124\] vssd1 vssd1
+ vccd1 vccd1 _06739_ sky130_fd_sc_hd__a32o_1
XFILLER_0_217_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16861_ net483 _00304_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1082 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18600_ clknet_leaf_69_clk _02029_ net604 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[127\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_189_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15812_ mix1.data_o\[106\] net751 _03830_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16792_ clknet_leaf_26_clk _00236_ net649 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[83\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18531_ clknet_leaf_62_clk _01960_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[58\]
+ sky130_fd_sc_hd__dfrtp_1
X_15743_ mix1.data_o\[73\] net770 _03797_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__mux2_1
X_12955_ _07781_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__clkbuf_1
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11906_ fifo_bank_register.bank\[5\]\[25\] _05323_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07228_ sky130_fd_sc_hd__mux2_1
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ clknet_leaf_34_clk _01892_ net662 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[102\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_213_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15674_ mix1.data_o\[40\] net726 _03764_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ fifo_bank_register.bank\[2\]\[104\] _05489_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07745_ sky130_fd_sc_hd__mux2_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_262 net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17413_ net523 _00856_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_273 addroundkey_data_o\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ _07190_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__clkbuf_1
X_14625_ fifo_bank_register.bank\[1\]\[118\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[118\]
+ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__a22o_1
XFILLER_0_213_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_284 mix1.data_o\[36\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18393_ clknet_leaf_1_clk _01823_ net620 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[78\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_295 sub1.data_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ net492 _00787_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14556_ fifo_bank_register.bank\[6\]\[110\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[110\]
+ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11768_ _07154_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10719_ mix1.data_o\[96\] _06129_ _06398_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13507_ _05249_ _05266_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__xor2_1
XFILLER_0_153_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17275_ net562 _00718_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_14487_ fifo_bank_register.bank\[0\]\[102\] _02820_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11699_ _07118_ vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16226_ _04111_ _04113_ _04151_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__or3b_2
X_13438_ _05499_ fifo_bank_register.bank\[0\]\[109\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16157_ addroundkey_round\[1\] vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13369_ _05430_ fifo_bank_register.bank\[0\]\[76\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _08000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_224_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15108_ _03099_ _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16088_ net200 ks1.key_reg\[48\] _03910_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15039_ addroundkey_data_o\[27\] _04378_ _05607_ _03311_ vssd1 vssd1 vccd1 vccd1
+ _03312_ sky130_fd_sc_hd__a211o_1
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09600_ _05496_ vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09531_ fifo_bank_register.bank\[9\]\[85\] _05449_ _05439_ vssd1 vssd1 vccd1 vccd1
+ _05450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09462_ net217 vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_188_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08413_ addroundkey_data_o\[48\] fifo_bank_register.data_out\[48\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09393_ _05356_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08344_ addroundkey_data_o\[15\] fifo_bank_register.data_out\[15\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__mux2_2
XFILLER_0_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_172_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08275_ net252 net253 net254 net251 vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_203_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09729_ round\[1\] _04613_ round\[2\] vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__and3_1
XFILLER_0_214_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12740_ _07668_ vssd1 vssd1 vccd1 vccd1 _01083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ fifo_bank_register.bank\[2\]\[2\] _05274_ _07629_ vssd1 vssd1 vccd1 vccd1
+ _07632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ fifo_bank_register.bank\[1\]\[94\] _02721_ _02722_ fifo_bank_register.bank\[8\]\[94\]
+ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_167_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11622_ _07077_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__clkbuf_1
X_15390_ _04369_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__buf_4
XFILLER_0_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ fifo_bank_register.bank\[7\]\[87\] _02623_ _02632_ fifo_bank_register.bank\[2\]\[87\]
+ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__a221o_1
X_11553_ fifo_bank_register.bank\[7\]\[115\] _05512_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ sub1.data_o\[75\] _06287_ _06239_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__mux2_1
X_17060_ net447 _00503_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14272_ fifo_bank_register.bank\[0\]\[79\] _02628_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11484_ fifo_bank_register.bank\[7\]\[82\] _05443_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07005_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16011_ _05547_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__xor2_2
X_13223_ _05284_ fifo_bank_register.bank\[0\]\[7\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ net221 ks1.key_reg\[67\] _06166_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13154_ _07886_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10366_ _05707_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_209_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ fifo_bank_register.bank\[5\]\[120\] _05522_ _07198_ vssd1 vssd1 vccd1 vccd1
+ _07332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _07794_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__buf_4
X_17962_ net452 _01405_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
X_10297_ _06090_ _05972_ sub1.data_o\[53\] _06079_ vssd1 vssd1 vccd1 vccd1 _06103_
+ sky130_fd_sc_hd__a31o_1
X_16913_ net545 _00356_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
X_12036_ fifo_bank_register.bank\[5\]\[87\] _05453_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17893_ net438 _01336_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16844_ net425 _00287_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16775_ clknet_leaf_67_clk _00219_ net610 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[66\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13987_ fifo_bank_register.bank\[6\]\[48\] _02313_ _02314_ fifo_bank_register.bank\[4\]\[48\]
+ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a22o_1
XFILLER_0_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18514_ clknet_leaf_62_clk _01943_ net598 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
X_15726_ mix1.data_o\[65\] net733 _03786_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__mux2_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ fifo_bank_register.bank\[1\]\[0\] _05248_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07773_ sky130_fd_sc_hd__mux2_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18445_ clknet_leaf_9_clk _01875_ net632 vssd1 vssd1 vccd1 vccd1 sub1.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15657_ mix1.data_o\[32\] net694 _03753_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__mux2_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12869_ fifo_bank_register.bank\[2\]\[96\] _05472_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07736_ sky130_fd_sc_hd__mux2_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14608_ fifo_bank_register.bank\[1\]\[116\] _02883_ _02884_ fifo_bank_register.bank\[8\]\[116\]
+ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__a22o_1
X_18376_ clknet_leaf_35_clk _01806_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[61\]
+ sky130_fd_sc_hd__dfrtp_4
X_15588_ mix1.data_o\[0\] _03170_ mix1.next_ready_o vssd1 vssd1 vccd1 vccd1 _03720_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17327_ net467 _00770_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14539_ _08076_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17258_ net422 _00701_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16209_ _04155_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17189_ net402 _00632_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08962_ mix1.data_o\[47\] _04693_ _04695_ mix1.data_o\[39\] vssd1 vssd1 vccd1 vccd1
+ _04986_ sky130_fd_sc_hd__a22o_1
XFILLER_0_227_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08893_ ks1.key_reg\[24\] _04729_ _04731_ net174 vssd1 vssd1 vccd1 vccd1 _04917_
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09514_ net236 vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09445_ _05391_ vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__clkbuf_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ fifo_bank_register.bank\[9\]\[35\] _05344_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05345_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08327_ _04476_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__buf_2
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ net23 net12 net33 net32 vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__or4_1
XFILLER_0_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ mix1.data_o\[46\] _05876_ _05993_ _05994_ sub1.data_o\[46\] vssd1 vssd1 vccd1
+ vccd1 _06033_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _05613_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput280 net280 vssd1 vssd1 vccd1 vccd1 data_o[118] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput291 net291 vssd1 vssd1 vccd1 vccd1 data_o[12] sky130_fd_sc_hd__clkbuf_4
XTAP_5923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10082_ net184 ks1.key_reg\[33\] _05762_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__mux2_1
XTAP_5934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13910_ _02306_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__clkbuf_1
XTAP_5978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14890_ addroundkey_data_o\[127\] _03054_ _03165_ vssd1 vssd1 vccd1 vccd1 _03166_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13841_ fifo_bank_register.bank\[9\]\[31\] _02226_ _02243_ _02244_ _02245_ vssd1
+ vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_138_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13772_ fifo_bank_register.bank\[6\]\[24\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__a22o_1
X_16560_ net473 _00008_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10984_ addroundkey_data_o\[121\] _06721_ _05696_ vssd1 vssd1 vccd1 vccd1 _06722_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15511_ sub1.data_o\[19\] sub1.data_o\[83\] _03671_ vssd1 vssd1 vccd1 vccd1 _03672_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12723_ _07659_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_1236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16491_ net728 _03402_ _04321_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18230_ clknet_leaf_38_clk _01661_ net668 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[60\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15442_ _03627_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__clkbuf_1
X_12654_ fifo_bank_register.bank\[3\]\[123\] _05528_ _07485_ vssd1 vssd1 vccd1 vccd1
+ _07622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_167_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11605_ fifo_bank_register.bank\[6\]\[11\] _05293_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18161_ clknet_leaf_49_clk _01592_ net611 vssd1 vssd1 vccd1 vccd1 ks1.col\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_217_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15373_ _03582_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__clkbuf_1
X_12585_ _07508_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17112_ net533 _00555_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_14324_ fifo_bank_register.bank\[5\]\[85\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[85\]
+ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11536_ fifo_bank_register.bank\[7\]\[107\] _05495_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07032_ sky130_fd_sc_hd__mux2_1
X_18092_ net460 _01535_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14255_ _08068_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17043_ net546 _00486_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11467_ fifo_bank_register.bank\[7\]\[74\] _05426_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _06996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _06766_ _07483_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10418_ net219 ks1.key_reg\[65\] _06166_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14186_ _02140_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__clkbuf_4
X_11398_ fifo_bank_register.bank\[7\]\[41\] _05357_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _07877_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10349_ _06150_ vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13068_ _07841_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17945_ net563 _01388_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12019_ fifo_bank_register.bank\[5\]\[79\] _05436_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17876_ net535 _01319_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16827_ clknet_leaf_8_clk _00271_ net633 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[118\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_220_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16758_ clknet_leaf_39_clk _00202_ net668 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[49\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_220_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_159_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15709_ mix1.data_o\[57\] net715 _03775_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16689_ clknet_leaf_50_clk _00136_ net615 vssd1 vssd1 vccd1 vccd1 addroundkey_round\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_186_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09230_ sub1.data_o\[118\] _05197_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__a21o_1
XFILLER_0_158_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18428_ clknet_leaf_15_clk _01858_ net637 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[113\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_150_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09161_ _05154_ _05171_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18359_ clknet_leaf_84_clk _01789_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[44\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_185_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09092_ _04367_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09994_ _05615_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_229_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ _04833_ _04967_ _04649_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__a21o_1
XFILLER_0_228_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_192_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ _04698_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_196_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09428_ net205 vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09359_ net181 vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_165_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12370_ _05516_ fifo_bank_register.bank\[4\]\[117\] _07464_ vssd1 vssd1 vccd1 vccd1
+ _07472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11321_ fifo_bank_register.bank\[7\]\[5\] _05280_ _06913_ vssd1 vssd1 vccd1 vccd1
+ _06919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ fifo_bank_register.bank\[0\]\[53\] _02422_ _02401_ vssd1 vssd1 vccd1 vccd1
+ _02423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11252_ _05483_ fifo_bank_register.bank\[8\]\[101\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10203_ sub1.data_o\[44\] _06017_ _05991_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11183_ _06845_ vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10134_ net188 ks1.key_reg\[37\] _05920_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__mux2_4
XTAP_5720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ net133 ks1.key_reg\[102\] _03902_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__mux2_2
XTAP_5731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17730_ net494 _01173_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14942_ _03089_ _03216_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__xnor2_2
X_10065_ _05575_ _05890_ _05891_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__a21o_1
XTAP_5764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ net571 _01104_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14873_ addroundkey_data_o\[72\] _03144_ _03145_ addroundkey_data_o\[40\] vssd1 vssd1
+ vccd1 vccd1 _03149_ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_187_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_159_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16612_ net563 _00060_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_199_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13824_ fifo_bank_register.bank\[5\]\[30\] _02228_ _02229_ fifo_bank_register.bank\[3\]\[30\]
+ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__a22o_1
X_17592_ net408 _01035_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[114\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_202_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16543_ sub1.data_o\[80\] sub1.data_o\[16\] _03574_ vssd1 vssd1 vccd1 vccd1 _04356_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1022 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13755_ fifo_bank_register.bank\[7\]\[22\] _02128_ _02139_ fifo_bank_register.bank\[2\]\[22\]
+ _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a221o_1
X_10967_ _06705_ _06706_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_202_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ fifo_bank_register.bank\[2\]\[19\] _05309_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07650_ sky130_fd_sc_hd__mux2_1
X_16474_ _03171_ _03539_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__or2_1
X_10898_ sub1.data_o\[113\] _06513_ _06642_ _06643_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06644_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13686_ fifo_bank_register.bank\[5\]\[16\] _08192_ _08193_ fifo_bank_register.bank\[3\]\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18213_ clknet_leaf_84_clk _01644_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[43\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15425_ sub1.data_o\[116\] sub1.data_o\[52\] _03609_ vssd1 vssd1 vccd1 vccd1 _03617_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_171_915 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12637_ _07613_ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18144_ clknet_leaf_53_clk sbox1.ah\[2\] net656 vssd1 vssd1 vccd1 vccd1 sbox1.ah_reg\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_14_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15356_ net724 _03529_ _03145_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12568_ _07577_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_198_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14307_ _02660_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__clkbuf_1
X_11519_ fifo_bank_register.bank\[7\]\[99\] _05478_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07023_ sky130_fd_sc_hd__mux2_1
X_18075_ net555 _01518_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[77\]
+ sky130_fd_sc_hd__dfxtp_1
X_15287_ _03475_ _03532_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__xnor2_2
X_12499_ fifo_bank_register.bank\[3\]\[49\] _05373_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17026_ net515 _00469_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14238_ fifo_bank_register.bank\[0\]\[75\] _02598_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14169_ fifo_bank_register.bank\[6\]\[68\] _02475_ _02476_ fifo_bank_register.bank\[4\]\[68\]
+ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__a22o_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_226_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ ks1.key_reg\[17\] _04742_ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a21oi_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17928_ net527 _01371_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[66\]
+ sky130_fd_sc_hd__dfxtp_1
X_08661_ addroundkey_data_o\[60\] mix1.data_o\[60\] _04663_ vssd1 vssd1 vccd1 vccd1
+ _04685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17859_ net496 _01302_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08592_ next_first_round_reg _04619_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_220_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_5__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_220_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09213_ _05170_ _05191_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09144_ _05109_ _05110_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09075_ sbox1.ah\[2\] _05088_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__nand2_1
XFILLER_0_170_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09977_ net172 ks1.key_reg\[22\] _05708_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__mux2_4
XTAP_5027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ addroundkey_data_o\[93\] mix1.data_o\[93\] _04657_ vssd1 vssd1 vccd1 vccd1
+ _04952_ sky130_fd_sc_hd__mux2_1
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08859_ _04879_ _04881_ _04882_ _04668_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__a22o_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11870_ _07208_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__clkbuf_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _05757_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__clkbuf_4
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10752_ sub1.data_o\[99\] _06511_ _06478_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__mux2_1
X_13540_ _08110_ vssd1 vssd1 vccd1 vccd1 _08111_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_223_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13471_ _05532_ fifo_bank_register.bank\[0\]\[125\] _07914_ vssd1 vssd1 vccd1 vccd1
+ _08053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10683_ _06416_ _06448_ _06449_ _06420_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15210_ _03470_ _03471_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12422_ _07500_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16190_ _04113_ _04125_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__or2_1
XFILLER_0_168_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15141_ _03407_ _03408_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__xnor2_2
X_12353_ _05499_ fifo_bank_register.bank\[4\]\[109\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07463_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11304_ _06908_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15072_ _03336_ _03343_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_50_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12284_ _05430_ fifo_bank_register.bank\[4\]\[76\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14023_ fifo_bank_register.bank\[9\]\[51\] _02388_ _02405_ _02406_ _02407_ vssd1
+ vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a2111o_1
X_11235_ _05466_ fifo_bank_register.bank\[8\]\[93\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06873_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11166_ _05396_ fifo_bank_register.bank\[8\]\[60\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10117_ mix1.data_o\[36\] _05576_ _05916_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__o21a_1
XTAP_5550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11097_ _06800_ vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__clkbuf_1
X_15974_ _03943_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__xor2_2
XTAP_5561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17713_ net462 _01156_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14925_ _05201_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__nand2_2
X_10048_ mix1.data_o\[30\] _05876_ _05821_ _05822_ sub1.data_o\[30\] vssd1 vssd1 vccd1
+ vccd1 _05877_ sky130_fd_sc_hd__a32o_1
XFILLER_0_101_1099 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold90 mix1.data_reg\[75\] vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17644_ net416 _01087_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14856_ sub1.data_o\[93\] _03108_ _03066_ sub1.data_o\[61\] vssd1 vssd1 vccd1 vccd1
+ _03132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_187_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13807_ fifo_bank_register.bank\[9\]\[28\] _02137_ _02212_ _02213_ _02214_ vssd1
+ vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_212_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17575_ net448 _01018_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[97\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14787_ _03062_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__clkbuf_4
X_11999_ _07276_ vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16526_ _04347_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13738_ _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16457_ net815 _04309_ _03957_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__mux2_1
X_13669_ _02091_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_213_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15408_ sub1.data_o\[79\] _03600_ _03595_ sub1.data_o\[15\] vssd1 vssd1 vccd1 vccd1
+ _03605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16388_ _04271_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_186_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18127_ clknet_leaf_20_clk _01570_ net640 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[81\]
+ sky130_fd_sc_hd__dfrtp_4
X_15339_ _03562_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18058_ net513 _01501_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09900_ mix1.data_o\[15\] _05677_ _05703_ _05704_ sub1.data_o\[15\] vssd1 vssd1 vccd1
+ vccd1 _05744_ sky130_fd_sc_hd__a32o_1
X_17009_ net392 _00452_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout506 net507 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09831_ _05682_ vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__clkbuf_1
Xfanout517 net520 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_2
XFILLER_0_226_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout528 net529 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__clkbuf_2
Xfanout539 net542 vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__buf_1
XFILLER_0_225_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09762_ _05620_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08713_ ks1.state\[0\] ks1.state\[2\] vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__nor2_1
X_09693_ sub1.data_o\[123\] _05196_ _04891_ vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08644_ _04363_ _04364_ _04365_ _04362_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__and4bb_4
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08575_ _04606_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_117_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_194_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09127_ sbox1.ah_reg\[1\] _05119_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09058_ _05060_ _04923_ _05072_ _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11020_ mix1.data_o\[126\] _05676_ _05758_ _05620_ sub1.data_o\[126\] vssd1 vssd1
+ vccd1 vccd1 _06753_ sky130_fd_sc_hd__a32o_1
XFILLER_0_124_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ fifo_bank_register.bank\[1\]\[16\] _05303_ _07783_ vssd1 vssd1 vccd1 vccd1
+ _07790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_172_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ sub1.data_o\[82\] _03010_ _03015_ sub1.next_ready_o vssd1 vssd1 vccd1 vccd1
+ _03016_ sky130_fd_sc_hd__a22o_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _07236_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__clkbuf_1
X_15690_ mix1.data_o\[48\] net741 _03764_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__mux2_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ fifo_bank_register.bank\[1\]\[120\] _08111_ _08114_ fifo_bank_register.bank\[8\]\[120\]
+ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__a22o_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ fifo_bank_register.bank\[5\]\[0\] _05248_ _07199_ vssd1 vssd1 vccd1 vccd1
+ _07200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _05623_ _06555_ _06559_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__o21ai_4
X_17360_ net496 _00803_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_11784_ fifo_bank_register.bank\[6\]\[96\] _05472_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07163_ sky130_fd_sc_hd__mux2_1
X_14572_ _02896_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__clkbuf_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16311_ net807 _04121_ _04222_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13523_ fifo_bank_register.read_ptr\[3\] fifo_bank_register.read_ptr\[2\] vssd1 vssd1
+ vccd1 vccd1 _08094_ sky130_fd_sc_hd__or2b_1
XFILLER_0_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10735_ _06381_ _06490_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_153_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17291_ net512 _00734_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[69\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16242_ _04185_ _04186_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__xor2_4
X_10666_ mix1.data_o\[90\] _06296_ _06320_ _06321_ sub1.data_o\[90\] vssd1 vssd1 vccd1
+ vccd1 _06435_ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13454_ _08044_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12405_ _07491_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_207_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16173_ _04123_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__clkbuf_1
X_13385_ _08008_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__clkbuf_1
X_10597_ sub1.data_o\[84\] _06371_ _06113_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ _03393_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12336_ _07454_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15055_ _03282_ _03326_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12267_ _05413_ fifo_bank_register.bank\[4\]\[68\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11218_ _05449_ fifo_bank_register.bank\[8\]\[85\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06864_ sky130_fd_sc_hd__mux2_1
X_14006_ fifo_bank_register.bank\[5\]\[50\] _02390_ _02391_ fifo_bank_register.bank\[3\]\[50\]
+ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__a22o_1
XFILLER_0_208_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12198_ _05344_ fifo_bank_register.bank\[4\]\[35\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11149_ _05380_ fifo_bank_register.bank\[8\]\[52\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06828_ sky130_fd_sc_hd__mux2_1
XTAP_6070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15957_ _03928_ _03929_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__xor2_1
XTAP_5391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput180 key_i[2] vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_4
XFILLER_0_218_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput191 key_i[3] vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__buf_4
X_14908_ sub1.data_o\[119\] _03077_ _03182_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_163_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _05553_ sub1.data_o\[65\] _05200_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17627_ net483 _01070_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14839_ _03111_ _03114_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__nor2_4
XFILLER_0_148_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08360_ _04494_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_148_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17558_ net540 _01001_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16509_ _04338_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08291_ net221 net220 net222 net223 vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__or4b_1
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17489_ net503 _00932_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_184_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_183_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_171_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09814_ sub1.data_o\[6\] _05666_ _05610_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__buf_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08627_ net129 mix1.ready_o _04650_ addroundkey_ready_o vssd1 vssd1 vccd1 vccd1 _04651_
+ sky130_fd_sc_hd__a22oi_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08558_ addroundkey_data_o\[117\] fifo_bank_register.data_out\[117\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__mux2_4
XFILLER_0_132_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_181_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08489_ addroundkey_data_o\[84\] fifo_bank_register.data_out\[84\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__mux2_4
XFILLER_0_135_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ net103 mix1.data_o\[77\] _06237_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10451_ _05757_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_165_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13170_ fifo_bank_register.bank\[1\]\[110\] _05501_ _07894_ vssd1 vssd1 vccd1 vccd1
+ _07895_ sky130_fd_sc_hd__mux2_1
X_10382_ net86 mix1.data_o\[61\] _06158_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_206_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12121_ _06766_ _06910_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_206_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12052_ _07304_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11003_ sub1.data_o\[124\] _06737_ _05609_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__mux2_1
X_16860_ net501 _00303_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_15811_ _03837_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16791_ clknet_leaf_24_clk _00235_ net649 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[82\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18530_ clknet_leaf_60_clk _01959_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[57\]
+ sky130_fd_sc_hd__dfrtp_1
X_15742_ _03801_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12954_ fifo_bank_register.bank\[1\]\[8\] _05286_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18461_ clknet_leaf_32_clk _01891_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[101\]
+ sky130_fd_sc_hd__dfrtp_4
X_11905_ _07227_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_217_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15673_ _03765_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__clkbuf_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12885_ _07744_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_241 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_200_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17412_ net523 _00855_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_252 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_263 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14624_ fifo_bank_register.bank\[6\]\[118\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[118\]
+ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a22o_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18392_ clknet_leaf_1_clk _01822_ net620 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[77\]
+ sky130_fd_sc_hd__dfrtp_4
X_11836_ fifo_bank_register.bank\[6\]\[121\] _05524_ _07055_ vssd1 vssd1 vccd1 vccd1
+ _07190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_274 addroundkey_data_o\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 mix1.data_o\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_296 sub1.data_o\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17343_ net490 _00786_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ _02148_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_184_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11767_ fifo_bank_register.bank\[6\]\[88\] _05455_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _08072_ _08081_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10718_ _06126_ _06479_ _06480_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17274_ net562 _00717_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ fifo_bank_register.bank\[9\]\[102\] _02793_ _02817_ _02818_ _02819_ vssd1
+ vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a2111o_1
X_11698_ fifo_bank_register.bank\[6\]\[55\] _05386_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16225_ _04171_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13437_ _08035_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10649_ _04609_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16156_ _04107_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13368_ _07999_ vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15107_ _03198_ _03376_ _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_80_1227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12319_ _07445_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_220_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16087_ _04044_ _04045_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__xor2_2
XFILLER_0_224_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13299_ _07963_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__clkbuf_1
X_15038_ addroundkey_data_o\[91\] _03064_ _03084_ addroundkey_data_o\[59\] vssd1 vssd1
+ vccd1 vccd1 _03311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16989_ net487 _00432_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09530_ net241 vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09461_ _05402_ vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_815 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_176_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ _04521_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09392_ fifo_bank_register.bank\[9\]\[40\] _05354_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08343_ _04485_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ net243 net245 net244 net242 vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_162_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_203_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09728_ round\[2\] _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__and2_1
X_09659_ net160 vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_195_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_215_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _07631_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11621_ fifo_bank_register.bank\[6\]\[19\] _05309_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_166_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14340_ fifo_bank_register.bank\[5\]\[87\] _02633_ _02634_ fifo_bank_register.bank\[3\]\[87\]
+ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11552_ _07040_ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ net101 mix1.data_o\[75\] _06237_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11483_ _07004_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__clkbuf_1
X_14271_ fifo_bank_register.bank\[9\]\[79\] _02550_ _02625_ _02626_ _02627_ vssd1
+ vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_107_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_190_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16010_ net135 ks1.key_reg\[104\] _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__mux2_1
X_10434_ _06171_ _06224_ _06225_ _06175_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__a22o_1
X_13222_ _07922_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ _06001_ _06161_ _06164_ _06005_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__a22o_1
X_13153_ fifo_bank_register.bank\[1\]\[102\] _05485_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _07331_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__clkbuf_1
X_13084_ _07849_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__clkbuf_1
X_17961_ net447 _01404_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10296_ sub1.data_o\[53\] _06101_ _05936_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__mux2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16912_ net545 _00355_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
X_12035_ _07295_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17892_ net438 _01335_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16843_ net421 _00286_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16774_ clknet_leaf_47_clk _00218_ net651 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[65\]
+ sky130_fd_sc_hd__dfrtp_4
X_13986_ fifo_bank_register.bank\[7\]\[48\] _02299_ _02308_ fifo_bank_register.bank\[2\]\[48\]
+ _02373_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18513_ clknet_leaf_59_clk _01942_ net605 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_15725_ _03792_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12937_ _07771_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18444_ clknet_leaf_8_clk _01874_ net632 vssd1 vssd1 vccd1 vccd1 sub1.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15656_ _03756_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__clkbuf_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _07735_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ fifo_bank_register.bank\[6\]\[116\] _02880_ _02881_ fifo_bank_register.bank\[4\]\[116\]
+ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a22o_1
X_18375_ clknet_leaf_38_clk _01805_ net669 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[60\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11819_ _07181_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__clkbuf_1
X_15587_ _03717_ _03709_ _05245_ _03719_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a31o_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12799_ _07699_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__clkbuf_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17326_ net462 _00769_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14538_ _02865_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17257_ net416 _00700_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_14469_ fifo_bank_register.bank\[9\]\[100\] _02793_ _02798_ _02801_ _02804_ vssd1
+ vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16208_ net248 ks1.key_reg\[91\] _03979_ vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__mux2_2
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17188_ net455 _00631_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ ks1.col\[22\] _04091_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__xor2_2
XFILLER_0_45_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_224_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08961_ _04975_ _04978_ _04981_ _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__or4_1
XFILLER_0_227_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08892_ _04741_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__inv_4
XFILLER_0_224_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09513_ _05437_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_189_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09444_ fifo_bank_register.bank\[9\]\[57\] _05390_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ net186 vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__buf_2
XFILLER_0_148_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08326_ addroundkey_data_o\[7\] fifo_bank_register.data_out\[7\] _04468_ vssd1 vssd1
+ vccd1 vccd1 _04476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08257_ _04398_ _04403_ _04408_ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10150_ sub1.data_o\[39\] _05969_ _05936_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput270 net270 vssd1 vssd1 vccd1 vccd1 data_o[109] sky130_fd_sc_hd__buf_2
XFILLER_0_203_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput281 net281 vssd1 vssd1 vccd1 vccd1 data_o[119] sky130_fd_sc_hd__clkbuf_4
Xoutput292 net292 vssd1 vssd1 vccd1 vccd1 data_o[13] sky130_fd_sc_hd__clkbuf_4
XTAP_5902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ _05899_ _05901_ _05906_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__o21ai_4
XTAP_5924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_226_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13840_ fifo_bank_register.bank\[1\]\[31\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[31\]
+ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_215_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ fifo_bank_register.bank\[7\]\[24\] _02128_ _02139_ fifo_bank_register.bank\[2\]\[24\]
+ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__a221o_1
XFILLER_0_173_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10983_ _06719_ _06720_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15510_ _05202_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ fifo_bank_register.bank\[2\]\[26\] _05325_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07659_ sky130_fd_sc_hd__mux2_1
X_16490_ _04328_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15441_ sub1.data_o\[26\] _05559_ _04879_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _07621_ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18160_ clknet_leaf_48_clk _01591_ net612 vssd1 vssd1 vccd1 vccd1 ks1.col\[30\] sky130_fd_sc_hd__dfrtp_2
X_11604_ _07068_ vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__clkbuf_1
X_15372_ sub1.data_o\[2\] _03580_ _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12584_ _07585_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__clkbuf_1
X_17111_ net532 _00554_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14323_ _02674_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18091_ net434 _01534_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_11535_ _07031_ vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17042_ net545 _00485_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14254_ fifo_bank_register.bank\[0\]\[77\] _02612_ _02563_ vssd1 vssd1 vccd1 vccd1
+ _02613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11466_ _06995_ vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13205_ _07912_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__clkbuf_1
X_10417_ _06171_ _06209_ _06210_ _06175_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11397_ _06959_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14185_ _02138_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13136_ fifo_bank_register.bank\[1\]\[94\] _05468_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07877_ sky130_fd_sc_hd__mux2_1
X_10348_ addroundkey_data_o\[57\] _06149_ _06064_ vssd1 vssd1 vccd1 vccd1 _06150_
+ sky130_fd_sc_hd__mux2_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_209_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ addroundkey_data_o\[51\] _06086_ _06064_ vssd1 vssd1 vccd1 vccd1 _06087_
+ sky130_fd_sc_hd__mux2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ fifo_bank_register.bank\[1\]\[61\] _05399_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17944_ net562 _01387_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[82\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12018_ _07286_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_218_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17875_ net506 _01318_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[13\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16826_ clknet_leaf_76_clk _00270_ net586 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[117\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_191_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16757_ clknet_leaf_66_clk _00201_ net603 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[48\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_177_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13969_ fifo_bank_register.bank\[7\]\[46\] _02299_ _02308_ fifo_bank_register.bank\[2\]\[46\]
+ _02358_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__a221o_1
XFILLER_0_220_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15708_ _03783_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16688_ clknet_leaf_49_clk ks1.next_ready_o net615 vssd1 vssd1 vccd1 vccd1 ks1.ready_o
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15639_ _03747_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18427_ clknet_leaf_15_clk _01857_ net636 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[112\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_111_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09160_ _05163_ _05170_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__xor2_4
XFILLER_0_111_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18358_ clknet_leaf_83_clk _01788_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[43\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17309_ net538 _00752_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[87\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09091_ _05100_ _05102_ vssd1 vssd1 vccd1 vccd1 sbox1.intermediate_to_invert_var\[0\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18289_ clknet_leaf_26_clk _01720_ net649 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[55\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_185_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ _05828_ vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_228_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08944_ _04833_ _04967_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__nor2_1
XFILLER_0_209_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ _04897_ _04898_ _04698_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ _05379_ vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_165_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09358_ _05332_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08309_ _04393_ _04436_ _04444_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__nor4_4
XFILLER_0_180_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09289_ _05285_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ _06918_ vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ _06881_ vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10202_ net67 mix1.data_o\[44\] _05989_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11182_ _05413_ fifo_bank_register.bank\[8\]\[68\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_197_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10133_ _05899_ _05948_ _05954_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_140_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15990_ _03959_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__clkbuf_1
XTAP_5721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10064_ _05201_ _05754_ sub1.data_o\[32\] _05585_ vssd1 vssd1 vccd1 vccd1 _05891_
+ sky130_fd_sc_hd__a31o_1
X_14941_ _03212_ _03215_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__nor2_4
XTAP_5754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17660_ net556 _01103_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ sub1.data_o\[104\] _03143_ _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_215_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16611_ net573 _00059_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
X_13823_ _02142_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17591_ net429 _01034_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_214_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16542_ _04355_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ fifo_bank_register.bank\[5\]\[22\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[22\]
+ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10966_ net151 ks1.key_reg\[119\] _04639_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12705_ _07649_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16473_ net705 _03060_ _03053_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13685_ _02105_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__clkbuf_1
X_10897_ mix1.data_o\[113\] _06494_ _05617_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__o21a_1
X_18212_ clknet_leaf_84_clk _01643_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[42\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15424_ _03603_ _04949_ _05196_ _03616_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12636_ fifo_bank_register.bank\[3\]\[114\] _05510_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_171_927 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18143_ clknet_leaf_53_clk sbox1.ah\[1\] net657 vssd1 vssd1 vccd1 vccd1 sbox1.ah_reg\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15355_ _03570_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_182_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12567_ fifo_bank_register.bank\[3\]\[81\] _05441_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14306_ _02659_ fifo_bank_register.data_out\[82\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18074_ net516 _01517_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[76\]
+ sky130_fd_sc_hd__dfxtp_2
X_11518_ _07022_ vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__clkbuf_1
X_15286_ _03380_ _03531_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12498_ _07540_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17025_ net572 _00468_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
X_14237_ fifo_bank_register.bank\[9\]\[75\] _02550_ _02595_ _02596_ _02597_ vssd1
+ vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_123_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11449_ _06986_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14168_ fifo_bank_register.bank\[7\]\[68\] _02461_ _02470_ fifo_bank_register.bank\[2\]\[68\]
+ _02535_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a221o_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13119_ fifo_bank_register.bank\[1\]\[86\] _05451_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _02146_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__clkbuf_4
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ net526 _01370_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[65\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08660_ _04362_ _04363_ _04365_ _04364_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__nor4b_4
X_17858_ net531 _01301_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16809_ clknet_leaf_81_clk _00253_ net586 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[100\]
+ sky130_fd_sc_hd__dfrtp_4
X_08591_ addroundkey_ready_o _04618_ _04611_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_220_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17789_ net571 _01232_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09212_ _05104_ _04946_ _05219_ _05221_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_228_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_1228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09143_ _05137_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09074_ _05067_ _05077_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_163_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09976_ _05712_ _05811_ _05812_ _05716_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a22o_1
XFILLER_0_228_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08927_ addroundkey_data_o\[69\] mix1.data_o\[69\] _04702_ vssd1 vssd1 vccd1 vccd1
+ _04951_ sky130_fd_sc_hd__mux2_1
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08858_ addroundkey_data_o\[72\] mix1.data_o\[72\] _04702_ vssd1 vssd1 vccd1 vccd1
+ _04882_ sky130_fd_sc_hd__mux2_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _04710_ _04811_ _04812_ _04684_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__a22o_1
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ sub1.data_o\[105\] _06572_ _06573_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__mux2_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10751_ net127 mix1.data_o\[99\] _06476_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_223_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13470_ _08052_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_211_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ mix1.data_o\[92\] _06296_ _06320_ _06321_ sub1.data_o\[92\] vssd1 vssd1 vccd1
+ vccd1 _06449_ sky130_fd_sc_hd__a32o_1
XFILLER_0_192_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12421_ fifo_bank_register.bank\[3\]\[12\] _05295_ _07497_ vssd1 vssd1 vccd1 vccd1
+ _07500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15140_ _03090_ _03216_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_168_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12352_ _07462_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11303_ _05534_ fifo_bank_register.bank\[8\]\[126\] _06768_ vssd1 vssd1 vccd1 vccd1
+ _06908_ sky130_fd_sc_hd__mux2_1
X_15071_ _03339_ _03342_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__nor2_8
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12283_ _07426_ vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__clkbuf_1
X_14022_ fifo_bank_register.bank\[1\]\[51\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[51\]
+ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a22o_1
X_11234_ _06872_ vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11165_ _06791_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__buf_4
XFILLER_0_207_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10116_ _05575_ _05937_ _05938_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__a21o_1
X_11096_ _05327_ fifo_bank_register.bank\[8\]\[27\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06800_ sky130_fd_sc_hd__mux2_1
X_15973_ net222 ks1.key_reg\[68\] _03906_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__mux2_1
XFILLER_0_207_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14924_ _03141_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__xnor2_2
X_10047_ _05585_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17712_ net464 _01155_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[106\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_222_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold80 mix1.data_reg\[69\] vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 mix1.data_reg\[88\] vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14855_ _03127_ _03130_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__nor2_8
X_17643_ net414 _01086_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_202_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13806_ fifo_bank_register.bank\[1\]\[28\] _02152_ _02154_ fifo_bank_register.bank\[8\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__a22o_1
X_17574_ net445 _01017_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[96\]
+ sky130_fd_sc_hd__dfxtp_1
X_14786_ _03061_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__buf_4
XFILLER_0_212_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11998_ fifo_bank_register.bank\[5\]\[69\] _05415_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16525_ net790 _03510_ _04343_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__mux2_1
X_13737_ _08113_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__buf_6
X_10949_ sub1.data_o\[118\] _06689_ _05608_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16456_ _04144_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13668_ _02090_ fifo_bank_register.data_out\[13\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _02091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15407_ _03603_ _03593_ _05236_ _03604_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__a31o_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ fifo_bank_register.bank\[3\]\[106\] _05493_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16387_ net844 _04157_ _04264_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__mux2_1
X_13599_ fifo_bank_register.bank\[0\]\[6\] _08163_ _08121_ vssd1 vssd1 vccd1 vccd1
+ _08164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18126_ clknet_leaf_20_clk _01569_ net640 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[80\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_182_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15338_ net764 _03502_ _03560_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ net574 _01500_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[59\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15269_ _03232_ _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17008_ net394 _00451_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[42\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_223_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09830_ addroundkey_data_o\[7\] _05681_ next_addroundkey_ready_o vssd1 vssd1 vccd1
+ vccd1 _05682_ sky130_fd_sc_hd__mux2_1
Xfanout507 net530 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__buf_2
Xfanout518 net520 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__buf_2
XFILLER_0_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_226_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09761_ _05619_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_226_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08712_ net161 ks1.key_reg\[12\] _04735_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09692_ _05561_ vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08643_ addroundkey_data_o\[76\] mix1.data_o\[76\] _04666_ vssd1 vssd1 vccd1 vccd1
+ _04667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08574_ addroundkey_data_o\[125\] fifo_bank_register.data_out\[125\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__mux2_2
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_194_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_61_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09126_ _05123_ _05136_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09057_ _04966_ _05055_ _04649_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ mix1.data_o\[20\] _05797_ _05703_ _05704_ sub1.data_o\[20\] vssd1 vssd1 vccd1
+ vccd1 _05798_ sky130_fd_sc_hd__a32o_1
XFILLER_0_102_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _07789_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ fifo_bank_register.bank\[5\]\[32\] _05338_ _07233_ vssd1 vssd1 vccd1 vccd1
+ _07236_ sky130_fd_sc_hd__mux2_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ fifo_bank_register.bank\[6\]\[120\] _08104_ _08107_ fifo_bank_register.bank\[4\]\[120\]
+ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__a22o_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _07198_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__buf_4
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ sub1.data_o\[103\] _06513_ _06557_ _06558_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06559_ sky130_fd_sc_hd__a221o_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _02895_ fifo_bank_register.data_out\[111\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02896_ sky130_fd_sc_hd__mux2_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _07162_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_clk clknet_3_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16310_ _04229_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__clkbuf_1
X_13522_ _08092_ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__clkbuf_4
X_10734_ sub1.data_o\[97\] _06341_ _06493_ _06495_ _06483_ vssd1 vssd1 vccd1 vccd1
+ _06496_ sky130_fd_sc_hd__a221o_1
X_17290_ net522 _00733_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ net251 ks1.key_reg\[94\] _03918_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__mux2_2
X_13453_ _05514_ fifo_bank_register.bank\[0\]\[116\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665_ sub1.data_o\[90\] _06433_ _06318_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_192_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12404_ fifo_bank_register.bank\[3\]\[4\] _05278_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16172_ ks1.key_reg\[24\] _04122_ _04106_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13384_ _05445_ fifo_bank_register.bank\[0\]\[83\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08008_ sky130_fd_sc_hd__mux2_1
X_10596_ net111 mix1.data_o\[84\] _06111_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15123_ net697 _03392_ _03171_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__mux2_1
X_12335_ _05480_ fifo_bank_register.bank\[4\]\[100\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15054_ _03233_ _03304_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_107_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12266_ _07417_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14005_ _02142_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11217_ _06863_ vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12197_ _07381_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11148_ _06827_ vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__clkbuf_1
XTAP_6071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11079_ _06790_ vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__clkbuf_1
X_15956_ net185 ks1.key_reg\[34\] _03910_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__mux2_1
Xinput170 key_i[20] vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_4
XTAP_5381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput181 key_i[30] vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_4
XTAP_5392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14907_ sub1.data_o\[23\] _04375_ _03058_ _03181_ vssd1 vssd1 vccd1 vccd1 _03182_
+ sky130_fd_sc_hd__a211o_1
Xinput192 key_i[40] vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__buf_4
X_15887_ _03877_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_203_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17626_ net512 _01069_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14838_ addroundkey_data_o\[117\] _03055_ _03113_ vssd1 vssd1 vccd1 vccd1 _03114_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17557_ net547 _01000_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
X_14769_ _03048_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_clk clknet_3_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16508_ net745 _03484_ _04332_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17488_ net493 _00931_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_08290_ net217 net216 net219 net218 vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16439_ net794 _04060_ _04295_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18109_ net454 _01552_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[111\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09813_ net95 mix1.data_o\[6\] _05604_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09744_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__buf_4
XFILLER_0_213_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09675_ _04649_ _05153_ _05545_ _05546_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_119_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _04617_ _04616_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__or2_4
XFILLER_0_210_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _04597_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__buf_1
XFILLER_0_221_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_34_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ _04561_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_175_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10450_ sub1.data_o\[69\] _06238_ _06239_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09109_ _05109_ _05110_ _05119_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10381_ _06179_ vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_1264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12120_ _07339_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12051_ fifo_bank_register.bank\[5\]\[94\] _05468_ _07299_ vssd1 vssd1 vccd1 vccd1
+ _07304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11002_ net28 mix1.data_o\[124\] _05603_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__mux2_1
X_15810_ mix1.data_o\[105\] net687 _03830_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__mux2_1
X_16790_ clknet_leaf_26_clk _00234_ net649 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[81\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_176_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_176_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15741_ mix1.data_o\[72\] net769 _03797_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__mux2_1
X_12953_ _07780_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__clkbuf_1
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ fifo_bank_register.bank\[5\]\[24\] _05321_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07227_ sky130_fd_sc_hd__mux2_1
X_15672_ mix1.data_o\[39\] net791 _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__mux2_1
X_18460_ clknet_leaf_32_clk _01890_ net661 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[100\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_213_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_220 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12884_ fifo_bank_register.bank\[2\]\[103\] _05487_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07744_ sky130_fd_sc_hd__mux2_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_185_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_197_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_185_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17411_ net524 _00854_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_14623_ fifo_bank_register.bank\[7\]\[118\] _02866_ _02875_ fifo_bank_register.bank\[2\]\[118\]
+ _02940_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__a221o_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_253 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_158_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18391_ clknet_leaf_0_clk _01821_ net620 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[76\]
+ sky130_fd_sc_hd__dfrtp_2
X_11835_ _07189_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__clkbuf_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_213_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_264 _04468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_275 addroundkey_data_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_286 mix1.data_o\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17342_ net441 _00785_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_297 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _02146_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _07153_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13505_ _08071_ _08074_ _08056_ vssd1 vssd1 vccd1 vccd1 _08081_ sky130_fd_sc_hd__a21oi_1
X_10717_ _06395_ _06342_ sub1.data_o\[96\] _06384_ vssd1 vssd1 vccd1 vccd1 _06480_
+ sky130_fd_sc_hd__a31o_1
X_17273_ net572 _00716_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14485_ fifo_bank_register.bank\[1\]\[102\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[102\]
+ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11697_ _07117_ vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16224_ ks1.key_reg\[28\] _04170_ _04106_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__mux2_1
X_13436_ _05497_ fifo_bank_register.bank\[0\]\[108\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08035_ sky130_fd_sc_hd__mux2_1
X_10648_ mix1.data_o\[88\] _06296_ _06320_ _06321_ sub1.data_o\[88\] vssd1 vssd1 vccd1
+ vccd1 _06419_ sky130_fd_sc_hd__a32o_1
XFILLER_0_183_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16155_ ks1.key_reg\[23\] _04105_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13367_ _05428_ fifo_bank_register.bank\[0\]\[75\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _07999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10579_ sub1.data_o\[82\] _06341_ _06354_ _06355_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06356_ sky130_fd_sc_hd__a221o_1
XFILLER_0_183_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15106_ _03198_ _03376_ _06630_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12318_ _05464_ fifo_bank_register.bank\[4\]\[92\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_1239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16086_ net236 ks1.key_reg\[80\] _03907_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13298_ _05359_ fifo_bank_register.bank\[0\]\[42\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15037_ sub1.data_o\[123\] _03057_ _03309_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12249_ _07408_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_223_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16988_ net501 _00431_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_218_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15939_ _04371_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__buf_4
XFILLER_0_211_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09460_ fifo_bank_register.bank\[9\]\[62\] _05401_ _05397_ vssd1 vssd1 vccd1 vccd1
+ _05402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08411_ addroundkey_data_o\[47\] fifo_bank_register.data_out\[47\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__mux2_4
XFILLER_0_114_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17609_ net475 _01052_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09391_ _05312_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__buf_4
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18589_ clknet_leaf_81_clk _02018_ net586 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[116\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08342_ addroundkey_data_o\[14\] fifo_bank_register.data_out\[14\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__mux2_2
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_157_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08273_ net248 net247 net249 net250 vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__or4b_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_196_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_195_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_227_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09727_ round\[1\] _04613_ _05574_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__or3_1
XFILLER_0_214_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09658_ _05535_ vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__clkbuf_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_195_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08609_ round\[3\] addroundkey_round\[3\] vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__xor2_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ net135 vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__buf_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _07076_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11551_ fifo_bank_register.bank\[7\]\[114\] _05510_ _07035_ vssd1 vssd1 vccd1 vccd1
+ _07040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10502_ _06286_ vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__clkbuf_1
X_14270_ fifo_bank_register.bank\[1\]\[79\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[79\]
+ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a22o_1
X_11482_ fifo_bank_register.bank\[7\]\[81\] _05441_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13221_ _05282_ fifo_bank_register.bank\[0\]\[6\] _07915_ vssd1 vssd1 vccd1 vccd1
+ _07922_ sky130_fd_sc_hd__mux2_1
X_10433_ mix1.data_o\[67\] _06217_ _06162_ _06163_ sub1.data_o\[67\] vssd1 vssd1 vccd1
+ vccd1 _06225_ sky130_fd_sc_hd__a32o_1
XFILLER_0_208_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13152_ _07885_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__clkbuf_1
X_10364_ mix1.data_o\[59\] _06138_ _06162_ _06163_ sub1.data_o\[59\] vssd1 vssd1 vccd1
+ vccd1 _06164_ sky130_fd_sc_hd__a32o_1
XFILLER_0_108_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ fifo_bank_register.bank\[5\]\[119\] _05520_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ fifo_bank_register.bank\[1\]\[69\] _05415_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07849_ sky130_fd_sc_hd__mux2_1
X_17960_ net447 _01403_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[98\]
+ sky130_fd_sc_hd__dfxtp_1
X_10295_ net77 mix1.data_o\[53\] _05934_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16911_ net552 _00354_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
X_12034_ fifo_bank_register.bank\[5\]\[86\] _05451_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07295_ sky130_fd_sc_hd__mux2_1
X_17891_ net492 _01334_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16842_ net420 _00285_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_205_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13985_ fifo_bank_register.bank\[5\]\[48\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[48\]
+ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__a22o_1
X_16773_ clknet_leaf_67_clk _00217_ net610 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[64\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18512_ clknet_leaf_66_clk _01941_ net604 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[39\]
+ sky130_fd_sc_hd__dfrtp_1
X_15724_ mix1.data_o\[64\] mix1.data_reg\[64\] _03786_ vssd1 vssd1 vccd1 vccd1 _03792_
+ sky130_fd_sc_hd__mux2_1
X_12936_ _07770_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__buf_4
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_198_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18443_ clknet_leaf_9_clk _01873_ net632 vssd1 vssd1 vccd1 vccd1 sub1.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15655_ mix1.data_o\[31\] _03537_ _03753_ vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__mux2_1
X_12867_ fifo_bank_register.bank\[2\]\[95\] _05470_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07735_ sky130_fd_sc_hd__mux2_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14606_ fifo_bank_register.bank\[7\]\[116\] _02866_ _02875_ fifo_bank_register.bank\[2\]\[116\]
+ _02925_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__a221o_1
X_11818_ fifo_bank_register.bank\[6\]\[112\] _05506_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_201_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18374_ clknet_leaf_38_clk _01804_ net668 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[59\]
+ sky130_fd_sc_hd__dfrtp_4
X_15586_ sub1.data_o\[15\] _03660_ _03710_ sub1.data_o\[79\] vssd1 vssd1 vccd1 vccd1
+ _03719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12798_ fifo_bank_register.bank\[2\]\[62\] _05401_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07699_ sky130_fd_sc_hd__mux2_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _02864_ fifo_bank_register.data_out\[108\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02865_ sky130_fd_sc_hd__mux2_1
X_17325_ net464 _00768_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
X_11749_ _07144_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17256_ net418 _00699_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
X_14468_ fifo_bank_register.bank\[1\]\[100\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[100\]
+ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_226_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13419_ _07937_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16207_ _04153_ _04154_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__xor2_4
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17187_ net402 _00630_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14399_ fifo_bank_register.bank\[5\]\[93\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[93\]
+ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16138_ net150 ks1.key_reg\[118\] _03976_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08960_ _04684_ _04982_ _04983_ _04689_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16069_ _04028_ _04029_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__xor2_4
XFILLER_0_227_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_5_clk clknet_3_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08891_ ks1.key_reg\[16\] _04726_ _04914_ net165 vssd1 vssd1 vccd1 vccd1 _04915_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_202_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09512_ fifo_bank_register.bank\[9\]\[79\] _05436_ _05418_ vssd1 vssd1 vccd1 vccd1
+ _05437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09443_ net210 vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_177_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09374_ _05343_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08325_ _04475_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__buf_2
XFILLER_0_157_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08256_ _04409_ _04410_ _04411_ _04412_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__or4_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput260 net260 vssd1 vssd1 vccd1 vccd1 data_o[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput271 net271 vssd1 vssd1 vccd1 vccd1 data_o[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput282 net282 vssd1 vssd1 vccd1 vccd1 data_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_203_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10080_ sub1.data_o\[33\] _05753_ _05904_ _05905_ _04611_ vssd1 vssd1 vccd1 vccd1
+ _05906_ sky130_fd_sc_hd__a221o_1
Xoutput293 net293 vssd1 vssd1 vccd1 vccd1 data_o[14] sky130_fd_sc_hd__buf_2
XTAP_5914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_214_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13770_ fifo_bank_register.bank\[5\]\[24\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[24\]
+ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10982_ net154 ks1.key_reg\[121\] _06579_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__mux2_1
X_12721_ _07658_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15440_ _03626_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_214_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_194_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ fifo_bank_register.bank\[3\]\[122\] _05526_ _07485_ vssd1 vssd1 vccd1 vccd1
+ _07621_ sky130_fd_sc_hd__mux2_1
XFILLER_0_167_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11603_ fifo_bank_register.bank\[6\]\[10\] _05290_ _07067_ vssd1 vssd1 vccd1 vccd1
+ _07068_ sky130_fd_sc_hd__mux2_1
X_15371_ _04368_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_148_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ fifo_bank_register.bank\[3\]\[89\] _05457_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17110_ net496 _00553_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14322_ _02673_ fifo_bank_register.data_out\[84\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18090_ net456 _01533_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[92\]
+ sky130_fd_sc_hd__dfxtp_2
X_11534_ fifo_bank_register.bank\[7\]\[106\] _05493_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17041_ net543 _00484_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14253_ fifo_bank_register.bank\[9\]\[77\] _02550_ _02609_ _02610_ _02611_ vssd1
+ vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_184_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11465_ fifo_bank_register.bank\[7\]\[73\] _05424_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _06995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13204_ fifo_bank_register.bank\[1\]\[127\] _05536_ _07771_ vssd1 vssd1 vccd1 vccd1
+ _07912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10416_ mix1.data_o\[65\] _06138_ _06162_ _06163_ sub1.data_o\[65\] vssd1 vssd1 vccd1
+ vccd1 _06210_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14184_ _02136_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_180_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11396_ fifo_bank_register.bank\[7\]\[40\] _05354_ _06958_ vssd1 vssd1 vccd1 vccd1
+ _06959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13135_ _07876_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__clkbuf_1
X_10347_ _06147_ _06148_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17943_ net565 _01386_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[81\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _07840_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_225_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10278_ _06084_ _06085_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12017_ fifo_bank_register.bank\[5\]\[78\] _05434_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1064 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17874_ net500 _01317_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16825_ clknet_leaf_8_clk _00269_ net632 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[116\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_206_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16756_ clknet_leaf_66_clk _00200_ net604 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[47\]
+ sky130_fd_sc_hd__dfrtp_4
X_13968_ fifo_bank_register.bank\[5\]\[46\] _02309_ _02310_ fifo_bank_register.bank\[3\]\[46\]
+ vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_159_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15707_ mix1.data_o\[56\] net756 _03775_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12919_ fifo_bank_register.bank\[2\]\[120\] _05522_ _07628_ vssd1 vssd1 vccd1 vccd1
+ _07762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13899_ fifo_bank_register.bank\[0\]\[38\] _02296_ _02239_ vssd1 vssd1 vccd1 vccd1
+ _02297_ sky130_fd_sc_hd__mux2_1
X_16687_ net443 _00135_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18426_ clknet_leaf_0_clk _01856_ net620 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[111\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_61_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15638_ mix1.data_o\[23\] _03510_ _03742_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_174_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18357_ clknet_leaf_84_clk _01787_ net581 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[42\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15569_ _04713_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17308_ net536 _00751_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[86\]
+ sky130_fd_sc_hd__dfxtp_1
X_09090_ _05068_ _05101_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__xnor2_1
X_18288_ clknet_leaf_26_clk _01719_ net649 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[54\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17239_ net497 _00682_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09992_ addroundkey_data_o\[23\] _05827_ _05793_ vssd1 vssd1 vccd1 vccd1 _05828_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08943_ _04923_ _04966_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_228_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08874_ addroundkey_data_o\[40\] _04693_ _04695_ addroundkey_data_o\[32\] vssd1 vssd1
+ vccd1 vccd1 _04898_ sky130_fd_sc_hd__a22o_1
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_220_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09426_ fifo_bank_register.bank\[9\]\[51\] _05378_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_176_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09357_ fifo_bank_register.bank\[9\]\[29\] _05331_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08308_ _04449_ _04454_ _04459_ _04464_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__or4_2
XFILLER_0_133_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09288_ fifo_bank_register.bank\[9\]\[7\] _05284_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_209_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ net70 net69 net72 net71 vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__or4_1
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11250_ _05480_ fifo_bank_register.bank\[8\]\[100\] _06880_ vssd1 vssd1 vccd1 vccd1
+ _06881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10201_ _06016_ vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11181_ _06844_ vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_219_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ sub1.data_o\[37\] _05753_ _05951_ _05953_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _05954_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10063_ sub1.data_o\[32\] _05889_ _05751_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__mux2_1
X_14940_ addroundkey_data_o\[96\] _03056_ _03214_ vssd1 vssd1 vccd1 vccd1 _03215_
+ sky130_fd_sc_hd__a21oi_2
XTAP_5744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14871_ sub1.data_o\[8\] _04379_ _03059_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_
+ sky130_fd_sc_hd__a211o_1
XTAP_5799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16610_ net557 _00058_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13822_ _02140_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__clkbuf_4
X_17590_ net412 _01033_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[112\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16541_ net706 _03537_ _03143_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__mux2_1
X_13753_ _02167_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__clkbuf_1
X_10965_ _05623_ _06700_ _06704_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ fifo_bank_register.bank\[2\]\[18\] _05307_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13684_ _02104_ fifo_bank_register.data_out\[15\] _08172_ vssd1 vssd1 vccd1 vccd1
+ _02105_ sky130_fd_sc_hd__mux2_1
X_16472_ _04319_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10896_ _06491_ _06640_ _06641_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18211_ clknet_leaf_12_clk _01642_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_222_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15423_ sub1.data_o\[19\] _03606_ _03615_ _03611_ vssd1 vssd1 vccd1 vccd1 _03616_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_182_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_167_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ _07612_ vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15354_ net742 _03527_ _03560_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18142_ clknet_leaf_53_clk sbox1.ah\[0\] net656 vssd1 vssd1 vccd1 vccd1 sbox1.ah_reg\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_939 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12566_ _07576_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11517_ fifo_bank_register.bank\[7\]\[98\] _05476_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07022_ sky130_fd_sc_hd__mux2_1
X_14305_ fifo_bank_register.bank\[0\]\[82\] _02658_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02659_ sky130_fd_sc_hd__mux2_1
X_15285_ _03124_ _03416_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_135_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18073_ net555 _01516_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12497_ fifo_bank_register.bank\[3\]\[48\] _05371_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14236_ fifo_bank_register.bank\[1\]\[75\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[75\]
+ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
X_17024_ net557 _00467_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11448_ fifo_bank_register.bank\[7\]\[65\] _05407_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ fifo_bank_register.bank\[5\]\[68\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[68\]
+ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11379_ fifo_bank_register.bank\[7\]\[32\] _05338_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _07867_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__clkbuf_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14098_ fifo_bank_register.bank\[7\]\[60\] _02461_ _02470_ fifo_bank_register.bank\[2\]\[60\]
+ _02473_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a221o_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ net512 _01369_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[64\]
+ sky130_fd_sc_hd__dfxtp_1
X_13049_ _07831_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17857_ net439 _01300_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[123\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16808_ clknet_leaf_4_clk _00252_ net591 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[99\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_206_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08590_ _04615_ _04616_ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__mux2_4
X_17788_ net570 _01231_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16739_ clknet_leaf_47_clk _00183_ net653 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09211_ sub1.data_o\[116\] _05197_ _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18409_ clknet_leaf_10_clk _01839_ net623 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[94\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_174_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09142_ _05145_ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09073_ _05084_ _05086_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_198_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09975_ mix1.data_o\[22\] _05797_ _05703_ _05704_ sub1.data_o\[22\] vssd1 vssd1 vccd1
+ vccd1 _05812_ sky130_fd_sc_hd__a32o_1
XTAP_5007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08926_ _04946_ _04947_ _04948_ _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__a22o_1
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08857_ addroundkey_data_o\[16\] mix1.data_o\[16\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04881_ sky130_fd_sc_hd__mux2_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08788_ addroundkey_data_o\[59\] mix1.data_o\[59\] _04805_ vssd1 vssd1 vccd1 vccd1
+ _04812_ sky130_fd_sc_hd__mux2_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _06510_ vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ net198 vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10681_ sub1.data_o\[92\] _06447_ _06318_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12420_ _07499_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ _05497_ fifo_bank_register.bank\[4\]\[108\] _07453_ vssd1 vssd1 vccd1 vccd1
+ _07462_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11302_ _06907_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15070_ addroundkey_data_o\[116\] _03057_ _03341_ vssd1 vssd1 vccd1 vccd1 _03342_
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12282_ _05428_ fifo_bank_register.bank\[4\]\[75\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07426_ sky130_fd_sc_hd__mux2_1
X_14021_ fifo_bank_register.bank\[6\]\[51\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[51\]
+ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ _05464_ fifo_bank_register.bank\[8\]\[92\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11164_ _06835_ vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10115_ _05913_ _05754_ sub1.data_o\[36\] _05902_ vssd1 vssd1 vccd1 vccd1 _05938_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ _06799_ vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__clkbuf_1
X_15972_ ks1.col\[4\] _03942_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__xor2_4
XTAP_5541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17711_ net467 _01154_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14923_ _03180_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__xnor2_4
X_10046_ sub1.data_o\[30\] _05874_ _05819_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__mux2_1
XTAP_5574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_216_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold70 mix1.data_reg\[53\] vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_203_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_175_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold81 mix1.data_reg\[106\] vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 mix1.data_reg\[38\] vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ net422 _01085_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[36\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_4873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14854_ addroundkey_data_o\[101\] _03055_ _03129_ vssd1 vssd1 vccd1 vccd1 _03130_
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_89_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13805_ fifo_bank_register.bank\[6\]\[28\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_188_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17573_ net400 _01016_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[95\]
+ sky130_fd_sc_hd__dfxtp_1
X_14785_ mix1.state\[0\] _03060_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__and2_2
X_11997_ _07275_ vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16524_ _04346_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__clkbuf_1
X_10948_ net21 mix1.data_o\[118\] _05602_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__mux2_1
X_13736_ _02151_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16455_ _04308_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__clkbuf_1
X_13667_ fifo_bank_register.bank\[0\]\[13\] _02089_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02090_ sky130_fd_sc_hd__mux2_1
X_10879_ addroundkey_data_o\[111\] _06626_ _06612_ vssd1 vssd1 vccd1 vccd1 _06627_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15406_ sub1.data_o\[78\] _03600_ _03595_ sub1.data_o\[14\] vssd1 vssd1 vccd1 vccd1
+ _03604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12618_ _07603_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__clkbuf_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ fifo_bank_register.bank\[9\]\[6\] _08090_ _08160_ _08161_ _08162_ vssd1 vssd1
+ vccd1 vccd1 _08163_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _04270_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18125_ net442 _01568_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[127\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15337_ _03561_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12549_ _07567_ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18056_ net557 _01499_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[58\]
+ sky130_fd_sc_hd__dfxtp_1
X_15268_ _03207_ _03273_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17007_ net389 _00450_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14219_ fifo_bank_register.bank\[6\]\[73\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[73\]
+ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15199_ _03420_ _03461_ _04617_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout508 net509 vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_2
Xfanout519 net520 vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_226_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09760_ _04625_ _05616_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__nand2_4
XFILLER_0_225_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08711_ _04724_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__buf_4
XFILLER_0_207_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17909_ net396 _01352_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[47\]
+ sky130_fd_sc_hd__dfxtp_1
X_09691_ sub1.data_o\[122\] _05560_ _04891_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_193_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08642_ _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__buf_4
XFILLER_0_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_179_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08573_ _04605_ vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_174_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09125_ _05128_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_165_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _04966_ _05055_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__nor2_1
XFILLER_0_170_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09958_ _05676_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__clkbuf_4
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ addroundkey_data_o\[117\] mix1.data_o\[117\] _04702_ vssd1 vssd1 vccd1 vccd1
+ _04933_ sky130_fd_sc_hd__mux2_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _05734_ vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__clkbuf_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _07235_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_169_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ mix1.data_o\[103\] _06494_ _06398_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14570_ fifo_bank_register.bank\[0\]\[111\] _02894_ _02887_ vssd1 vssd1 vccd1 vccd1
+ _02895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ fifo_bank_register.bank\[6\]\[95\] _05470_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10733_ mix1.data_o\[97\] _06494_ _06398_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__o21a_1
X_13521_ _08091_ vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ _08043_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__clkbuf_1
X_16240_ _04183_ _04184_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10664_ net118 mix1.data_o\[90\] _06316_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12403_ _07490_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16171_ _04918_ _04121_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__xnor2_1
X_13383_ _08007_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__clkbuf_1
X_10595_ _06370_ vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_180_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15122_ _03140_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__xor2_4
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12334_ _07364_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__buf_4
XFILLER_0_50_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15053_ _03325_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12265_ _05411_ fifo_bank_register.bank\[4\]\[67\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14004_ _02140_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11216_ _05447_ fifo_bank_register.bank\[8\]\[84\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06863_ sky130_fd_sc_hd__mux2_1
X_12196_ _05342_ fifo_bank_register.bank\[4\]\[34\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_6050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11147_ _05378_ fifo_bank_register.bank\[8\]\[51\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06827_ sky130_fd_sc_hd__mux2_1
XTAP_6061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11078_ _05309_ fifo_bank_register.bank\[8\]\[19\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06790_ sky130_fd_sc_hd__mux2_1
X_15955_ _03926_ _03927_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__xor2_1
XFILLER_0_223_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput160 key_i[127] vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_4
XFILLER_0_216_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput171 key_i[21] vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_4
XTAP_5393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14906_ sub1.data_o\[87\] _03062_ _03091_ sub1.data_o\[55\] vssd1 vssd1 vccd1 vccd1
+ _03181_ sky130_fd_sc_hd__a22o_1
X_10029_ sub1.data_o\[28\] _05859_ _05819_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__mux2_1
Xinput182 key_i[31] vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xinput193 key_i[41] vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_4
X_15886_ sub1.data_o\[96\] _03874_ _03876_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__mux2_1
XTAP_4670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17625_ net501 _01068_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
X_14837_ addroundkey_data_o\[21\] _04376_ _05606_ _03112_ vssd1 vssd1 vccd1 vccd1
+ _03113_ sky130_fd_sc_hd__a211o_1
XFILLER_0_188_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17556_ net517 _00999_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
X_14768_ ks1.col\[20\] _05217_ _00007_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16507_ _04337_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13719_ _02135_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__clkbuf_1
X_17487_ net480 _00930_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14699_ fifo_bank_register.bank\[0\]\[127\] _03007_ _08120_ vssd1 vssd1 vccd1 vccd1
+ _03008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16438_ _04299_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16369_ _04260_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18108_ net470 _01551_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[110\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039_ net399 _01482_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[41\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09812_ _05665_ vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_185_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09743_ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09674_ _05152_ _05242_ _05060_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_193_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_179_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08625_ _04624_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__nand2_4
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08556_ addroundkey_data_o\[116\] fifo_bank_register.data_out\[116\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__mux2_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08487_ addroundkey_data_o\[83\] fifo_bank_register.data_out\[83\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_175_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_165_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_220_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09108_ _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__buf_2
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10380_ addroundkey_data_o\[60\] _06178_ _06169_ vssd1 vssd1 vccd1 vccd1 _06179_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_1276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09039_ _04967_ _05054_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12050_ _07303_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11001_ _06736_ vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15740_ _03800_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__clkbuf_1
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12952_ fifo_bank_register.bank\[1\]\[7\] _05284_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07780_ sky130_fd_sc_hd__mux2_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _07226_ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__clkbuf_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _03741_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__buf_4
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _07743_ vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__clkbuf_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_185_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17410_ net515 _00853_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_232 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ fifo_bank_register.bank\[5\]\[118\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[118\]
+ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__a22o_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_243 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18390_ clknet_leaf_84_clk _01820_ net619 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[75\]
+ sky130_fd_sc_hd__dfrtp_4
X_11834_ fifo_bank_register.bank\[6\]\[120\] _05522_ _07055_ vssd1 vssd1 vccd1 vccd1
+ _07189_ sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_265 _04490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_276 addroundkey_data_o\[23\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_287 sub1.data_o\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17341_ net429 _00784_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_298 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14553_ fifo_bank_register.bank\[7\]\[110\] _02866_ _02875_ fifo_bank_register.bank\[2\]\[110\]
+ _02878_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__a221o_1
X_11765_ fifo_bank_register.bank\[6\]\[87\] _05453_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07153_ sky130_fd_sc_hd__mux2_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ sub1.data_o\[96\] _06477_ _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13504_ _05262_ _08064_ _08080_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17272_ net555 _00715_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11696_ fifo_bank_register.bank\[6\]\[54\] _05384_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07117_ sky130_fd_sc_hd__mux2_1
X_14484_ fifo_bank_register.bank\[6\]\[102\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[102\]
+ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16223_ _04748_ _04169_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ sub1.data_o\[88\] _06417_ _06318_ vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__mux2_1
X_13435_ _08034_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13366_ _07998_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__clkbuf_1
X_16154_ _03957_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__buf_4
X_10578_ mix1.data_o\[82\] _06129_ _06093_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15105_ _03374_ _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12317_ _07444_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13297_ _07962_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__clkbuf_1
X_16085_ ks1.col\[16\] _04043_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ sub1.data_o\[27\] _04378_ _03059_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12248_ _05394_ fifo_bank_register.bank\[4\]\[59\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_220_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12179_ _05325_ fifo_bank_register.bank\[4\]\[26\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16987_ net483 _00430_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_208_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15938_ _04920_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__or2_1
XFILLER_0_190_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_210_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15869_ sub1.data_o\[89\] _05553_ _04888_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_203_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08410_ _04520_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_188_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17608_ net475 _01051_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ net192 vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__buf_2
X_18588_ clknet_leaf_74_clk _02017_ net588 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_176_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08341_ _04484_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_19_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17539_ net526 _00982_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08272_ net147 net146 net149 net148 vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_229_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_172_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_227_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09726_ _04614_ _05575_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09657_ fifo_bank_register.bank\[9\]\[126\] _05534_ _05269_ vssd1 vssd1 vccd1 vccd1
+ _05535_ sky130_fd_sc_hd__mux2_1
XFILLER_0_222_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ round\[0\] addroundkey_round\[0\] vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__xor2_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09588_ _05488_ vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_195_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08539_ addroundkey_data_o\[108\] fifo_bank_register.data_out\[108\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__mux2_2
XFILLER_0_195_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_194_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_182_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11550_ _07039_ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10501_ addroundkey_data_o\[74\] _06285_ _06248_ vssd1 vssd1 vccd1 vccd1 _06286_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11481_ _07003_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _07921_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10432_ sub1.data_o\[67\] _06223_ _06160_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13151_ fifo_bank_register.bank\[1\]\[101\] _05483_ _07883_ vssd1 vssd1 vccd1 vccd1
+ _07885_ sky130_fd_sc_hd__mux2_1
X_10363_ _05620_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12102_ _07330_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13082_ _07848_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__clkbuf_1
X_10294_ _06100_ vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12033_ _07294_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__clkbuf_1
X_16910_ net555 _00353_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[72\]
+ sky130_fd_sc_hd__dfxtp_1
X_17890_ net485 _01333_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ net420 _00284_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16772_ clknet_leaf_47_clk _00216_ net651 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[63\]
+ sky130_fd_sc_hd__dfrtp_4
X_13984_ _02372_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18511_ clknet_leaf_62_clk _01940_ net598 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[38\]
+ sky130_fd_sc_hd__dfrtp_1
X_15723_ _03791_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__clkbuf_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12935_ _05267_ _07483_ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__and2_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ clknet_leaf_1_clk _01872_ net620 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[127\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _03755_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__clkbuf_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _07734_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14605_ fifo_bank_register.bank\[5\]\[116\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[116\]
+ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__a22o_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18373_ clknet_leaf_37_clk _01803_ net668 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[58\]
+ sky130_fd_sc_hd__dfrtp_4
X_11817_ _07180_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__clkbuf_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _03717_ _03709_ _05236_ _03718_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a31o_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12797_ _07698_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ net464 _00767_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[102\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ fifo_bank_register.bank\[0\]\[108\] _02863_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02864_ sky130_fd_sc_hd__mux2_1
X_11748_ fifo_bank_register.bank\[6\]\[79\] _05436_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17255_ net424 _00698_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[33\]
+ sky130_fd_sc_hd__dfxtp_1
X_14467_ _02153_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_183_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11679_ fifo_bank_register.bank\[6\]\[46\] _05367_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16206_ net156 ks1.key_reg\[123\] _04742_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__mux2_2
XFILLER_0_113_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13418_ _08025_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__clkbuf_1
X_17186_ net410 _00629_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14398_ _02741_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16137_ net698 _03901_ _04089_ _04090_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a22o_1
X_13349_ _07989_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_224_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16068_ net233 ks1.key_reg\[78\] _03907_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__mux2_2
XFILLER_0_110_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15019_ sub1.data_o\[19\] _03208_ _03081_ _03291_ vssd1 vssd1 vccd1 vccd1 _03292_
+ sky130_fd_sc_hd__a211o_1
X_08890_ ks1.key_reg\[16\] _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__or3_1
XFILLER_0_202_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_196_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09511_ net234 vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__buf_2
XFILLER_0_211_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09442_ _05389_ vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_182_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_177_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09373_ fifo_bank_register.bank\[9\]\[34\] _05342_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_177_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08324_ addroundkey_data_o\[6\] fifo_bank_register.data_out\[6\] _04468_ vssd1 vssd1
+ vccd1 vccd1 _04475_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08255_ net110 net109 net112 net111 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_172_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_203_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_203_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput261 net261 vssd1 vssd1 vccd1 vccd1 data_o[100] sky130_fd_sc_hd__clkbuf_4
Xoutput272 net272 vssd1 vssd1 vccd1 vccd1 data_o[110] sky130_fd_sc_hd__buf_2
XFILLER_0_218_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput283 net283 vssd1 vssd1 vccd1 vccd1 data_o[120] sky130_fd_sc_hd__clkbuf_4
Xoutput294 net294 vssd1 vssd1 vccd1 vccd1 data_o[15] sky130_fd_sc_hd__clkbuf_4
XTAP_5904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_5926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_173_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _04613_ _04627_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10981_ _06583_ _06717_ _06718_ _06587_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__a22o_1
XFILLER_0_214_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12720_ fifo_bank_register.bank\[2\]\[25\] _05323_ _07652_ vssd1 vssd1 vccd1 vccd1
+ _07658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_210_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12651_ _07620_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_214_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ _07055_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__buf_4
X_15370_ sub1.data_o\[34\] sub1.data_o\[98\] _03574_ vssd1 vssd1 vccd1 vccd1 _03580_
+ sky130_fd_sc_hd__mux2_1
X_12582_ _07584_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14321_ fifo_bank_register.bank\[0\]\[84\] _02672_ _02644_ vssd1 vssd1 vccd1 vccd1
+ _02673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11533_ _07030_ vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17040_ net546 _00483_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_1295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14252_ fifo_bank_register.bank\[1\]\[77\] _02559_ _02560_ fifo_bank_register.bank\[8\]\[77\]
+ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__a22o_1
X_11464_ _06994_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ sub1.data_o\[65\] _06208_ _06160_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__mux2_1
X_13203_ _07911_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11395_ _06935_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__buf_4
X_14183_ _02549_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_221_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13134_ fifo_bank_register.bank\[1\]\[93\] _05466_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07876_ sky130_fd_sc_hd__mux2_1
X_10346_ net210 ks1.key_reg\[57\] _05997_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ net566 _01385_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[80\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ fifo_bank_register.bank\[1\]\[60\] _05396_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07840_ sky130_fd_sc_hd__mux2_1
X_10277_ net204 ks1.key_reg\[51\] _05920_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__mux2_4
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12016_ _07285_ vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_224_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17873_ net533 _01316_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[11\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_217_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16824_ clknet_leaf_29_clk _00268_ net635 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_219_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16755_ clknet_leaf_66_clk _00199_ net603 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[46\]
+ sky130_fd_sc_hd__dfrtp_4
X_13967_ _02357_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15706_ _03782_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__clkbuf_1
X_12918_ _07761_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16686_ net495 _00134_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[126\]
+ sky130_fd_sc_hd__dfxtp_1
X_13898_ fifo_bank_register.bank\[9\]\[38\] _02226_ _02293_ _02294_ _02295_ vssd1
+ vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18425_ clknet_leaf_3_clk _01855_ net583 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[110\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_119_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15637_ _03746_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__clkbuf_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_159_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12849_ _07725_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__clkbuf_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18356_ clknet_leaf_12_clk _01786_ net621 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[41\]
+ sky130_fd_sc_hd__dfrtp_4
X_15568_ _03700_ _04935_ _05245_ _03708_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a31o_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17307_ net540 _00750_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[85\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_946 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14519_ fifo_bank_register.bank\[0\]\[106\] _02848_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02849_ sky130_fd_sc_hd__mux2_1
X_18287_ clknet_leaf_26_clk _01718_ net649 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[53\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15499_ _04369_ _04777_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17238_ net493 _00681_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17169_ net552 _00612_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09991_ _05824_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ _04648_ _04955_ _04965_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08873_ mix1.data_o\[40\] _04693_ _04695_ mix1.data_o\[32\] vssd1 vssd1 vccd1 vccd1
+ _04897_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_212_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09425_ net204 vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__buf_2
XFILLER_0_192_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09356_ net179 vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__buf_2
XFILLER_0_118_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08307_ _04460_ _04461_ _04462_ _04463_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__or4_1
X_09287_ net235 vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08238_ net61 net60 net64 net63 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10200_ addroundkey_data_o\[43\] _06015_ _05980_ vssd1 vssd1 vccd1 vccd1 _06016_
+ sky130_fd_sc_hd__mux2_1
X_11180_ _05411_ fifo_bank_register.bank\[8\]\[67\] _06836_ vssd1 vssd1 vccd1 vccd1
+ _06844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_197_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10131_ mix1.data_o\[37\] _05952_ _05916_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__o21a_1
XTAP_5701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_206_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10062_ net54 mix1.data_o\[32\] _05749_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14870_ sub1.data_o\[72\] _03144_ _03145_ sub1.data_o\[40\] vssd1 vssd1 vccd1 vccd1
+ _03146_ sky130_fd_sc_hd__a22o_1
XTAP_5789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_216_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13821_ _02138_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16540_ _04354_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_168_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13752_ _02166_ fifo_bank_register.data_out\[21\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10964_ sub1.data_o\[119\] _05613_ _06702_ _06703_ _04610_ vssd1 vssd1 vccd1 vccd1
+ _06704_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12703_ _07648_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__clkbuf_1
X_16471_ net849 _04318_ _03957_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ fifo_bank_register.bank\[0\]\[15\] _02103_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02104_ sky130_fd_sc_hd__mux2_1
X_10895_ _06630_ _06514_ sub1.data_o\[113\] _05675_ vssd1 vssd1 vccd1 vccd1 _06641_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18210_ clknet_leaf_14_clk _01641_ net629 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[40\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15422_ sub1.data_o\[115\] sub1.data_o\[51\] _03609_ vssd1 vssd1 vccd1 vccd1 _03615_
+ sky130_fd_sc_hd__mux2_1
X_12634_ fifo_bank_register.bank\[3\]\[113\] _05508_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18141_ clknet_leaf_53_clk sbox1.next_alph\[3\] net657 vssd1 vssd1 vccd1 vccd1 sbox1.alph\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_15353_ _03569_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12565_ fifo_bank_register.bank\[3\]\[80\] _05438_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_182_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14304_ fifo_bank_register.bank\[9\]\[82\] _02631_ _02655_ _02656_ _02657_ vssd1
+ vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a2111o_1
X_11516_ _07021_ vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18072_ net549 _01515_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[74\]
+ sky130_fd_sc_hd__dfxtp_2
X_15284_ _03530_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_202_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ _07539_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17023_ net550 _00466_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14235_ fifo_bank_register.bank\[6\]\[75\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[75\]
+ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
XFILLER_0_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11447_ _06985_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11378_ _06949_ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__clkbuf_1
X_14166_ _02534_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13117_ fifo_bank_register.bank\[1\]\[85\] _05449_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07867_ sky130_fd_sc_hd__mux2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ net208 ks1.key_reg\[55\] _06097_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__mux2_4
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ fifo_bank_register.bank\[5\]\[60\] _02471_ _02472_ fifo_bank_register.bank\[3\]\[60\]
+ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__a22o_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ net524 _01368_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_13048_ fifo_bank_register.bank\[1\]\[52\] _05380_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_206_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17856_ net493 _01299_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[122\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16807_ clknet_leaf_74_clk _00251_ net591 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[98\]
+ sky130_fd_sc_hd__dfrtp_4
X_17787_ net562 _01230_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[53\]
+ sky130_fd_sc_hd__dfxtp_1
X_14999_ _03269_ _03272_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__nor2_4
XFILLER_0_156_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16738_ clknet_leaf_51_clk _00182_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16669_ net458 _00117_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_220_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_202_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09210_ sub1.data_o\[20\] _05200_ _05203_ sub1.data_o\[84\] vssd1 vssd1 vccd1 vccd1
+ _05220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18408_ clknet_leaf_10_clk _01838_ net623 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[93\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ _05148_ _05151_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_134_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18339_ clknet_leaf_35_clk _01769_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_173_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09072_ _05058_ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09974_ sub1.data_o\[22\] _05810_ _05701_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08925_ _04710_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_228_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08856_ _04805_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__buf_4
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08787_ addroundkey_data_o\[11\] mix1.data_o\[11\] _04665_ vssd1 vssd1 vccd1 vccd1
+ _04811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09408_ _05366_ vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__clkbuf_1
X_10680_ net120 mix1.data_o\[92\] _06316_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_211_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ fifo_bank_register.bank\[9\]\[23\] _05319_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ _07461_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11301_ _05532_ fifo_bank_register.bank\[8\]\[125\] _06768_ vssd1 vssd1 vccd1 vccd1
+ _06907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12281_ _07425_ vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11232_ _06871_ vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__clkbuf_1
X_14020_ fifo_bank_register.bank\[7\]\[51\] _02380_ _02389_ fifo_bank_register.bank\[2\]\[51\]
+ _02404_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a221o_1
XFILLER_0_181_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11163_ _05394_ fifo_bank_register.bank\[8\]\[59\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10114_ sub1.data_o\[36\] _05935_ _05936_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__mux2_1
XTAP_5520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11094_ _05325_ fifo_bank_register.bank\[8\]\[26\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06799_ sky130_fd_sc_hd__mux2_1
X_15971_ net131 ks1.key_reg\[100\] _03905_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__mux2_2
XFILLER_0_207_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17710_ net462 _01153_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14922_ _03188_ _03196_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__xor2_2
X_10045_ net52 mix1.data_o\[30\] _05817_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__mux2_1
XTAP_5564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold60 mix1.data_reg\[46\] vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold71 mix1.data_reg\[48\] vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold82 mix1.data_reg\[90\] vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17641_ net416 _01084_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14853_ addroundkey_data_o\[5\] _03100_ _05606_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_
+ sky130_fd_sc_hd__a211o_1
Xhold93 mix1.data_reg\[51\] vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_188_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_165_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13804_ fifo_bank_register.bank\[7\]\[28\] _02128_ _02139_ fifo_bank_register.bank\[2\]\[28\]
+ _02211_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a221o_1
X_17572_ net448 _01015_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_203_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14784_ mix1.state\[1\] vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__inv_2
X_11996_ fifo_bank_register.bank\[5\]\[68\] _05413_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16523_ net779 _03507_ _04343_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13735_ _08110_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__buf_6
XFILLER_0_202_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10947_ _06688_ vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_196_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16454_ ks1.key_reg\[121\] _04307_ _03957_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_195_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13666_ fifo_bank_register.bank\[9\]\[13\] _08190_ _02086_ _02087_ _02088_ vssd1
+ vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_112_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10878_ _06624_ _06625_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__xor2_1
XFILLER_0_171_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15405_ _05103_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__clkbuf_4
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12617_ fifo_bank_register.bank\[3\]\[105\] _05491_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07603_ sky130_fd_sc_hd__mux2_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ ks1.key_reg\[90\] _04269_ _04264_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_213_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13597_ fifo_bank_register.bank\[1\]\[6\] _08112_ _08115_ fifo_bank_register.bank\[8\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _08162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_171_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18124_ net531 _01567_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[126\]
+ sky130_fd_sc_hd__dfxtp_1
X_15336_ net763 _03497_ _03560_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12548_ fifo_bank_register.bank\[3\]\[72\] _05422_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18055_ net549 _01498_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[57\]
+ sky130_fd_sc_hd__dfxtp_1
X_15267_ _03517_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__clkbuf_1
X_12479_ _07530_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 _02138_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17006_ net392 _00449_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[40\]
+ sky130_fd_sc_hd__dfxtp_1
X_14218_ fifo_bank_register.bank\[7\]\[73\] _02542_ _02551_ fifo_bank_register.bank\[2\]\[73\]
+ _02580_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__a221o_1
X_15198_ _03459_ _03460_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14149_ _02519_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__clkbuf_1
Xfanout509 net510 vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08710_ ks1.key_reg\[4\] _04726_ _04733_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__a21oi_1
X_17908_ net390 _01351_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[46\]
+ sky130_fd_sc_hd__dfxtp_1
X_09690_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__buf_4
X_08641_ _04655_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__buf_4
X_17839_ net468 _01282_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[105\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08572_ addroundkey_data_o\[124\] fifo_bank_register.data_out\[124\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__mux2_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09124_ sbox1.alph\[2\] _05134_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_228_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ sbox1.ah\[1\] _05071_ vssd1 vssd1 vccd1 vccd1 sbox1.next_alph\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_26_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_217_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_204_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09957_ sub1.data_o\[20\] _05795_ _05701_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ addroundkey_data_o\[85\] mix1.data_o\[85\] _04880_ vssd1 vssd1 vccd1 vccd1
+ _04932_ sky130_fd_sc_hd__mux2_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09888_ addroundkey_data_o\[13\] _05733_ _05697_ vssd1 vssd1 vccd1 vccd1 _05734_
+ sky130_fd_sc_hd__mux2_1
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08839_ _04721_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__inv_2
XFILLER_0_213_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _05267_ _06910_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _06491_ _06555_ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a21o_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_184_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11781_ _07161_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__clkbuf_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13520_ _05262_ _08056_ _08066_ vssd1 vssd1 vccd1 vccd1 _08091_ sky130_fd_sc_hd__nor3_1
XFILLER_0_83_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10732_ _04626_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13451_ _05512_ fifo_bank_register.bank\[0\]\[115\] _08037_ vssd1 vssd1 vccd1 vccd1
+ _08043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10663_ _06432_ vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_193_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ fifo_bank_register.bank\[3\]\[3\] _05276_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16170_ _04119_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__xor2_1
X_10594_ addroundkey_data_o\[83\] _06369_ _06327_ vssd1 vssd1 vccd1 vccd1 _06370_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_1260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13382_ _05443_ fifo_bank_register.bank\[0\]\[82\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08007_ sky130_fd_sc_hd__mux2_1
X_15121_ _03389_ _03390_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_180_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12333_ _07452_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15052_ mix1.data_reg\[67\] _03324_ _03171_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12264_ _07416_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14003_ _02138_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__clkbuf_4
X_11215_ _06862_ vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__clkbuf_1
X_12195_ _07380_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _06826_ vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__clkbuf_1
XTAP_6051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_208_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11077_ _06789_ vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__clkbuf_1
X_15954_ net220 ks1.key_reg\[66\] _03907_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__mux2_1
XTAP_6095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput150 key_i[118] vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__buf_4
XFILLER_0_218_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput161 key_i[12] vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_4
XTAP_5383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905_ _03107_ _03179_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__xnor2_4
X_10028_ net49 mix1.data_o\[28\] _05817_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__mux2_1
Xinput172 key_i[22] vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_4
XTAP_5394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_216_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15885_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__clkbuf_4
Xinput183 key_i[32] vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
Xinput194 key_i[42] vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_215_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_188_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14836_ addroundkey_data_o\[85\] _03108_ _03066_ addroundkey_data_o\[53\] vssd1 vssd1
+ vccd1 vccd1 _03112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17624_ net503 _01067_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[18\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ net544 _00998_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_169_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14767_ _03047_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11979_ _07221_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16506_ net711 _03477_ _04332_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__mux2_1
X_13718_ _02134_ fifo_bank_register.data_out\[19\] _02119_ vssd1 vssd1 vccd1 vccd1
+ _02135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17486_ net492 _00929_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14698_ fifo_bank_register.bank\[9\]\[127\] _08089_ _03004_ _03005_ _03006_ vssd1
+ vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_183_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16437_ net814 _04052_ _04295_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ fifo_bank_register.bank\[1\]\[11\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16368_ net808 _04070_ _04252_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18107_ net459 _01550_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[109\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_147_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15319_ net723 _03446_ _03549_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16299_ net833 _04064_ _04222_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ net415 _01481_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09811_ addroundkey_data_o\[5\] _05664_ next_addroundkey_ready_o vssd1 vssd1 vccd1
+ vccd1 _05665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_226_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09742_ _04624_ _04615_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09673_ _05152_ _05242_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_171_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08555_ _04596_ vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_166_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_193_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08486_ _04560_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_212_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09107_ _05113_ _05114_ _05115_ _05116_ _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_165_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09038_ _04971_ _05057_ vssd1 vssd1 vccd1 vccd1 sbox1.ah\[0\] sky130_fd_sc_hd__xor2_4
XFILLER_0_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_229_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11000_ addroundkey_data_o\[123\] _06735_ _05696_ vssd1 vssd1 vccd1 vccd1 _06736_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_229_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _07779_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__clkbuf_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11902_ fifo_bank_register.bank\[5\]\[23\] _05319_ _07222_ vssd1 vssd1 vccd1 vccd1
+ _07226_ sky130_fd_sc_hd__mux2_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15670_ _03763_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__clkbuf_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 net151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12882_ fifo_bank_register.bank\[2\]\[102\] _05485_ _07740_ vssd1 vssd1 vccd1 vccd1
+ _07743_ sky130_fd_sc_hd__mux2_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_212_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _02939_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__clkbuf_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_158_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11833_ _07188_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__clkbuf_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_255 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_266 _04501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_277 addroundkey_data_o\[39\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17340_ net408 _00783_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_200_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ fifo_bank_register.bank\[5\]\[110\] _02876_ _02877_ fifo_bank_register.bank\[3\]\[110\]
+ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a22o_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_288 sub1.data_o\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _07152_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_299 net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_172_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13503_ _08056_ _08075_ _08078_ _08079_ _08064_ vssd1 vssd1 vccd1 vccd1 _08080_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _05608_ vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__buf_4
X_17271_ net407 _00714_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14483_ fifo_bank_register.bank\[7\]\[102\] _02785_ _02794_ fifo_bank_register.bank\[2\]\[102\]
+ _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__a221o_1
X_11695_ _07116_ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16222_ _04167_ _04168_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__xor2_2
XFILLER_0_153_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ _05495_ fifo_bank_register.bank\[0\]\[107\] _08026_ vssd1 vssd1 vccd1 vccd1
+ _08034_ sky130_fd_sc_hd__mux2_1
X_10646_ net115 mix1.data_o\[88\] _06316_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_183_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_973 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ _05000_ _04104_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13365_ _05426_ fifo_bank_register.bank\[0\]\[74\] _07993_ vssd1 vssd1 vccd1 vccd1
+ _07998_ sky130_fd_sc_hd__mux2_1
X_10577_ _06126_ _06352_ _06353_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__a21o_1
XFILLER_0_183_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15104_ _03307_ _03352_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ _05462_ fifo_bank_register.bank\[4\]\[91\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07444_ sky130_fd_sc_hd__mux2_1
X_16084_ net144 ks1.key_reg\[112\] _03902_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_210_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13296_ _05357_ fifo_bank_register.bank\[0\]\[41\] _07960_ vssd1 vssd1 vccd1 vccd1
+ _07962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15035_ sub1.data_o\[91\] _03064_ _03068_ sub1.data_o\[59\] vssd1 vssd1 vccd1 vccd1
+ _03308_ sky130_fd_sc_hd__a22o_1
X_12247_ _07407_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_208_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12178_ _07371_ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11129_ _06817_ vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16986_ net508 _00429_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_194_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_218_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15937_ _03909_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__xor2_1
XTAP_5191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_161_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15868_ _03866_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_189_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14819_ sub1.data_o\[109\] _03078_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__a21oi_2
X_17607_ net492 _01050_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15799_ _03831_ vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__clkbuf_1
X_18587_ clknet_leaf_75_clk _02016_ net587 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_175_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08340_ addroundkey_data_o\[13\] fifo_bank_register.data_out\[13\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17538_ net513 _00981_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_191_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08271_ net143 net144 net145 net142 vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__or4bb_1
X_17469_ net435 _00912_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_229_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_172_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_162_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_229_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ _05585_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_179_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09656_ net159 vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__clkbuf_4
X_08607_ round\[1\] addroundkey_round\[1\] vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__xor2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ fifo_bank_register.bank\[9\]\[103\] _05487_ _05481_ vssd1 vssd1 vccd1 vccd1
+ _05488_ sky130_fd_sc_hd__mux2_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _04587_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08469_ _04551_ vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10500_ _06283_ _06284_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__xor2_1
XFILLER_0_163_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11480_ fifo_bank_register.bank\[7\]\[80\] _05438_ _07002_ vssd1 vssd1 vccd1 vccd1
+ _07003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_190_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10431_ net92 mix1.data_o\[67\] _06158_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13150_ _07884_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__clkbuf_1
X_10362_ _05757_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12101_ fifo_bank_register.bank\[5\]\[118\] _05518_ _07321_ vssd1 vssd1 vccd1 vccd1
+ _07330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_1373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10293_ addroundkey_data_o\[52\] _06099_ _06064_ vssd1 vssd1 vccd1 vccd1 _06100_
+ sky130_fd_sc_hd__mux2_1
X_13081_ fifo_bank_register.bank\[1\]\[68\] _05413_ _07839_ vssd1 vssd1 vccd1 vccd1
+ _07848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_218_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ fifo_bank_register.bank\[5\]\[85\] _05449_ _07288_ vssd1 vssd1 vccd1 vccd1
+ _07294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ net420 _00283_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_205_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout670 net259 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__buf_4
X_16771_ clknet_leaf_48_clk _00215_ net611 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[62\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13983_ _02370_ fifo_bank_register.data_out\[47\] _02371_ vssd1 vssd1 vccd1 vccd1
+ _02372_ sky130_fd_sc_hd__mux2_1
XFILLER_0_219_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15722_ mix1.data_o\[63\] mix1.data_reg\[63\] _03786_ vssd1 vssd1 vccd1 vccd1 _03791_
+ sky130_fd_sc_hd__mux2_1
X_18510_ clknet_leaf_62_clk _01939_ net600 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_12934_ _07769_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15653_ mix1.data_o\[30\] _03533_ _03753_ vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__mux2_1
X_18441_ clknet_leaf_1_clk _01871_ net624 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[126\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ fifo_bank_register.bank\[2\]\[94\] _05468_ _07729_ vssd1 vssd1 vccd1 vccd1
+ _07734_ sky130_fd_sc_hd__mux2_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_200_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_205_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _02924_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__clkbuf_1
X_18372_ clknet_leaf_37_clk _01802_ net667 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[57\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_185_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11816_ fifo_bank_register.bank\[6\]\[111\] _05504_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07180_ sky130_fd_sc_hd__mux2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15584_ sub1.data_o\[14\] _03660_ _03710_ sub1.data_o\[78\] vssd1 vssd1 vccd1 vccd1
+ _03718_ sky130_fd_sc_hd__a22o_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_200_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12796_ fifo_bank_register.bank\[2\]\[61\] _05399_ _07696_ vssd1 vssd1 vccd1 vccd1
+ _07698_ sky130_fd_sc_hd__mux2_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_157_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ net446 _00766_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[101\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_173_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ fifo_bank_register.bank\[9\]\[108\] _02793_ _02860_ _02861_ _02862_ vssd1
+ vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a2111o_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _07143_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17254_ net419 _00697_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[32\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14466_ _02151_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11678_ _07107_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16205_ ks1.col\[27\] _04152_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_226_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_183_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13417_ _05478_ fifo_bank_register.bank\[0\]\[99\] _08015_ vssd1 vssd1 vccd1 vccd1
+ _08025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17185_ net401 _00628_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10629_ _04638_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_221_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14397_ _02740_ fifo_bank_register.data_out\[92\] _02695_ vssd1 vssd1 vccd1 vccd1
+ _02741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16136_ _04957_ _04088_ _03914_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13348_ _05409_ fifo_bank_register.bank\[0\]\[66\] _07982_ vssd1 vssd1 vccd1 vccd1
+ _07989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16067_ _05235_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__xor2_4
XFILLER_0_122_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13279_ _05340_ fifo_bank_register.bank\[0\]\[33\] _07949_ vssd1 vssd1 vccd1 vccd1
+ _07953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_224_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15018_ sub1.data_o\[83\] _03209_ _03084_ sub1.data_o\[51\] vssd1 vssd1 vccd1 vccd1
+ _03291_ sky130_fd_sc_hd__a22o_1
XFILLER_0_209_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16969_ net475 _00412_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_224_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09510_ _05435_ vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09441_ fifo_bank_register.bank\[9\]\[56\] _05388_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09372_ net185 vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_192_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08323_ _04474_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08254_ net105 net104 net108 net107 vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_166_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_162_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput262 net262 vssd1 vssd1 vccd1 vccd1 data_o[101] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_203_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput273 net273 vssd1 vssd1 vccd1 vccd1 data_o[111] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput284 net284 vssd1 vssd1 vccd1 vccd1 data_o[121] sky130_fd_sc_hd__clkbuf_4
Xoutput295 net295 vssd1 vssd1 vccd1 vccd1 data_o[16] sky130_fd_sc_hd__clkbuf_4
XTAP_5905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_214_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09708_ _05198_ _04629_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10980_ mix1.data_o\[121\] _05676_ _06575_ _06576_ sub1.data_o\[121\] vssd1 vssd1
+ vccd1 vccd1 _06718_ sky130_fd_sc_hd__a32o_1
XFILLER_0_186_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09639_ fifo_bank_register.bank\[9\]\[120\] _05522_ _05269_ vssd1 vssd1 vccd1 vccd1
+ _05523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_168_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ fifo_bank_register.bank\[3\]\[121\] _05524_ _07485_ vssd1 vssd1 vccd1 vccd1
+ _07620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_210_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11601_ _07066_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ fifo_bank_register.bank\[3\]\[88\] _05455_ _07575_ vssd1 vssd1 vccd1 vccd1
+ _07584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ fifo_bank_register.bank\[9\]\[84\] _02631_ _02669_ _02670_ _02671_ vssd1
+ vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a2111o_1
X_11532_ fifo_bank_register.bank\[7\]\[105\] _05491_ _07024_ vssd1 vssd1 vccd1 vccd1
+ _07030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14251_ fifo_bank_register.bank\[6\]\[77\] _02556_ _02557_ fifo_bank_register.bank\[4\]\[77\]
+ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_184_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11463_ fifo_bank_register.bank\[7\]\[72\] _05422_ _06991_ vssd1 vssd1 vccd1 vccd1
+ _06994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_180_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13202_ fifo_bank_register.bank\[1\]\[126\] _05534_ _07771_ vssd1 vssd1 vccd1 vccd1
+ _07911_ sky130_fd_sc_hd__mux2_1
X_10414_ net90 mix1.data_o\[65\] _06158_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__mux2_1
X_14182_ _02548_ fifo_bank_register.data_out\[69\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02549_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11394_ _06957_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13133_ _07875_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__clkbuf_1
X_10345_ _06001_ _06145_ _06146_ _06005_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _07794_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__buf_4
X_17941_ net549 _01384_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[79\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_221_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_195_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10276_ _06076_ _06078_ _06083_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__o21ai_1
X_12015_ fifo_bank_register.bank\[5\]\[77\] _05432_ _07277_ vssd1 vssd1 vccd1 vccd1
+ _07285_ sky130_fd_sc_hd__mux2_1
X_17872_ net500 _01315_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[10\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_206_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16823_ clknet_leaf_8_clk _00267_ net633 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[114\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_205_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_191_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_206_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_215_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13966_ _02356_ fifo_bank_register.data_out\[45\] _02290_ vssd1 vssd1 vccd1 vccd1
+ _02357_ sky130_fd_sc_hd__mux2_1
X_16754_ clknet_leaf_64_clk _00198_ net603 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[45\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_191_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_221_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15705_ mix1.data_o\[55\] net734 _03775_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__mux2_1
X_12917_ fifo_bank_register.bank\[2\]\[119\] _05520_ _07751_ vssd1 vssd1 vccd1 vccd1
+ _07761_ sky130_fd_sc_hd__mux2_1
X_16685_ net497 _00133_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
X_13897_ fifo_bank_register.bank\[1\]\[38\] _02235_ _02236_ fifo_bank_register.bank\[8\]\[38\]
+ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18424_ clknet_leaf_83_clk _01854_ net584 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[109\]
+ sky130_fd_sc_hd__dfrtp_2
X_15636_ mix1.data_o\[22\] _03507_ _03742_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ fifo_bank_register.bank\[2\]\[86\] _05451_ _07718_ vssd1 vssd1 vccd1 vccd1
+ _07725_ sky130_fd_sc_hd__mux2_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_201_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15567_ sub1.data_o\[71\] _03691_ _03707_ _03594_ vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_174_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18355_ clknet_leaf_14_clk _01785_ net627 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[40\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ fifo_bank_register.bank\[2\]\[53\] _05382_ _07685_ vssd1 vssd1 vccd1 vccd1
+ _07689_ sky130_fd_sc_hd__mux2_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17306_ net536 _00749_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[84\]
+ sky130_fd_sc_hd__dfxtp_1
X_14518_ fifo_bank_register.bank\[9\]\[106\] _02793_ _02845_ _02846_ _02847_ vssd1
+ vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18286_ clknet_leaf_26_clk _01717_ net642 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[52\]
+ sky130_fd_sc_hd__dfrtp_4
X_15498_ _03652_ _04784_ _05245_ _03662_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17237_ net506 _00680_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_14449_ fifo_bank_register.bank\[5\]\[99\] _02714_ _02715_ fifo_bank_register.bank\[3\]\[99\]
+ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17168_ net546 _00611_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[74\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16119_ _04074_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17099_ net473 _00542_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_09990_ net173 ks1.key_reg\[23\] _05825_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__mux2_4
XFILLER_0_122_1112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08941_ _04916_ _04957_ _04959_ _04911_ _04964_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a221o_2
XFILLER_0_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_200_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_209_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _04883_ _04887_ _04892_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__or4_1
XFILLER_0_209_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_211_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_220_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09424_ _05377_ vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_165_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09355_ _05330_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_212_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08306_ net186 net185 net187 net188 vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__or4b_1
X_09286_ _05283_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08237_ net66 net65 net68 net67 vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__or4_4
XFILLER_0_90_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_219_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10130_ _04626_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_219_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10061_ _05888_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__clkbuf_1
XTAP_5724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13820_ _02136_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_214_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_203_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13751_ fifo_bank_register.bank\[0\]\[21\] _02165_ _02158_ vssd1 vssd1 vccd1 vccd1
+ _02166_ sky130_fd_sc_hd__mux2_1
X_10963_ mix1.data_o\[119\] _04626_ _05617_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_82_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12702_ fifo_bank_register.bank\[2\]\[17\] _05305_ _07640_ vssd1 vssd1 vccd1 vccd1
+ _07648_ sky130_fd_sc_hd__mux2_1
X_16470_ _04195_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__inv_2
XFILLER_0_168_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13682_ fifo_bank_register.bank\[9\]\[15\] _08190_ _02100_ _02101_ _02102_ vssd1
+ vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_214_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10894_ sub1.data_o\[113\] _06639_ _06478_ vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15421_ _03603_ _04949_ _05560_ _03614_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12633_ _07611_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15352_ net743 _03525_ _03560_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_182_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18140_ clknet_leaf_53_clk sbox1.next_alph\[2\] net657 vssd1 vssd1 vccd1 vccd1 sbox1.alph\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12564_ _07508_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_164_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14303_ fifo_bank_register.bank\[1\]\[82\] _02640_ _02641_ fifo_bank_register.bank\[8\]\[82\]
+ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_164_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11515_ fifo_bank_register.bank\[7\]\[97\] _05474_ _07013_ vssd1 vssd1 vccd1 vccd1
+ _07021_ sky130_fd_sc_hd__mux2_1
X_18071_ net554 _01514_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[73\]
+ sky130_fd_sc_hd__dfxtp_1
X_15283_ net773 _03529_ _03144_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12495_ fifo_bank_register.bank\[3\]\[47\] _05369_ _07531_ vssd1 vssd1 vccd1 vccd1
+ _07539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17022_ net571 _00465_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[56\]
+ sky130_fd_sc_hd__dfxtp_1
X_14234_ fifo_bank_register.bank\[7\]\[75\] _02542_ _02551_ fifo_bank_register.bank\[2\]\[75\]
+ _02594_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11446_ fifo_bank_register.bank\[7\]\[64\] _05405_ _06980_ vssd1 vssd1 vccd1 vccd1
+ _06985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14165_ _02532_ fifo_bank_register.data_out\[67\] _02533_ vssd1 vssd1 vccd1 vccd1
+ _02534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11377_ fifo_bank_register.bank\[7\]\[31\] _05336_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13116_ _07866_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__clkbuf_1
X_10328_ _06076_ _06125_ _06131_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__o21ai_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _02142_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__clkbuf_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_221_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ net523 _01367_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_13047_ _07830_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__clkbuf_1
X_10259_ _05913_ _05972_ sub1.data_o\[50\] _05902_ vssd1 vssd1 vccd1 vccd1 _06068_
+ sky130_fd_sc_hd__a31o_1
X_17855_ net491 _01298_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_227_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16806_ clknet_leaf_80_clk _00250_ net578 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[97\]
+ sky130_fd_sc_hd__dfrtp_4
X_17786_ net563 _01229_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_14998_ addroundkey_data_o\[114\] _03079_ _03271_ vssd1 vssd1 vccd1 vccd1 _03272_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16737_ clknet_leaf_52_clk _00181_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_1258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13949_ fifo_bank_register.bank\[0\]\[43\] _02341_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_163_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_73_clk clknet_3_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_202_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16668_ net453 _00116_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[108\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18407_ clknet_leaf_25_clk _01837_ net650 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[92\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_159_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_201_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15619_ _03736_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16599_ net415 _00047_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_174_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _05149_ _05150_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18338_ clknet_leaf_35_clk _01768_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09071_ _05016_ _05067_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18269_ clknet_leaf_34_clk _01700_ net662 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_163_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_163_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_204_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09973_ net43 mix1.data_o\[22\] _05699_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_217_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_204_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08924_ addroundkey_data_o\[13\] mix1.data_o\[13\] _04657_ vssd1 vssd1 vccd1 vccd1
+ _04948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_216_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08855_ _04661_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__buf_4
XFILLER_0_225_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08786_ _04706_ _04808_ _04809_ _04675_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a22o_1
XFILLER_0_212_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_170_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_174_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_64_clk clknet_3_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09407_ fifo_bank_register.bank\[9\]\[45\] _05365_ _05355_ vssd1 vssd1 vccd1 vccd1
+ _05366_ sky130_fd_sc_hd__mux2_1
XFILLER_0_211_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09338_ net173 vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09269_ net169 vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_161_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_181_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11300_ _06906_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__clkbuf_1
X_12280_ _05426_ fifo_bank_register.bank\[4\]\[74\] _07420_ vssd1 vssd1 vccd1 vccd1
+ _07425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11231_ _05462_ fifo_bank_register.bank\[8\]\[91\] _06869_ vssd1 vssd1 vccd1 vccd1
+ _06871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11162_ _06834_ vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10113_ _05608_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__buf_4
XFILLER_0_105_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11093_ _06798_ vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__clkbuf_1
X_15970_ _03941_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__clkbuf_1
XTAP_5521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14921_ _03124_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__xnor2_4
X_10044_ _05873_ vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__clkbuf_1
XTAP_5554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold50 mix1.data_reg\[71\] vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_215_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold61 mix1.data_reg\[79\] vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 mix1.data_reg\[60\] vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17640_ net418 _01083_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_5598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold83 mix1.data_reg\[50\] vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ addroundkey_data_o\[69\] _03108_ _03066_ addroundkey_data_o\[37\] vssd1 vssd1
+ vccd1 vccd1 _03128_ sky130_fd_sc_hd__a22o_1
Xhold94 mix1.data_reg\[52\] vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13803_ fifo_bank_register.bank\[5\]\[28\] _02141_ _02143_ fifo_bank_register.bank\[3\]\[28\]
+ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__a22o_1
X_14783_ _03058_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__buf_4
X_17571_ net400 _01014_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_11995_ _07274_ vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_55_clk clknet_3_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16522_ _04345_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__clkbuf_1
X_13734_ fifo_bank_register.bank\[6\]\[20\] _02147_ _02149_ fifo_bank_register.bank\[4\]\[20\]
+ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a22o_1
X_10946_ addroundkey_data_o\[117\] _06687_ _06612_ vssd1 vssd1 vccd1 vccd1 _06688_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_196_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13665_ fifo_bank_register.bank\[1\]\[13\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__a22o_1
X_16453_ _04130_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10877_ net143 ks1.key_reg\[111\] _06579_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _03019_ _03593_ _05228_ _03602_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12616_ _07602_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__clkbuf_1
X_16384_ _04146_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__inv_2
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ fifo_bank_register.bank\[6\]\[6\] _08105_ _08108_ fifo_bank_register.bank\[4\]\[6\]
+ vssd1 vssd1 vccd1 vccd1 _08161_ sky130_fd_sc_hd__a22o_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15335_ _03145_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18123_ net531 _01566_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[125\]
+ sky130_fd_sc_hd__dfxtp_1
X_12547_ _07566_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_227_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15266_ net785 _03516_ _03498_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__mux2_1
X_18054_ net574 _01497_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[56\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_124_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12478_ fifo_bank_register.bank\[3\]\[39\] _05352_ _07520_ vssd1 vssd1 vccd1 vccd1
+ _07530_ sky130_fd_sc_hd__mux2_1
XANTENNA_3 _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17005_ net414 _00448_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14217_ fifo_bank_register.bank\[5\]\[73\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[73\]
+ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11429_ fifo_bank_register.bank\[7\]\[56\] _05388_ _06969_ vssd1 vssd1 vccd1 vccd1
+ _06976_ sky130_fd_sc_hd__mux2_1
X_15197_ _03322_ _03443_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14148_ _02518_ fifo_bank_register.data_out\[65\] _02452_ vssd1 vssd1 vccd1 vccd1
+ _02519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14079_ fifo_bank_register.bank\[1\]\[58\] _02397_ _02398_ fifo_bank_register.bank\[8\]\[58\]
+ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a22o_1
XFILLER_0_225_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17907_ net406 _01350_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_225_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_207_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08640_ addroundkey_data_o\[20\] mix1.data_o\[20\] _04663_ vssd1 vssd1 vccd1 vccd1
+ _04664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_179_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17838_ net463 _01281_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[104\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_222_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_179_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08571_ _04604_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__buf_1
X_17769_ net428 _01212_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[35\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_228_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09123_ _05119_ _05131_ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__a21o_2
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_161_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09054_ _05015_ _05065_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_206_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_198_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09956_ net41 mix1.data_o\[20\] _05699_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08907_ _04884_ _04929_ _04930_ _04675_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _05731_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__xor2_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ ks1.key_reg\[14\] _04725_ _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_225_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _04721_ _04759_ _04761_ _04645_ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__o221a_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_clk clknet_3_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10800_ _06395_ _06514_ sub1.data_o\[103\] _05675_ vssd1 vssd1 vccd1 vccd1 _06556_
+ sky130_fd_sc_hd__a31o_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11780_ fifo_bank_register.bank\[6\]\[94\] _05468_ _07156_ vssd1 vssd1 vccd1 vccd1
+ _07161_ sky130_fd_sc_hd__mux2_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_178_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731_ _06491_ _06490_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13450_ _08042_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10662_ addroundkey_data_o\[89\] _06430_ _06431_ vssd1 vssd1 vccd1 vccd1 _06432_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12401_ _07489_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_192_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_180_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13381_ _08006_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__clkbuf_1
X_10593_ _06367_ _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__xnor2_1
X_15120_ _03179_ _03195_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_1_1272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12332_ _05478_ fifo_bank_register.bank\[4\]\[99\] _07442_ vssd1 vssd1 vccd1 vccd1
+ _07452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15051_ _03290_ _03323_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_107_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12263_ _05409_ fifo_bank_register.bank\[4\]\[66\] _07409_ vssd1 vssd1 vccd1 vccd1
+ _07416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_181_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14002_ _02136_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__clkbuf_4
X_11214_ _05445_ fifo_bank_register.bank\[8\]\[83\] _06858_ vssd1 vssd1 vccd1 vccd1
+ _06862_ sky130_fd_sc_hd__mux2_1
X_12194_ _05340_ fifo_bank_register.bank\[4\]\[33\] _07376_ vssd1 vssd1 vccd1 vccd1
+ _07380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_222_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11145_ _05375_ fifo_bank_register.bank\[8\]\[50\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06826_ sky130_fd_sc_hd__mux2_1
XTAP_6041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_6052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11076_ _05307_ fifo_bank_register.bank\[8\]\[18\] _06780_ vssd1 vssd1 vccd1 vccd1
+ _06789_ sky130_fd_sc_hd__mux2_1
X_15953_ ks1.col\[2\] _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__xor2_4
XTAP_6096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_223_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput140 key_i[109] vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_8
XTAP_5362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput151 key_i[119] vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_8
XTAP_5373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10027_ _05858_ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__clkbuf_1
X_14904_ _03175_ _03178_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__nor2_8
Xinput162 key_i[13] vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__buf_4
XFILLER_0_204_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput173 key_i[23] vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_4
Xinput184 key_i[33] vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_4
XTAP_5395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15884_ _04368_ _04716_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_208_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput195 key_i[43] vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_4
XTAP_4672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17623_ net497 _01066_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_215_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14835_ sub1.data_o\[117\] _03055_ _03110_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_clk clknet_3_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_176_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17554_ net543 _00997_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[76\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_187_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11978_ _07265_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__clkbuf_1
X_14766_ ks1.col\[19\] _05172_ _00007_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _04336_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__clkbuf_1
X_10929_ _05574_ _06670_ _06671_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13717_ fifo_bank_register.bank\[0\]\[19\] _02133_ _02068_ vssd1 vssd1 vccd1 vccd1
+ _02134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_188_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17485_ net479 _00928_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_14697_ fifo_bank_register.bank\[1\]\[127\] _08111_ _08114_ fifo_bank_register.bank\[8\]\[127\]
+ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16436_ _04298_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__clkbuf_1
X_13648_ fifo_bank_register.bank\[6\]\[11\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a22o_1
XFILLER_0_229_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_183_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13579_ fifo_bank_register.bank\[7\]\[4\] _08078_ _08093_ fifo_bank_register.bank\[2\]\[4\]
+ _08145_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__a221o_1
X_16367_ _04259_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_171_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_204_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18106_ net450 _01549_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[108\]
+ sky130_fd_sc_hd__dfxtp_1
X_15318_ _03551_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__clkbuf_1
X_16298_ _04223_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_164_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18037_ net415 _01480_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[39\]
+ sky130_fd_sc_hd__dfxtp_1
X_15249_ _03139_ _03379_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__xor2_4
XFILLER_0_169_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09810_ _05662_ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_226_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ round\[3\] _05568_ net258 _05581_ _05600_ vssd1 vssd1 vccd1 vccd1 _00152_
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_201_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_226_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09672_ addroundkey_round\[3\] _04637_ _04642_ _05544_ vssd1 vssd1 vccd1 vccd1 _00139_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_207_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08623_ _04371_ _04645_ _04646_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_19_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ addroundkey_data_o\[115\] fifo_bank_register.data_out\[115\] _04589_ vssd1
+ vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__mux2_4
XFILLER_0_210_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_171_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_212_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08485_ addroundkey_data_o\[82\] fifo_bank_register.data_out\[82\] _04556_ vssd1
+ vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_175_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_174_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_220_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09106_ sbox1.inversion_to_invert_var\[0\] _05105_ sbox1.inversion_to_invert_var\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__and3b_1
XFILLER_0_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ _05058_ vssd1 vssd1 vccd1 vccd1 sbox1.ah\[3\] sky130_fd_sc_hd__inv_2
XFILLER_0_14_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_217_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09939_ mix1.data_o\[18\] _05576_ _05758_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__o21a_1
X_12950_ fifo_bank_register.bank\[1\]\[6\] _05282_ _07772_ vssd1 vssd1 vccd1 vccd1
+ _07779_ sky130_fd_sc_hd__mux2_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11901_ _07225_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__clkbuf_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _07742_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__clkbuf_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 net155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11832_ fifo_bank_register.bank\[6\]\[119\] _05520_ _07178_ vssd1 vssd1 vccd1 vccd1
+ _07188_ sky130_fd_sc_hd__mux2_1
X_14620_ _02937_ fifo_bank_register.data_out\[117\] _02938_ vssd1 vssd1 vccd1 vccd1
+ _02939_ sky130_fd_sc_hd__mux2_1
XANTENNA_223 net220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_213_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 net244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _02142_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__clkbuf_4
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 _04748_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_278 addroundkey_data_o\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ fifo_bank_register.bank\[6\]\[86\] _05451_ _07145_ vssd1 vssd1 vccd1 vccd1
+ _07152_ sky130_fd_sc_hd__mux2_1
XFILLER_0_200_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_289 sub1.data_o\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ net124 mix1.data_o\[96\] _06476_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__mux2_1
X_13502_ fifo_bank_register.read_ptr\[0\] fifo_bank_register.read_ptr\[1\] _05262_
+ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ net397 _00713_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ fifo_bank_register.bank\[5\]\[102\] _02795_ _02796_ fifo_bank_register.bank\[3\]\[102\]
+ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__a22o_1
XFILLER_0_181_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11694_ fifo_bank_register.bank\[6\]\[53\] _05382_ _07112_ vssd1 vssd1 vccd1 vccd1
+ _07116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16221_ net214 ks1.key_reg\[60\] _03982_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__mux2_1
X_13433_ _08033_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__clkbuf_1
X_10645_ _05614_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16152_ _04102_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__xor2_1
XFILLER_0_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13364_ _07997_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__clkbuf_1
X_10576_ _06090_ _06342_ sub1.data_o\[82\] _06079_ vssd1 vssd1 vccd1 vccd1 _06353_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_107_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_228_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15103_ _03246_ _03373_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12315_ _07443_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__clkbuf_1
X_16083_ _04042_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__clkbuf_1
X_13295_ _07961_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15034_ _03297_ _03306_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__xnor2_2
X_12246_ _05392_ fifo_bank_register.bank\[4\]\[58\] _07398_ vssd1 vssd1 vccd1 vccd1
+ _07407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12177_ _05323_ fifo_bank_register.bank\[4\]\[25\] _07365_ vssd1 vssd1 vccd1 vccd1
+ _07371_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11128_ _05359_ fifo_bank_register.bank\[8\]\[42\] _06814_ vssd1 vssd1 vccd1 vccd1
+ _06817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_208_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16985_ net502 _00428_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_219_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_5170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11059_ _06768_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__buf_4
X_15936_ net183 ks1.key_reg\[32\] _03910_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__mux2_1
XTAP_5181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_218_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15867_ sub1.data_o\[88\] _05547_ _04888_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_189_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17606_ net475 _01049_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_176_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14818_ sub1.data_o\[13\] _04376_ _03081_ _03093_ vssd1 vssd1 vccd1 vccd1 _03094_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18586_ clknet_leaf_76_clk _02015_ net589 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[113\]
+ sky130_fd_sc_hd__dfrtp_1
X_15798_ mix1.data_o\[99\] net719 _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__mux2_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ net570 _00980_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14749_ _03038_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_191_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_171_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_157_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08270_ _04425_ _04426_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17468_ net456 _00911_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[118\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_229_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16419_ _04289_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17399_ net408 _00842_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[4\]\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_172_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_8_clk clknet_3_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_227_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_226_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09724_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09655_ _05533_ vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_210_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08606_ _04631_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.clk sky130_fd_sc_hd__clkbuf_2
XFILLER_0_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ net134 vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__buf_2
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_194_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ addroundkey_data_o\[107\] fifo_bank_register.data_out\[107\] _04578_ vssd1
+ vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__mux2_2
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08468_ addroundkey_data_o\[74\] fifo_bank_register.data_out\[74\] _04545_ vssd1
+ vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__mux2_2
XFILLER_0_65_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08399_ addroundkey_data_o\[41\] fifo_bank_register.data_out\[41\] _04512_ vssd1
+ vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__mux2_2
XFILLER_0_68_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ _06222_ vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_208_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10361_ sub1.data_o\[59\] _06159_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12100_ _07329_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13080_ _07847_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10292_ _06096_ _06098_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12031_ _07293_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_178_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_218_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout660 net670 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_219_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16770_ clknet_leaf_48_clk _00214_ net610 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[61\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13982_ _08068_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__buf_8
XFILLER_0_219_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_176_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15721_ _03790_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ fifo_bank_register.bank\[2\]\[127\] _05536_ _07628_ vssd1 vssd1 vccd1 vccd1
+ _07769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_213_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ clknet_leaf_35_clk _01870_ net665 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[125\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15652_ _03754_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_185_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ _07733_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__clkbuf_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_200_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _02923_ fifo_bank_register.data_out\[115\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18371_ clknet_leaf_37_clk _01801_ net667 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[56\]
+ sky130_fd_sc_hd__dfrtp_4
X_11815_ _07179_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__clkbuf_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_201_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_157_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15583_ _05103_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__clkbuf_4
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _07697_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__clkbuf_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_173_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_200_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17322_ net452 _00765_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[100\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11746_ fifo_bank_register.bank\[6\]\[78\] _05434_ _07134_ vssd1 vssd1 vccd1 vccd1
+ _07143_ sky130_fd_sc_hd__mux2_1
X_14534_ fifo_bank_register.bank\[1\]\[108\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[108\]
+ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_165_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17253_ net424 _00696_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ fifo_bank_register.bank\[6\]\[45\] _05365_ _07101_ vssd1 vssd1 vccd1 vccd1
+ _07107_ sky130_fd_sc_hd__mux2_1
X_14465_ fifo_bank_register.bank\[6\]\[100\] _02799_ _02800_ fifo_bank_register.bank\[4\]\[100\]
+ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_183_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16204_ _04111_ _04140_ _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10628_ _06381_ _06394_ _06400_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13416_ _08024_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_226_1329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17184_ net409 _00627_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[90\]
+ sky130_fd_sc_hd__dfxtp_1
X_14396_ fifo_bank_register.bank\[0\]\[92\] _02739_ _02725_ vssd1 vssd1 vccd1 vccd1
+ _02740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13347_ _07988_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__clkbuf_1
X_16135_ _04957_ _04088_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__or2_1
X_10559_ addroundkey_data_o\[80\] _06337_ _06327_ vssd1 vssd1 vccd1 vccd1 _06338_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_161_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13278_ _07952_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__clkbuf_1
X_16066_ net142 ks1.key_reg\[110\] _03979_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__mux2_2
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15017_ _03287_ _03288_ _03289_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_121_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12229_ _07364_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__buf_4
XFILLER_0_208_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_202_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_209_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16968_ net476 _00411_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15919_ _03717_ _04943_ _05219_ _03897_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a31o_1
X_16899_ net527 _00342_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[8\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_190_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09440_ net209 vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__buf_2
XFILLER_0_91_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09371_ _05341_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18569_ clknet_leaf_64_clk _01998_ net599 vssd1 vssd1 vccd1 vccd1 ks1.key_reg\[96\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_192_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ addroundkey_data_o\[5\] fifo_bank_register.data_out\[5\] _04468_ vssd1 vssd1
+ vccd1 vccd1 _04474_ sky130_fd_sc_hd__mux2_2
XFILLER_0_191_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08253_ net97 net96 net99 net98 vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__or4_2
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_162_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput263 net263 vssd1 vssd1 vccd1 vccd1 data_o[102] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput274 net274 vssd1 vssd1 vccd1 vccd1 data_o[112] sky130_fd_sc_hd__buf_2
XFILLER_0_199_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput285 net285 vssd1 vssd1 vccd1 vccd1 data_o[122] sky130_fd_sc_hd__clkbuf_4
XTAP_5906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput296 net296 vssd1 vssd1 vccd1 vccd1 data_o[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_227_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_226_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_199_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_227_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09707_ _05570_ vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09638_ net153 vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_179_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_210_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_168_947 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09569_ _05475_ vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11600_ fifo_bank_register.bank\[6\]\[9\] _05288_ _07056_ vssd1 vssd1 vccd1 vccd1
+ _07066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_194_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ _07583_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11531_ _07029_ vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14250_ fifo_bank_register.bank\[7\]\[77\] _02542_ _02551_ fifo_bank_register.bank\[2\]\[77\]
+ _02608_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__a221o_1
XFILLER_0_190_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11462_ _06993_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_184_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_208_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13201_ _07910_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__clkbuf_1
X_10413_ _06207_ vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14181_ fifo_bank_register.bank\[0\]\[69\] _02547_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_180_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11393_ fifo_bank_register.bank\[7\]\[39\] _05352_ _06947_ vssd1 vssd1 vccd1 vccd1
+ _06957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13132_ fifo_bank_register.bank\[1\]\[92\] _05464_ _07872_ vssd1 vssd1 vccd1 vccd1
+ _07875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10344_ mix1.data_o\[57\] _06138_ _05993_ _05994_ sub1.data_o\[57\] vssd1 vssd1 vccd1
+ vccd1 _06146_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17940_ net525 _01383_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[78\]
+ sky130_fd_sc_hd__dfxtp_1
X_13063_ _07838_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__clkbuf_1
X_10275_ sub1.data_o\[51\] _05971_ _06081_ _06082_ _05941_ vssd1 vssd1 vccd1 vccd1
+ _06083_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12014_ _07284_ vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__clkbuf_1
X_17871_ net426 _01314_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[9\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_178_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16822_ clknet_leaf_75_clk _00266_ net587 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[113\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_206_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_219_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout490 net498 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__buf_2
XFILLER_0_191_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16753_ clknet_leaf_65_clk _00197_ net603 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[44\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_219_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13965_ fifo_bank_register.bank\[0\]\[45\] _02355_ _02320_ vssd1 vssd1 vccd1 vccd1
+ _02356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15704_ _03781_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_191_1369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12916_ _07760_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__clkbuf_1
X_16684_ net495 _00132_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13896_ fifo_bank_register.bank\[6\]\[38\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[38\]
+ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_213_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18423_ clknet_leaf_83_clk _01853_ net582 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[108\]
+ sky130_fd_sc_hd__dfrtp_2
X_15635_ _03745_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_186_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12847_ _07724_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__clkbuf_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18354_ clknet_leaf_15_clk _01784_ net629 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15566_ sub1.data_o\[103\] sub1.data_o\[39\] _03574_ vssd1 vssd1 vccd1 vccd1 _03707_
+ sky130_fd_sc_hd__mux2_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _07688_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__clkbuf_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ net539 _00748_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[83\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_189_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14517_ fifo_bank_register.bank\[1\]\[106\] _02802_ _02803_ fifo_bank_register.bank\[8\]\[106\]
+ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__a22o_1
X_18285_ clknet_leaf_26_clk _01716_ net649 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[51\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_56_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11729_ _07078_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__buf_4
X_15497_ sub1.data_o\[111\] _03660_ _03653_ sub1.data_o\[47\] vssd1 vssd1 vccd1 vccd1
+ _03662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_182_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ net506 _00679_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[5\]\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14448_ _08181_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ net554 _00610_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[73\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14379_ _02157_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16118_ ks1.key_reg\[19\] _04073_ _03958_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17098_ net474 _00541_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08940_ _04721_ _04961_ _04963_ _04750_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__a2bb2o_1
X_16049_ _05218_ _04011_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_209_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08871_ _04684_ _04893_ _04894_ _04689_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_208_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_223_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_224_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_211_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_189_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09423_ fifo_bank_register.bank\[9\]\[50\] _05375_ _05376_ vssd1 vssd1 vccd1 vccd1
+ _05377_ sky130_fd_sc_hd__mux2_1
XFILLER_0_176_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09354_ fifo_bank_register.bank\[9\]\[28\] _05329_ _05313_ vssd1 vssd1 vccd1 vccd1
+ _05330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08305_ net182 net184 net183 net181 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_117_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09285_ fifo_bank_register.bank\[9\]\[6\] _05282_ _05270_ vssd1 vssd1 vccd1 vccd1
+ _05283_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08236_ _04380_ _04382_ _04387_ _04392_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__or4_4
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_160_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_166_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_160_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_219_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_5703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ addroundkey_data_o\[31\] _05887_ _05872_ vssd1 vssd1 vccd1 vccd1 _05888_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_5714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_5725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_227_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_214_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_216_1317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_214_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10962_ _05574_ _06700_ _06701_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__a21o_1
X_13750_ fifo_bank_register.bank\[9\]\[21\] _02137_ _02162_ _02163_ _02164_ vssd1
+ vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ _07647_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10893_ net16 mix1.data_o\[113\] _06476_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13681_ fifo_bank_register.bank\[1\]\[15\] _08199_ _08200_ fifo_bank_register.bank\[8\]\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_214_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_195_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15420_ sub1.data_o\[18\] _03606_ _03613_ _03611_ vssd1 vssd1 vccd1 vccd1 _03614_
+ sky130_fd_sc_hd__a22o_1
X_12632_ fifo_bank_register.bank\[3\]\[112\] _05506_ _07608_ vssd1 vssd1 vccd1 vccd1
+ _07611_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15351_ _03568_ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__clkbuf_1
X_12563_ _07574_ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_164_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_202_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11514_ _07020_ vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__clkbuf_1
X_14302_ fifo_bank_register.bank\[6\]\[82\] _02637_ _02638_ fifo_bank_register.bank\[4\]\[82\]
+ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18070_ net557 _01513_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[72\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15282_ _03464_ _03479_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_151_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12494_ _07538_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_202_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17021_ net570 _00464_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_184_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _06984_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14233_ fifo_bank_register.bank\[5\]\[75\] _02552_ _02553_ fifo_bank_register.bank\[3\]\[75\]
+ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14164_ _08068_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11376_ _06948_ vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_221_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10327_ sub1.data_o\[55\] _05971_ _06128_ _06130_ _06118_ vssd1 vssd1 vccd1 vccd1
+ _06131_ sky130_fd_sc_hd__a221o_1
X_13115_ fifo_bank_register.bank\[1\]\[84\] _05447_ _07861_ vssd1 vssd1 vccd1 vccd1
+ _07866_ sky130_fd_sc_hd__mux2_1
X_14095_ _02140_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_221_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_219_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ net527 _01366_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_13046_ fifo_bank_register.bank\[1\]\[51\] _05378_ _07828_ vssd1 vssd1 vccd1 vccd1
+ _07830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_221_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10258_ sub1.data_o\[50\] _06066_ _05936_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__mux2_1
X_17854_ net471 _01297_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[120\]
+ sky130_fd_sc_hd__dfxtp_1
X_10189_ _06001_ _06003_ _06004_ _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_206_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_205_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16805_ clknet_leaf_80_clk _00249_ net578 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[96\]
+ sky130_fd_sc_hd__dfrtp_4
X_17785_ net573 _01228_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_227_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_191_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14997_ addroundkey_data_o\[18\] _03208_ _03086_ _03270_ vssd1 vssd1 vccd1 vccd1
+ _03271_ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_221_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16736_ clknet_leaf_43_clk _00180_ net655 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[27\]
+ sky130_fd_sc_hd__dfrtp_2
X_13948_ fifo_bank_register.bank\[9\]\[43\] _02307_ _02338_ _02339_ _02340_ vssd1
+ vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_191_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_186_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_158_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16667_ net451 _00115_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_186_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13879_ fifo_bank_register.bank\[6\]\[36\] _02232_ _02233_ fifo_bank_register.bank\[4\]\[36\]
+ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a22o_1
XFILLER_0_201_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18406_ clknet_leaf_25_clk _01836_ net648 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[91\]
+ sky130_fd_sc_hd__dfrtp_4
X_15618_ mix1.data_o\[14\] _03477_ _03730_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_186_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16598_ net428 _00046_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[9\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18337_ clknet_leaf_35_clk _01767_ net664 vssd1 vssd1 vccd1 vccd1 mix1.data_o\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15549_ _03668_ _04935_ _05554_ _03695_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09070_ _05082_ _05083_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__nor2_1
X_18268_ clknet_leaf_33_clk _01699_ net663 vssd1 vssd1 vccd1 vccd1 sub1.data_o\[34\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17219_ net496 _00662_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[6\]\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18199_ clknet_leaf_10_clk _01630_ net623 vssd1 vssd1 vccd1 vccd1 mix1.data_reg\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_163_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_198_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_229_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09972_ _05809_ vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_200_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08923_ addroundkey_data_o\[109\] mix1.data_o\[109\] _04702_ vssd1 vssd1 vccd1 vccd1
+ _04947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_209_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_225_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08854_ addroundkey_data_o\[120\] mix1.data_o\[120\] _04658_ vssd1 vssd1 vccd1 vccd1
+ _04878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_225_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_196_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ addroundkey_data_o\[27\] mix1.data_o\[27\] _04805_ vssd1 vssd1 vccd1 vccd1
+ _04809_ sky130_fd_sc_hd__mux2_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_224_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_170_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_211_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_196_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_211_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_177_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_220_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09406_ net197 vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_177_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_211_1269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09337_ _05318_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_192_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_164_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09268_ _05271_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_209_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08219_ _04376_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09199_ sbox1.alph\[2\] _05127_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_205_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_181_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11230_ _06870_ vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11161_ _05392_ fifo_bank_register.bank\[8\]\[58\] _06825_ vssd1 vssd1 vccd1 vccd1
+ _06834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_222_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_219_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10112_ net58 mix1.data_o\[36\] _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__mux2_1
XTAP_5500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_179_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11092_ _05323_ fifo_bank_register.bank\[8\]\[25\] _06792_ vssd1 vssd1 vccd1 vccd1
+ _06798_ sky130_fd_sc_hd__mux2_1
XTAP_5511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_228_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_5533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10043_ addroundkey_data_o\[29\] _05871_ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_
+ sky130_fd_sc_hd__mux2_1
X_14920_ _03191_ _03194_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__nor2_8
XTAP_5544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold40 mix1.data_reg\[54\] vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold51 ks1.key_reg\[105\] vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold62 mix1.data_reg\[42\] vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_5588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold73 mix1.data_reg\[59\] vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14851_ sub1.data_o\[101\] _03055_ _03126_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__a21oi_4
XTAP_5599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold84 mix1.data_reg\[41\] vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_4876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold95 mix1.data_reg\[126\] vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _02210_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_215_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17570_ net403 _01013_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_216_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14782_ _04658_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__buf_4
X_11994_ fifo_bank_register.bank\[5\]\[67\] _05411_ _07266_ vssd1 vssd1 vccd1 vccd1
+ _07274_ sky130_fd_sc_hd__mux2_1
X_16521_ net776 _03505_ _04343_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__mux2_1
X_13733_ _02148_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__clkbuf_4
X_10945_ _06685_ _06686_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_196_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ _04215_ _04117_ _04306_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__o21ai_1
X_13664_ fifo_bank_register.bank\[6\]\[13\] _08196_ _08197_ fifo_bank_register.bank\[4\]\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__a22o_1
X_10876_ _06583_ _06622_ _06623_ _06587_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_183_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15403_ sub1.data_o\[77\] _03600_ _03595_ sub1.data_o\[13\] vssd1 vssd1 vccd1 vccd1
+ _03602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_220_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12615_ fifo_bank_register.bank\[3\]\[104\] _05489_ _07597_ vssd1 vssd1 vccd1 vccd1
+ _07602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_183_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16383_ _04268_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__clkbuf_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13595_ fifo_bank_register.bank\[7\]\[6\] _08078_ _08093_ fifo_bank_register.bank\[2\]\[6\]
+ _08159_ vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__a221o_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18122_ net531 _01565_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _03559_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_164_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12546_ fifo_bank_register.bank\[3\]\[71\] _05420_ _07564_ vssd1 vssd1 vccd1 vccd1
+ _07566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18053_ net574 _01496_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15265_ _03423_ _03438_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__xnor2_4
X_12477_ _07529_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__clkbuf_1
X_17004_ net418 _00447_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[7\]\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_4 _02151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_227_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14216_ _02579_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__clkbuf_1
X_11428_ _06975_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__clkbuf_1
X_15196_ _03394_ _03458_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_158_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11359_ _06939_ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__clkbuf_1
X_14147_ fifo_bank_register.bank\[0\]\[65\] _02517_ _02482_ vssd1 vssd1 vccd1 vccd1
+ _02518_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14078_ fifo_bank_register.bank\[6\]\[58\] _02394_ _02395_ fifo_bank_register.bank\[4\]\[58\]
+ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_225_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_158_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_184_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13029_ fifo_bank_register.bank\[1\]\[43\] _05361_ _07817_ vssd1 vssd1 vccd1 vccd1
+ _07821_ sky130_fd_sc_hd__mux2_1
X_17906_ net389 _01349_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[0\]\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_207_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17837_ net458 _01280_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_206_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08570_ addroundkey_data_o\[123\] fifo_bank_register.data_out\[123\] _04467_ vssd1
+ vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_178_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17768_ net430 _01211_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[1\]\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16719_ clknet_leaf_51_clk _00163_ net654 vssd1 vssd1 vccd1 vccd1 addroundkey_data_o\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17699_ net400 _01142_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[93\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09122_ sbox1.inversion_to_invert_var\[3\] _05114_ _05117_ _05129_ _05132_ vssd1
+ vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__o221a_1
XFILLER_0_161_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_228_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_162_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_199_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _05070_ vssd1 vssd1 vccd1 vccd1 sbox1.next_alph\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_170_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_198_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_204_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09955_ _05794_ vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_217_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_218_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08906_ addroundkey_data_o\[29\] mix1.data_o\[29\] _04702_ vssd1 vssd1 vccd1 vccd1
+ _04930_ sky130_fd_sc_hd__mux2_1
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ net162 ks1.key_reg\[13\] _05708_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__mux2_2
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ ks1.key_reg\[14\] _04729_ _04731_ net163 vssd1 vssd1 vccd1 vccd1 _04861_
+ sky130_fd_sc_hd__o31a_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_197_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _04763_ _04791_ _04648_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__o21ai_2
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_212_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08699_ addroundkey_start_i _04641_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_178_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10730_ _06395_ _06342_ sub1.data_o\[97\] _06384_ vssd1 vssd1 vccd1 vccd1 _06492_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_177_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_165_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10661_ _05792_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__buf_4
XFILLER_0_211_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_193_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12400_ fifo_bank_register.bank\[3\]\[2\] _05274_ _07486_ vssd1 vssd1 vccd1 vccd1
+ _07489_ sky130_fd_sc_hd__mux2_1
X_13380_ _05441_ fifo_bank_register.bank\[0\]\[81\] _08004_ vssd1 vssd1 vccd1 vccd1
+ _08006_ sky130_fd_sc_hd__mux2_1
X_10592_ net239 ks1.key_reg\[83\] _06097_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__mux2_4
XFILLER_0_90_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_180_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12331_ _07451_ vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15050_ _03307_ _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__xnor2_2
X_12262_ _07415_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_1285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14001_ _02387_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__clkbuf_1
X_11213_ _06861_ vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_1273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12193_ _07379_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_222_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11144_ _06791_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__buf_4
XTAP_6020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_207_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_6064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11075_ _06788_ vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__clkbuf_1
X_15952_ net255 ks1.key_reg\[98\] _03902_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__mux2_2
XTAP_6075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput130 key_i[0] vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
Xinput141 key_i[10] vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_4
XTAP_6097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_5363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput152 key_i[11] vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_4
X_10026_ addroundkey_data_o\[27\] _05857_ _05793_ vssd1 vssd1 vccd1 vccd1 _05858_
+ sky130_fd_sc_hd__mux2_1
X_14903_ addroundkey_data_o\[126\] _03078_ _03177_ vssd1 vssd1 vccd1 vccd1 _03178_
+ sky130_fd_sc_hd__a21oi_2
XTAP_5374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_170_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput163 key_i[14] vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_222_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15883_ _05547_ sub1.data_o\[64\] _05200_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__mux2_1
XTAP_4640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput174 key_i[24] vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_8
XTAP_4651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_215_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_5396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput185 key_i[34] vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_4
XTAP_4662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput196 key_i[44] vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_4
X_17622_ net496 _01065_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[2\]\[16\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_192_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14834_ sub1.data_o\[21\] _03100_ _03058_ _03109_ vssd1 vssd1 vccd1 vccd1 _03110_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_204_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ net543 _00996_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[75\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _03046_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__clkbuf_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11977_ fifo_bank_register.bank\[5\]\[59\] _05394_ _07255_ vssd1 vssd1 vccd1 vccd1
+ _07265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16504_ net787 _03467_ _04332_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__mux2_1
X_13716_ fifo_bank_register.bank\[9\]\[19\] _08190_ _02130_ _02131_ _02132_ vssd1
+ vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a2111o_1
X_10928_ _06630_ _06514_ sub1.data_o\[116\] _05675_ vssd1 vssd1 vccd1 vccd1 _06671_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_156_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17484_ net479 _00927_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.bank\[3\]\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_224_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14696_ fifo_bank_register.bank\[6\]\[127\] _08104_ _08107_ fifo_bank_register.bank\[4\]\[127\]
+ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_168_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16435_ ks1.key_reg\[112\] _04044_ _04295_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__mux2_1
X_13647_ fifo_bank_register.bank\[7\]\[11\] _08182_ _08191_ fifo_bank_register.bank\[2\]\[11\]
+ _02071_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__a221o_1
X_10859_ _06583_ _06607_ _06608_ _06587_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_229_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ net843 _04062_ _04252_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
X_13578_ fifo_bank_register.bank\[5\]\[4\] _08097_ _08100_ fifo_bank_register.bank\[3\]\[4\]
+ vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18105_ net451 _01548_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[107\]
+ sky130_fd_sc_hd__dfxtp_1
X_15317_ net732 _03435_ _03549_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12529_ fifo_bank_register.bank\[3\]\[63\] _05403_ _07553_ vssd1 vssd1 vccd1 vccd1
+ _07557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16297_ net834 _04056_ _04222_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_164_1341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18036_ net407 _01479_ vssd1 vssd1 vccd1 vccd1 fifo_bank_register.data_out\[38\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_112_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15248_ _03503_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_160_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15179_ _03297_ _03443_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_201_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09740_ _05595_ _05597_ _05599_ _05568_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__o211a_1
XFILLER_0_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
.ends

