magic
tech sky130A
magscale 1 2
timestamp 1698718705
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 14 2128 99254 97424
<< metal2 >>
rect 18 99200 74 100000
rect 1950 99200 2006 100000
rect 3882 99200 3938 100000
rect 6458 99200 6514 100000
rect 8390 99200 8446 100000
rect 10322 99200 10378 100000
rect 12254 99200 12310 100000
rect 14186 99200 14242 100000
rect 16762 99200 16818 100000
rect 18694 99200 18750 100000
rect 20626 99200 20682 100000
rect 22558 99200 22614 100000
rect 24490 99200 24546 100000
rect 27066 99200 27122 100000
rect 28998 99200 29054 100000
rect 30930 99200 30986 100000
rect 32862 99200 32918 100000
rect 34794 99200 34850 100000
rect 37370 99200 37426 100000
rect 39302 99200 39358 100000
rect 41234 99200 41290 100000
rect 43166 99200 43222 100000
rect 45742 99200 45798 100000
rect 47674 99200 47730 100000
rect 49606 99200 49662 100000
rect 51538 99200 51594 100000
rect 53470 99200 53526 100000
rect 56046 99200 56102 100000
rect 57978 99200 58034 100000
rect 59910 99200 59966 100000
rect 61842 99200 61898 100000
rect 63774 99200 63830 100000
rect 66350 99200 66406 100000
rect 68282 99200 68338 100000
rect 70214 99200 70270 100000
rect 72146 99200 72202 100000
rect 74078 99200 74134 100000
rect 76654 99200 76710 100000
rect 78586 99200 78642 100000
rect 80518 99200 80574 100000
rect 82450 99200 82506 100000
rect 84382 99200 84438 100000
rect 86958 99200 87014 100000
rect 88890 99200 88946 100000
rect 90822 99200 90878 100000
rect 92754 99200 92810 100000
rect 94686 99200 94742 100000
rect 97262 99200 97318 100000
rect 99194 99200 99250 100000
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 5814 0 5870 800
rect 7746 0 7802 800
rect 10322 0 10378 800
rect 12254 0 12310 800
rect 14186 0 14242 800
rect 16118 0 16174 800
rect 18050 0 18106 800
rect 20626 0 20682 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 28354 0 28410 800
rect 30930 0 30986 800
rect 32862 0 32918 800
rect 34794 0 34850 800
rect 36726 0 36782 800
rect 38658 0 38714 800
rect 41234 0 41290 800
rect 43166 0 43222 800
rect 45098 0 45154 800
rect 47030 0 47086 800
rect 48962 0 49018 800
rect 51538 0 51594 800
rect 53470 0 53526 800
rect 55402 0 55458 800
rect 57334 0 57390 800
rect 59266 0 59322 800
rect 61842 0 61898 800
rect 63774 0 63830 800
rect 65706 0 65762 800
rect 67638 0 67694 800
rect 70214 0 70270 800
rect 72146 0 72202 800
rect 74078 0 74134 800
rect 76010 0 76066 800
rect 77942 0 77998 800
rect 80518 0 80574 800
rect 82450 0 82506 800
rect 84382 0 84438 800
rect 86314 0 86370 800
rect 88246 0 88302 800
rect 90822 0 90878 800
rect 92754 0 92810 800
rect 94686 0 94742 800
rect 96618 0 96674 800
rect 98550 0 98606 800
<< obsm2 >>
rect 130 99144 1894 99362
rect 2062 99144 3826 99362
rect 3994 99144 6402 99362
rect 6570 99144 8334 99362
rect 8502 99144 10266 99362
rect 10434 99144 12198 99362
rect 12366 99144 14130 99362
rect 14298 99144 16706 99362
rect 16874 99144 18638 99362
rect 18806 99144 20570 99362
rect 20738 99144 22502 99362
rect 22670 99144 24434 99362
rect 24602 99144 27010 99362
rect 27178 99144 28942 99362
rect 29110 99144 30874 99362
rect 31042 99144 32806 99362
rect 32974 99144 34738 99362
rect 34906 99144 37314 99362
rect 37482 99144 39246 99362
rect 39414 99144 41178 99362
rect 41346 99144 43110 99362
rect 43278 99144 45686 99362
rect 45854 99144 47618 99362
rect 47786 99144 49550 99362
rect 49718 99144 51482 99362
rect 51650 99144 53414 99362
rect 53582 99144 55990 99362
rect 56158 99144 57922 99362
rect 58090 99144 59854 99362
rect 60022 99144 61786 99362
rect 61954 99144 63718 99362
rect 63886 99144 66294 99362
rect 66462 99144 68226 99362
rect 68394 99144 70158 99362
rect 70326 99144 72090 99362
rect 72258 99144 74022 99362
rect 74190 99144 76598 99362
rect 76766 99144 78530 99362
rect 78698 99144 80462 99362
rect 80630 99144 82394 99362
rect 82562 99144 84326 99362
rect 84494 99144 86902 99362
rect 87070 99144 88834 99362
rect 89002 99144 90766 99362
rect 90934 99144 92698 99362
rect 92866 99144 94630 99362
rect 94798 99144 97206 99362
rect 97374 99144 99138 99362
rect 20 856 99248 99144
rect 130 711 1894 856
rect 2062 711 3826 856
rect 3994 711 5758 856
rect 5926 711 7690 856
rect 7858 711 10266 856
rect 10434 711 12198 856
rect 12366 711 14130 856
rect 14298 711 16062 856
rect 16230 711 17994 856
rect 18162 711 20570 856
rect 20738 711 22502 856
rect 22670 711 24434 856
rect 24602 711 26366 856
rect 26534 711 28298 856
rect 28466 711 30874 856
rect 31042 711 32806 856
rect 32974 711 34738 856
rect 34906 711 36670 856
rect 36838 711 38602 856
rect 38770 711 41178 856
rect 41346 711 43110 856
rect 43278 711 45042 856
rect 45210 711 46974 856
rect 47142 711 48906 856
rect 49074 711 51482 856
rect 51650 711 53414 856
rect 53582 711 55346 856
rect 55514 711 57278 856
rect 57446 711 59210 856
rect 59378 711 61786 856
rect 61954 711 63718 856
rect 63886 711 65650 856
rect 65818 711 67582 856
rect 67750 711 70158 856
rect 70326 711 72090 856
rect 72258 711 74022 856
rect 74190 711 75954 856
rect 76122 711 77886 856
rect 78054 711 80462 856
rect 80630 711 82394 856
rect 82562 711 84326 856
rect 84494 711 86258 856
rect 86426 711 88190 856
rect 88358 711 90766 856
rect 90934 711 92698 856
rect 92866 711 94630 856
rect 94798 711 96562 856
rect 96730 711 98494 856
rect 98662 711 99248 856
<< metal3 >>
rect 99200 98608 100000 98728
rect 0 97928 800 98048
rect 99200 96568 100000 96688
rect 0 95888 800 96008
rect 99200 93848 100000 93968
rect 0 93168 800 93288
rect 99200 91808 100000 91928
rect 0 91128 800 91248
rect 99200 89768 100000 89888
rect 0 89088 800 89208
rect 99200 87728 100000 87848
rect 0 87048 800 87168
rect 99200 85688 100000 85808
rect 0 85008 800 85128
rect 99200 82968 100000 83088
rect 0 82288 800 82408
rect 99200 80928 100000 81048
rect 0 80248 800 80368
rect 99200 78888 100000 79008
rect 0 78208 800 78328
rect 99200 76848 100000 76968
rect 0 76168 800 76288
rect 99200 74808 100000 74928
rect 0 74128 800 74248
rect 99200 72088 100000 72208
rect 0 71408 800 71528
rect 99200 70048 100000 70168
rect 0 69368 800 69488
rect 99200 68008 100000 68128
rect 0 67328 800 67448
rect 99200 65968 100000 66088
rect 0 65288 800 65408
rect 99200 63928 100000 64048
rect 0 62568 800 62688
rect 99200 61208 100000 61328
rect 0 60528 800 60648
rect 99200 59168 100000 59288
rect 0 58488 800 58608
rect 99200 57128 100000 57248
rect 0 56448 800 56568
rect 99200 55088 100000 55208
rect 0 54408 800 54528
rect 99200 53048 100000 53168
rect 0 51688 800 51808
rect 99200 50328 100000 50448
rect 0 49648 800 49768
rect 99200 48288 100000 48408
rect 0 47608 800 47728
rect 99200 46248 100000 46368
rect 0 45568 800 45688
rect 99200 44208 100000 44328
rect 0 43528 800 43648
rect 99200 42168 100000 42288
rect 0 40808 800 40928
rect 99200 39448 100000 39568
rect 0 38768 800 38888
rect 99200 37408 100000 37528
rect 0 36728 800 36848
rect 99200 35368 100000 35488
rect 0 34688 800 34808
rect 99200 33328 100000 33448
rect 0 32648 800 32768
rect 99200 31288 100000 31408
rect 0 29928 800 30048
rect 99200 28568 100000 28688
rect 0 27888 800 28008
rect 99200 26528 100000 26648
rect 0 25848 800 25968
rect 99200 24488 100000 24608
rect 0 23808 800 23928
rect 99200 22448 100000 22568
rect 0 21768 800 21888
rect 99200 19728 100000 19848
rect 0 19048 800 19168
rect 99200 17688 100000 17808
rect 0 17008 800 17128
rect 99200 15648 100000 15768
rect 0 14968 800 15088
rect 99200 13608 100000 13728
rect 0 12928 800 13048
rect 99200 11568 100000 11688
rect 0 10888 800 11008
rect 99200 8848 100000 8968
rect 0 8168 800 8288
rect 99200 6808 100000 6928
rect 0 6128 800 6248
rect 99200 4768 100000 4888
rect 0 4088 800 4208
rect 99200 2728 100000 2848
rect 0 2048 800 2168
rect 99200 688 100000 808
<< obsm3 >>
rect 798 98528 99120 98701
rect 798 98128 99200 98528
rect 880 97848 99200 98128
rect 798 96768 99200 97848
rect 798 96488 99120 96768
rect 798 96088 99200 96488
rect 880 95808 99200 96088
rect 798 94048 99200 95808
rect 798 93768 99120 94048
rect 798 93368 99200 93768
rect 880 93088 99200 93368
rect 798 92008 99200 93088
rect 798 91728 99120 92008
rect 798 91328 99200 91728
rect 880 91048 99200 91328
rect 798 89968 99200 91048
rect 798 89688 99120 89968
rect 798 89288 99200 89688
rect 880 89008 99200 89288
rect 798 87928 99200 89008
rect 798 87648 99120 87928
rect 798 87248 99200 87648
rect 880 86968 99200 87248
rect 798 85888 99200 86968
rect 798 85608 99120 85888
rect 798 85208 99200 85608
rect 880 84928 99200 85208
rect 798 83168 99200 84928
rect 798 82888 99120 83168
rect 798 82488 99200 82888
rect 880 82208 99200 82488
rect 798 81128 99200 82208
rect 798 80848 99120 81128
rect 798 80448 99200 80848
rect 880 80168 99200 80448
rect 798 79088 99200 80168
rect 798 78808 99120 79088
rect 798 78408 99200 78808
rect 880 78128 99200 78408
rect 798 77048 99200 78128
rect 798 76768 99120 77048
rect 798 76368 99200 76768
rect 880 76088 99200 76368
rect 798 75008 99200 76088
rect 798 74728 99120 75008
rect 798 74328 99200 74728
rect 880 74048 99200 74328
rect 798 72288 99200 74048
rect 798 72008 99120 72288
rect 798 71608 99200 72008
rect 880 71328 99200 71608
rect 798 70248 99200 71328
rect 798 69968 99120 70248
rect 798 69568 99200 69968
rect 880 69288 99200 69568
rect 798 68208 99200 69288
rect 798 67928 99120 68208
rect 798 67528 99200 67928
rect 880 67248 99200 67528
rect 798 66168 99200 67248
rect 798 65888 99120 66168
rect 798 65488 99200 65888
rect 880 65208 99200 65488
rect 798 64128 99200 65208
rect 798 63848 99120 64128
rect 798 62768 99200 63848
rect 880 62488 99200 62768
rect 798 61408 99200 62488
rect 798 61128 99120 61408
rect 798 60728 99200 61128
rect 880 60448 99200 60728
rect 798 59368 99200 60448
rect 798 59088 99120 59368
rect 798 58688 99200 59088
rect 880 58408 99200 58688
rect 798 57328 99200 58408
rect 798 57048 99120 57328
rect 798 56648 99200 57048
rect 880 56368 99200 56648
rect 798 55288 99200 56368
rect 798 55008 99120 55288
rect 798 54608 99200 55008
rect 880 54328 99200 54608
rect 798 53248 99200 54328
rect 798 52968 99120 53248
rect 798 51888 99200 52968
rect 880 51608 99200 51888
rect 798 50528 99200 51608
rect 798 50248 99120 50528
rect 798 49848 99200 50248
rect 880 49568 99200 49848
rect 798 48488 99200 49568
rect 798 48208 99120 48488
rect 798 47808 99200 48208
rect 880 47528 99200 47808
rect 798 46448 99200 47528
rect 798 46168 99120 46448
rect 798 45768 99200 46168
rect 880 45488 99200 45768
rect 798 44408 99200 45488
rect 798 44128 99120 44408
rect 798 43728 99200 44128
rect 880 43448 99200 43728
rect 798 42368 99200 43448
rect 798 42088 99120 42368
rect 798 41008 99200 42088
rect 880 40728 99200 41008
rect 798 39648 99200 40728
rect 798 39368 99120 39648
rect 798 38968 99200 39368
rect 880 38688 99200 38968
rect 798 37608 99200 38688
rect 798 37328 99120 37608
rect 798 36928 99200 37328
rect 880 36648 99200 36928
rect 798 35568 99200 36648
rect 798 35288 99120 35568
rect 798 34888 99200 35288
rect 880 34608 99200 34888
rect 798 33528 99200 34608
rect 798 33248 99120 33528
rect 798 32848 99200 33248
rect 880 32568 99200 32848
rect 798 31488 99200 32568
rect 798 31208 99120 31488
rect 798 30128 99200 31208
rect 880 29848 99200 30128
rect 798 28768 99200 29848
rect 798 28488 99120 28768
rect 798 28088 99200 28488
rect 880 27808 99200 28088
rect 798 26728 99200 27808
rect 798 26448 99120 26728
rect 798 26048 99200 26448
rect 880 25768 99200 26048
rect 798 24688 99200 25768
rect 798 24408 99120 24688
rect 798 24008 99200 24408
rect 880 23728 99200 24008
rect 798 22648 99200 23728
rect 798 22368 99120 22648
rect 798 21968 99200 22368
rect 880 21688 99200 21968
rect 798 19928 99200 21688
rect 798 19648 99120 19928
rect 798 19248 99200 19648
rect 880 18968 99200 19248
rect 798 17888 99200 18968
rect 798 17608 99120 17888
rect 798 17208 99200 17608
rect 880 16928 99200 17208
rect 798 15848 99200 16928
rect 798 15568 99120 15848
rect 798 15168 99200 15568
rect 880 14888 99200 15168
rect 798 13808 99200 14888
rect 798 13528 99120 13808
rect 798 13128 99200 13528
rect 880 12848 99200 13128
rect 798 11768 99200 12848
rect 798 11488 99120 11768
rect 798 11088 99200 11488
rect 880 10808 99200 11088
rect 798 9048 99200 10808
rect 798 8768 99120 9048
rect 798 8368 99200 8768
rect 880 8088 99200 8368
rect 798 7008 99200 8088
rect 798 6728 99120 7008
rect 798 6328 99200 6728
rect 880 6048 99200 6328
rect 798 4968 99200 6048
rect 798 4688 99120 4968
rect 798 4288 99200 4688
rect 880 4008 99200 4288
rect 798 2928 99200 4008
rect 798 2648 99120 2928
rect 798 2248 99200 2648
rect 880 1968 99200 2248
rect 798 888 99200 1968
rect 798 715 99120 888
<< metal4 >>
rect 1944 2128 2264 97424
rect 19944 2128 20264 97424
rect 37944 2128 38264 97424
rect 55944 2128 56264 97424
rect 73944 2128 74264 97424
rect 91944 2128 92264 97424
<< obsm4 >>
rect 19747 2347 19864 97069
rect 20344 2347 37864 97069
rect 38344 2347 55864 97069
rect 56344 2347 71149 97069
<< labels >>
rlabel metal3 s 99200 42168 100000 42288 6 clk
port 1 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 decrypt
port 2 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 desIn[0]
port 3 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 desIn[10]
port 4 nsew signal input
rlabel metal3 s 99200 72088 100000 72208 6 desIn[11]
port 5 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 desIn[12]
port 6 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 desIn[13]
port 7 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 desIn[14]
port 8 nsew signal input
rlabel metal3 s 99200 28568 100000 28688 6 desIn[15]
port 9 nsew signal input
rlabel metal2 s 84382 99200 84438 100000 6 desIn[16]
port 10 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 desIn[17]
port 11 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 desIn[18]
port 12 nsew signal input
rlabel metal3 s 99200 24488 100000 24608 6 desIn[19]
port 13 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 desIn[1]
port 14 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 desIn[20]
port 15 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 desIn[21]
port 16 nsew signal input
rlabel metal2 s 8390 99200 8446 100000 6 desIn[22]
port 17 nsew signal input
rlabel metal2 s 20626 99200 20682 100000 6 desIn[23]
port 18 nsew signal input
rlabel metal3 s 99200 74808 100000 74928 6 desIn[24]
port 19 nsew signal input
rlabel metal2 s 53470 99200 53526 100000 6 desIn[25]
port 20 nsew signal input
rlabel metal3 s 99200 59168 100000 59288 6 desIn[26]
port 21 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 desIn[27]
port 22 nsew signal input
rlabel metal2 s 57978 99200 58034 100000 6 desIn[28]
port 23 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 desIn[29]
port 24 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 desIn[2]
port 25 nsew signal input
rlabel metal3 s 99200 76848 100000 76968 6 desIn[30]
port 26 nsew signal input
rlabel metal3 s 99200 13608 100000 13728 6 desIn[31]
port 27 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 desIn[32]
port 28 nsew signal input
rlabel metal2 s 63774 99200 63830 100000 6 desIn[33]
port 29 nsew signal input
rlabel metal2 s 14186 99200 14242 100000 6 desIn[34]
port 30 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 desIn[35]
port 31 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 desIn[36]
port 32 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 desIn[37]
port 33 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 desIn[38]
port 34 nsew signal input
rlabel metal3 s 99200 87728 100000 87848 6 desIn[39]
port 35 nsew signal input
rlabel metal3 s 99200 98608 100000 98728 6 desIn[3]
port 36 nsew signal input
rlabel metal3 s 99200 53048 100000 53168 6 desIn[40]
port 37 nsew signal input
rlabel metal2 s 51538 99200 51594 100000 6 desIn[41]
port 38 nsew signal input
rlabel metal2 s 86958 99200 87014 100000 6 desIn[42]
port 39 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 desIn[43]
port 40 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 desIn[44]
port 41 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 desIn[45]
port 42 nsew signal input
rlabel metal2 s 92754 99200 92810 100000 6 desIn[46]
port 43 nsew signal input
rlabel metal3 s 99200 11568 100000 11688 6 desIn[47]
port 44 nsew signal input
rlabel metal3 s 99200 4768 100000 4888 6 desIn[48]
port 45 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 desIn[49]
port 46 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 desIn[4]
port 47 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 desIn[50]
port 48 nsew signal input
rlabel metal3 s 99200 31288 100000 31408 6 desIn[51]
port 49 nsew signal input
rlabel metal2 s 34794 99200 34850 100000 6 desIn[52]
port 50 nsew signal input
rlabel metal2 s 78586 99200 78642 100000 6 desIn[53]
port 51 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 desIn[54]
port 52 nsew signal input
rlabel metal2 s 30930 99200 30986 100000 6 desIn[55]
port 53 nsew signal input
rlabel metal2 s 37370 99200 37426 100000 6 desIn[56]
port 54 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 desIn[57]
port 55 nsew signal input
rlabel metal3 s 99200 17688 100000 17808 6 desIn[58]
port 56 nsew signal input
rlabel metal2 s 39302 99200 39358 100000 6 desIn[59]
port 57 nsew signal input
rlabel metal3 s 99200 89768 100000 89888 6 desIn[5]
port 58 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 desIn[60]
port 59 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 desIn[61]
port 60 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 desIn[62]
port 61 nsew signal input
rlabel metal3 s 99200 48288 100000 48408 6 desIn[63]
port 62 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 desIn[6]
port 63 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 desIn[7]
port 64 nsew signal input
rlabel metal3 s 99200 8848 100000 8968 6 desIn[8]
port 65 nsew signal input
rlabel metal2 s 47674 99200 47730 100000 6 desIn[9]
port 66 nsew signal input
rlabel metal2 s 90822 99200 90878 100000 6 desOut_ff[0]
port 67 nsew signal output
rlabel metal3 s 99200 93848 100000 93968 6 desOut_ff[10]
port 68 nsew signal output
rlabel metal2 s 88890 99200 88946 100000 6 desOut_ff[11]
port 69 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 desOut_ff[12]
port 70 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 desOut_ff[13]
port 71 nsew signal output
rlabel metal2 s 18694 99200 18750 100000 6 desOut_ff[14]
port 72 nsew signal output
rlabel metal2 s 80518 99200 80574 100000 6 desOut_ff[15]
port 73 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 desOut_ff[16]
port 74 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 desOut_ff[17]
port 75 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 desOut_ff[18]
port 76 nsew signal output
rlabel metal2 s 27066 99200 27122 100000 6 desOut_ff[19]
port 77 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 desOut_ff[1]
port 78 nsew signal output
rlabel metal3 s 99200 50328 100000 50448 6 desOut_ff[20]
port 79 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 desOut_ff[21]
port 80 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 desOut_ff[22]
port 81 nsew signal output
rlabel metal2 s 10322 99200 10378 100000 6 desOut_ff[23]
port 82 nsew signal output
rlabel metal2 s 32862 99200 32918 100000 6 desOut_ff[24]
port 83 nsew signal output
rlabel metal2 s 3882 99200 3938 100000 6 desOut_ff[25]
port 84 nsew signal output
rlabel metal3 s 99200 65968 100000 66088 6 desOut_ff[26]
port 85 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 desOut_ff[27]
port 86 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 desOut_ff[28]
port 87 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 desOut_ff[29]
port 88 nsew signal output
rlabel metal3 s 99200 80928 100000 81048 6 desOut_ff[2]
port 89 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 desOut_ff[30]
port 90 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 desOut_ff[31]
port 91 nsew signal output
rlabel metal2 s 76654 99200 76710 100000 6 desOut_ff[32]
port 92 nsew signal output
rlabel metal3 s 99200 2728 100000 2848 6 desOut_ff[33]
port 93 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 desOut_ff[34]
port 94 nsew signal output
rlabel metal3 s 99200 688 100000 808 6 desOut_ff[35]
port 95 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 desOut_ff[36]
port 96 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 desOut_ff[37]
port 97 nsew signal output
rlabel metal3 s 99200 55088 100000 55208 6 desOut_ff[38]
port 98 nsew signal output
rlabel metal2 s 74078 99200 74134 100000 6 desOut_ff[39]
port 99 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 desOut_ff[3]
port 100 nsew signal output
rlabel metal2 s 28998 99200 29054 100000 6 desOut_ff[40]
port 101 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 desOut_ff[41]
port 102 nsew signal output
rlabel metal3 s 99200 96568 100000 96688 6 desOut_ff[42]
port 103 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 desOut_ff[43]
port 104 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 desOut_ff[44]
port 105 nsew signal output
rlabel metal3 s 99200 85688 100000 85808 6 desOut_ff[45]
port 106 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 desOut_ff[46]
port 107 nsew signal output
rlabel metal3 s 99200 35368 100000 35488 6 desOut_ff[47]
port 108 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 desOut_ff[48]
port 109 nsew signal output
rlabel metal3 s 99200 57128 100000 57248 6 desOut_ff[49]
port 110 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 desOut_ff[4]
port 111 nsew signal output
rlabel metal2 s 61842 99200 61898 100000 6 desOut_ff[50]
port 112 nsew signal output
rlabel metal3 s 99200 61208 100000 61328 6 desOut_ff[51]
port 113 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 desOut_ff[52]
port 114 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 desOut_ff[53]
port 115 nsew signal output
rlabel metal2 s 41234 99200 41290 100000 6 desOut_ff[54]
port 116 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 desOut_ff[55]
port 117 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 desOut_ff[56]
port 118 nsew signal output
rlabel metal2 s 97262 99200 97318 100000 6 desOut_ff[57]
port 119 nsew signal output
rlabel metal3 s 99200 39448 100000 39568 6 desOut_ff[58]
port 120 nsew signal output
rlabel metal2 s 43166 99200 43222 100000 6 desOut_ff[59]
port 121 nsew signal output
rlabel metal2 s 59910 99200 59966 100000 6 desOut_ff[5]
port 122 nsew signal output
rlabel metal2 s 56046 99200 56102 100000 6 desOut_ff[60]
port 123 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 desOut_ff[61]
port 124 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 desOut_ff[62]
port 125 nsew signal output
rlabel metal3 s 99200 15648 100000 15768 6 desOut_ff[63]
port 126 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 desOut_ff[6]
port 127 nsew signal output
rlabel metal3 s 99200 82968 100000 83088 6 desOut_ff[7]
port 128 nsew signal output
rlabel metal2 s 22558 99200 22614 100000 6 desOut_ff[8]
port 129 nsew signal output
rlabel metal2 s 66350 99200 66406 100000 6 desOut_ff[9]
port 130 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 finish
port 131 nsew signal output
rlabel metal3 s 99200 26528 100000 26648 6 init
port 132 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 key[0]
port 133 nsew signal input
rlabel metal2 s 24490 99200 24546 100000 6 key[10]
port 134 nsew signal input
rlabel metal3 s 99200 44208 100000 44328 6 key[11]
port 135 nsew signal input
rlabel metal2 s 1950 99200 2006 100000 6 key[12]
port 136 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 key[13]
port 137 nsew signal input
rlabel metal3 s 99200 78888 100000 79008 6 key[14]
port 138 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 key[15]
port 139 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 key[16]
port 140 nsew signal input
rlabel metal3 s 99200 33328 100000 33448 6 key[17]
port 141 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 key[18]
port 142 nsew signal input
rlabel metal3 s 99200 6808 100000 6928 6 key[19]
port 143 nsew signal input
rlabel metal2 s 6458 99200 6514 100000 6 key[1]
port 144 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 key[20]
port 145 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 key[21]
port 146 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 key[22]
port 147 nsew signal input
rlabel metal3 s 99200 22448 100000 22568 6 key[23]
port 148 nsew signal input
rlabel metal3 s 99200 91808 100000 91928 6 key[24]
port 149 nsew signal input
rlabel metal3 s 99200 63928 100000 64048 6 key[25]
port 150 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 key[26]
port 151 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 key[27]
port 152 nsew signal input
rlabel metal3 s 99200 37408 100000 37528 6 key[28]
port 153 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 key[29]
port 154 nsew signal input
rlabel metal3 s 99200 70048 100000 70168 6 key[2]
port 155 nsew signal input
rlabel metal2 s 99194 99200 99250 100000 6 key[30]
port 156 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 key[31]
port 157 nsew signal input
rlabel metal2 s 94686 99200 94742 100000 6 key[32]
port 158 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 key[33]
port 159 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 key[34]
port 160 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 key[35]
port 161 nsew signal input
rlabel metal2 s 18 0 74 800 6 key[36]
port 162 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 key[37]
port 163 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 key[38]
port 164 nsew signal input
rlabel metal2 s 12254 99200 12310 100000 6 key[39]
port 165 nsew signal input
rlabel metal2 s 49606 99200 49662 100000 6 key[3]
port 166 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 key[40]
port 167 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 key[41]
port 168 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 key[42]
port 169 nsew signal input
rlabel metal2 s 68282 99200 68338 100000 6 key[43]
port 170 nsew signal input
rlabel metal2 s 45742 99200 45798 100000 6 key[44]
port 171 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 key[45]
port 172 nsew signal input
rlabel metal2 s 82450 99200 82506 100000 6 key[46]
port 173 nsew signal input
rlabel metal3 s 99200 19728 100000 19848 6 key[47]
port 174 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 key[48]
port 175 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 key[49]
port 176 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 key[4]
port 177 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 key[50]
port 178 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 key[51]
port 179 nsew signal input
rlabel metal3 s 99200 68008 100000 68128 6 key[52]
port 180 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 key[53]
port 181 nsew signal input
rlabel metal2 s 72146 99200 72202 100000 6 key[54]
port 182 nsew signal input
rlabel metal2 s 70214 99200 70270 100000 6 key[55]
port 183 nsew signal input
rlabel metal2 s 18 99200 74 100000 6 key[5]
port 184 nsew signal input
rlabel metal2 s 16762 99200 16818 100000 6 key[6]
port 185 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 key[7]
port 186 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 key[8]
port 187 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 key[9]
port 188 nsew signal input
rlabel metal3 s 99200 46248 100000 46368 6 reset
port 189 nsew signal input
rlabel metal4 s 1944 2128 2264 97424 6 vccd1
port 190 nsew power bidirectional
rlabel metal4 s 37944 2128 38264 97424 6 vccd1
port 190 nsew power bidirectional
rlabel metal4 s 73944 2128 74264 97424 6 vccd1
port 190 nsew power bidirectional
rlabel metal4 s 19944 2128 20264 97424 6 vssd1
port 191 nsew ground bidirectional
rlabel metal4 s 55944 2128 56264 97424 6 vssd1
port 191 nsew ground bidirectional
rlabel metal4 s 91944 2128 92264 97424 6 vssd1
port 191 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13726218
string GDS_FILE /home/baungarten/Desktop/HW_TI_Encryption/openlane/DES_Trojan/runs/23_10_30_20_08/results/signoff/des_Trojan.magic.gds
string GDS_START 935854
<< end >>

